`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UeUQOSqc517u4Gp21W1qcB44JkXjttQw3I9etxLnnrt3tkJ0d4uxhbBwSkc7IM9w0xxr7owGLR37
1Ii0/OYJsQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kOXgzYTJC4GxJCP3UAJekjjYLOXKC9b70sFPvaIFCHz6zbI3mz+JUFPTpADGukAuJQCKiXWwYOBZ
MmBb8JugLkKE+O1iqIjgnplEt9Bnnc0cPnUeT9o1Q0bWLLOKk75pVanxsTWyvGhO5t3dBcHf76mm
DceLRrUeM7AAXcHNQP8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JeQtyj3Kal6oTj33H4A+stJ+V3DCiNJv8J7k4H0+dLfFYYJJ3jbUoUt90xE3PJrsmjZDUKwDIVOX
HWBDaCL3u44dq/L0M441Q3RfpW9QQqU0ai34/xEtkAvplg6Oe3ludzsYQZ7T2bjYDyh8NSDEu4PD
/ngBWkp/hfXUBkMQq3g=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D+mEShAo+idVddojD4Ocf30d3PeQsjyupmNQjqsNdbpJFSb9AWyTI4HLKIImT0S50Zgb6LGKxa9h
26g8vXL3CdbVdP5O8FpM1809Abu5sfhEOCwdvtKWRwLRZt1+A/6C8nMHuYTLwrt4lXg1bU5c54n9
i12z+RFxTTeQUgM++Sl/RYKl7QJ7e+6a2bvs7RCI+NDk3Qaeos9nT6roJnfx2wpYOF4jStxFa2up
F5q2mhYTDOmLHpkBQCKAWc41vFlv1ZeWkv5nIa97hTbbuUW8GmJEmxKYO5Ix08oKP4QxHuiNF++X
v0t8M5z/+3rsLJl0oKiKofyP/dx+okR3PXDIyw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tcnuNu53+hchNr+pZ1NtakfiTYoR6SYivYJdM66R8/4XDELZLm46FZjh8e2MDPfDIe0TPxgXssIK
JBpdVvHEF3sN4ne8BH5Hig1m+5eYblKUujpGtmIpXovQKiu33+xi9YvN+S91R0i8O+wIG5Y8ZtSd
416fkpAXIqKUgtlCKXBPfNKh6pXB2wSYbWz3TlPOiCZhgXOn24ftBdQmq794Zo6QdyiBWEIqcHvf
cGxpfdy9soUWUFDgRcMQziQpv5Bf40FoOoFPc0PTxzAfe1PMhPuWIOtJwU7v2ehiljl8zfvKr43F
vafnOBmYmG/WIJ2D8gT8zcjKCOuzkEZD4/6LHw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CtAJ5i2Ss06xmVLrV4Tdrt3cQho/pCz9fbTCKJxQdDrBclu8FdA7n6uV/sbGH0tMaSievrFx2Jcw
lrfRQgsQbFyxSpn5PUFRabLV3UXwVpPqRPFv60hHW8dL6EBKTJRiEKGMFV/9GNtBclnQParE68gy
UWIYfWYlfU8odNKh63v3UlbKBdSSTudb0Ul16UHMxR9rOEcIVol8aLIxFF0XFN3SbjvZQYMrSrda
mdPrPZ6RZeEOu+2fjH5DVxI6YAiec9k48XHplaRfVHc5p6pbC8oywpPPg+e3mzZanroV2DYjAywn
LeUIPZxac7VkB/2/ioqm/Wqs+AR5+6YLStbDqg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558368)
`protect data_block
v96vx+Xnz5A/5tWt543ByRzuBusLYDqbkrt6yfkEXdK2qaUgm2Bn7IgeE1LGB1KJTnHGvrg3CGgP
qyDz5+jXkDYzZRQM9N8C1PU/R0a4RxEY0vuaAnwXZtoEVR7m6h2+0IeOoBQwqUPHpY6hevZPXY5o
fvJRJ98ZvjhPUZ2/a64Ou7qVTrhOvL7WkXvoe6RZK7zk3n/1Mu052YFDS+IGu0pix6f6BaLlg2YR
WQXFz4KDxpswDig/vWv1L/k7PYWyhUx7LvlvOSzhgfKBsoVO5lUneCjVfJdse1x4wRgCUyKo7iLO
Kovcw1MOsel+Xgq9WdCu4GF9H3+VZWTScbkXI54E51mMCcafDhLlxc4cHPPK0FTXTHMUKWGCqJuu
tky/LMRE5c1+Z+juXOnhAiX7+8CI2ZTkopQd4pNSrKXWpWuMVO53Pnt7pLhYJZaJUH5UIEiwii0j
v5tsDySGFMm8sB0QDSRw9wVj3UsXjyo5jqt+fzcRPzY/0ZWTOpE3cduYDDYpPcyw6AUjnNbK2Jxs
pIOyrFBOy+V8MaIM5Wqbl5zrOHIR/QpPOGwLCrDk4Ulj3JDUy2DBQvfeV6vr7boPK85ntIhe0+Vf
aBvypRZmGXP88HrIW41XysykSCxpZmVzjnA6jx/uludh6bsioqlcjIepIv3D9nLHyE9x3S1fqZQd
m6fglG4xSpmYO184R8nJs3btNH5RVAaHy21RqlaySqhQtlJba7JD0nu02dKuXInLvaA/PA2psrkx
sAOUjqa2nKvmUalIJEQhyR0g4oG6wOdmY4/6m1jFauZUC9DH8dihiu7zqZ2DZ4Zf/OJZM7PVURRl
8cJCYhMSsvy6hG6aFQtdN4HRypaoVdhV3pIr+FIIrZHPg1VS6ImHWgiNUTpUyuNlL17pcmOVk9QU
Tz1hJ9aNESM/XHKyxqLg0SpjL+SmPJhh0RkUAXFbtCbVBdCQ2grMq6HIk99iJQjsDSYbRlfupvHs
cxOfD/3cn41dCzi5fscveEc6f58a6oYogutOekbDyZoDPvQDoY7G90YrJLYWXMbVG9CwlS9n3QvH
Tqh8r8ALNV8zyUNDg5uUR+dSYg+K9AHtHKTfIPrvpsQMmfjPP9RKXD4zYLu4WkLSk70K10zfsN6s
wUYIYfz/8uMh6j3W89RjL9d/BCjFCA3BkE1qu80ULFuh1XXJgirS5FLQWSK+FpnzMpI8o09PVdNJ
qUF22+Fv0FscYXwO/y272/DATloJ2a3X9kVbSYzn9k1odkb9m208a7WAZeGcCo0B9R/kzlniHovu
WtlpkLUBIvCgiPCUukiozJICXGimts2DZUBxPVIxvrAvHUgFg2fb6AbZQKVvl0H0S+4iX6ordzr6
ZzMoF27ADvwhYhjdar8gAvcKn+Jl97BV37UywiRJABUpOV7VdQCacRra1yvVnIE4Z44Ve1SdYP5j
lLgGTpSpc/fViWF85s8ffoG0EcF5KNN100CMednuay4eoPBGpD5vixM5qzjfbaT4rmG/SFzwMBk9
QMSeyFi/v8i5rBaSE6SpdfkUpRQVgkhle5m3hyyjOuCYoupOvu6QGZKpj59dqebPuZ+FvfGzbJcQ
wngxZfqceKnn48tmPD/hjj3iWBWooR+VaAyuZIzKC4HicL5iW9MV9orGhmb1FQ+NA3wrMWR92GQU
0kdfRSeHQi3Jdb1x45PShHW3GqAD1Fx5ZUqw+GTxa4HQAsOSDsWhU1HEN2rAQJnQFCZOUTUkWMJ7
5ogdo47sLbw3kXpxTS+bzAR1iRzSsvCOVaqFBwH8xgwgRscvqtW90KF/KbM5veb3OG+4bgCLzAvd
ujcQ7nsSi7m2xHI7beqFaBFqIA2zgNMnM/ZI2IJEQogLM89sKSwHtrGkD8cpzzkfUskHb7uG3D6H
4bBFYx35PU4Fli2Vk4tFcO9xpbzm5ph15SGKX/sOeZeSrBkToB/A67Ao5ulpcO6RL4osox0Z5bmZ
Tc9ZYlcKD+TXmzjAIFxzILjMYmEbu8G0t7mkEErZd/yA3gdDYJHqVhkOfz+FYa/orA0JEc5oegOO
M9NllKWwhJ0fsefFZPKpPPEy28ole8CxR+18GlBJBznklusWV38L0pN3OOA6lAi7qK8sCkOH7GbO
kg9JwkVpaW05K8q11M6qcks+bxzxT+e1a4irc249B6Ha+b6KyzymJD5wGN0dG8PJ6CWxpj/Qu+I1
mb8owaMdZRusskm7mPEEuIhVF5HpjWQ4HaAPlgKeM8jEQKV8gObl2s2Ypyfjivpp9omdnx8whnSh
WG0xkhg6OarDI1osiUGKHJFZK/D8iJCaOVgcQuMbXkwFLNOovnnFuYlLb3y0wPTkgXUTi/xUACTA
CVAPIOb70SyQSGWPyLV0+h0h8nENoMxu2s2k1HoiopFVpV3RK5/dhzYkCAyy9FKT6e+zWr231Noz
wc3URTt+b0DqNLbPd9Fr6Wj/rxYW59eF6562sz8HeUF9I98WBxkSpFaX22dwCkpzdyZO23LD7STx
wV3eUBsBEHIKfEap3w2mPJRIg1KSLFz1JDuHUERWcXFI5gYj3+7jYoFn2ovm+chogx/L+WlyREz2
HpCBMg/pIwEJDgiYwNjrvZuc9JvmOvbnIUf+v40YkFN+HS/JmVqSMngvlvO0mAiZfVrMM+KMbGPe
cgXeymuazZt+WV/HhtmP4+G8wL+o1LXvvlz+GnFuOHocY6ma2eQp/3A9E0XNyx/T+WOPA0LCTVtb
eSBDCKuBGRJxF2RY0eNlIDfYo0326gbeZONZbchwYIbZa80u/ktFFyuqipqs6J7+tygRIXjU70PH
t/ZIMFiWOAlzJoifCB6MaG/WC18mKdmpdm1pD/n1UZn3k2mc3tiuj3jHNWvdKaSUCHiXObUNU65K
KHE7qQ6yJDM9pSdqZwPQ3J3c0JxGctLzjNc0tS5IAW+PEgDMdSUPjoX8govh2GKUq2L44kMnFYAO
zM7Q8k5mbZ6xECcdpABzJSfDJxvwaLKRWfSvxc1vt8s84YDW6EzTwOG/k48qXzRXGWYzFzCZdN5k
Wbj2pj8JdFatAQjZbmTrq88T2GBiBp26BmUB7eG84H+D6MO/vfSpWN8/inr/PWOeqhxS3B8kMoJN
xf6btafYyryCOSrhnKVSJMl96G6SCZjbq02R3Tg5grMd2ddSi7bMzAqQppt3mPu7P5t738aTzyYJ
LJ9uGjvuTS6qdF+deFu1viX6PaBPVkjedA71uIUil9DMjHdSF4hWZWCtV/or6BoybnYx1hjiFGup
T8XXgtFjU1iRALc5/tonuNylAzPwSTsq1jt3KGX6LANcaGlcGgILHsfkTqN3cnFXxD8YvWxzcFJd
f03KBfHRo1gc2NphU96lOUPCChVnQFfrE/jYbv8qWJahzgU8Nz+dnuQs4wZS4WIH6OgEz3nmUayw
E/Jcx+Kv0I80oUzE8TfSXoBPqsqxeyEBLeD7wueevp+E+mnAiohOd1vDLlz31Sr7psHdsQKvzbE7
kzQF7xktd73peNOtz5y3gZh5K6votTkmjJrs+INwYoEx3JOQVL72DBzXh7az9q2DcIZkuf7B621C
2sg4dFlUiGGlamYmFFOaUNIQ0OA0uGeWOBMpt8TjBy7vyIAiQOLqehwBXva5zmD8fFWcgVBE/qbw
/KtoJYRBWOAYJEg3XbAd1yCxDtG1tLSNGSDHj7sJc2NVh4feK8/GLE9x7Tu2RR3AfgWVo/6Ss7C7
8pq49B4BHgAtssT8JJQ9NhCZTLE5oOszge7vkzqX0rqVOrSQYIgZav4yWN/wA0v4D2Jl3WHHu+qs
5kqvBX6Fr2dsl+Inqa7VwPShSfj4/iWbgag4c6INcPhIPMkmt+6XvwQQkpPSdoaMdBOLfPVNzwEJ
gdpkSaC7ucXZlX3gtS5Ym3BlPiUwIT6OM3RdAqQz72IclKhO+30qoLwAYlvwvuyiING/+Jm9reDM
jOBImD9ggN4XlAuItuZQ/PqhsHtYL6oClwmx9xpgtz8MBo8bpIao+wyUEoe1HeBDqbZbZLKlhHDE
2/U67m6N6fkzXdPrjVUj9aTHgwSzo7U3K8oM9jo7p+Sk6ncagUGGXzqaYalnkLJpn47m/MG36i+X
4AJRccIJHDjRgYVy3bnWE4Ctg91/6O5H3aD429jp7Ck3TmFL9cvnoJDvV/FyedZKr1Xy1Bq8JxZV
kMBkguO03a3cYRoelY2dl/LnqU7AE7RiNZJFG7XP0XcCHOw68j2wDcJxbixRf88+4eAVhKWYnsTy
xB9/vgcJLoXDFi8D92yGtLrGmxHVuhMKUgLAIQpYeKpLDg89LTD3Afr/cfWIQXdkgr11km8IOojb
W/qgk9AQlKgwqR15QK6l3if3/6yM7LnvS1nLTOqSOhD9FZY4u+K+hBbR1K7xFgPx8mzq8f6Fb4UO
dMDUfjlnzkEgyZhfsept8EnFKGZGyebcJSarAoqA5eA7CZE+YKCfk8QJN5Tb1Pni0uap3JgftLRC
7q45JTRMrj7+O2c6f+nFv0sP1AI9a2MHVOvnmFJKRm3DIPdXyc4mvYGjCLmO3X6BjoW7by/NFSMD
A35JwcXr7QDPZnnSMTDcxx/jm6LxBpZmI4HyTve8rcLh4sNaM476hda6b6jp/iWUIv0q0pQW2hhz
A1sBx2GdsgtSh/s8eSn9yQ/9/ylOWgQXP1oJGJv3qYZPV9tcaf2EeGub5kVzL+FpVSrKAfOwe9lv
hgbBViVuQpPfYG0ppeCGPM45EIys70TXbXg4Lz2vHLURUKcvQj4ARpCGqIaBPaay9j8BEMJpJi8w
CWFvWf1T2UfeDDAHcEKGQJ26O03JTTk+3zqCmfZDzKFeM/KrhYyta9j9mHACFLrCXGG2ic43dgBU
qYHnIresZKF3smBE5wYWosjkGVVOrVHiA+xaUAjb/tOJb02+njcWik7CPUqYQZFfLjbdLmjpKvy1
Zo+tR/PZUOEomACCz2mt2xj0kz6yEJ6RitWHyUD27DVWWHtw7YQRrRoFmLnuBWh5xWN0BmrMkhb0
bDKOVTvyE22verW48RtIatO+mkM6ceyeYnX+VHihsGrPPrSVPgtCllMJxdLmH0vZpkAuDKwptc0e
43cskdgDECnOxM4aeP692qzwpRHAkWQ5JF3iRqQVpvOuRD/HEy7mZJ5qM7FTnbeuoUMJQqztUPj3
HvRGnsdsnwBNs4h3DecIeNG2XzrK1quW6Zfj2EhYofSyy6sYvNs4t08YyXgk5elmU2LZYF0Q4MTv
BPAqZMqSxss7REIDsESVFo0tFBwjdt5Ra6w+I3glWphGrmXvGgr4Q1QNGZLNT0sx2XR732VlHqoy
5pJifaLLe3nRHUVSpZGCPWQ2LbdtgnqX2O5J9nXzu37ib+2Q7VBO5nxKPnjO4FaoLlkHFLgk9SKT
I5xN2ii1Mcu2qx58+N88YuOHCxRR7wQentbYqc7m6wSw7bixSt3nkqfpPTqi/rWNzneQ9FmJ+nNw
n90R8D5AQQibnieECmWHwTUvT3340hpWdGo7fXAxjsfJZON7UqrJKiu0taPFMt7Kk3YasLMPzkg5
8Zox0wlKe7AO9shXFaxuW8J7bxod5FAa0IngjiwGzcnIZx1I/TyWAqlKxIU1Uh4YAws374aRo4fv
Z590Ys3RwcQKW1FPkqpf0kiRuNaOndA5oT+v7cj0TfAtY8jv0ILk13MAUBbRlc23aPe183Rb+AAK
ZS2TWboHytRZoOqV6tLjinkQ82eph9t7f8QzW7vorylCizyRfUk4jDA6tx3nBFrDkQEQoAwT6zeZ
eiWDQcz7fcBZo/WxtbV7dspXEbjpsLYKyO2ah025kgUaaNRVBfpM16Lapol66efrDFZVF+13yRy+
lZ8PV/yFnM/kyl6YECb0tP6fBdp50m4WRFTwLBi/RPW4WDbOZITyT3L149hny4T9mXygtef7dLYp
AS78uAyVcS2GDwPkSePm7UH5UmE1N740M2KRU342D6gC38vxozNAOKxREjno+hCfAV22xzJixrBf
OXaC+v9SKsjb9nRYC5xMIKKEjv1Rw1gdK5Kc06YxUC8hiV2RTa0EUqpHx8rLn/WmcToJYDkAZe/S
ON0SoMRT3WV3DeygdggU537TmeciAqq/YxqQgyxnVJ612LM4x8XNUeh+opCu9E+TrommlHepGVMO
mYSDFSgDoAT8rm3vfZHs/JeW4fc8OZF3Y2jIxcPd8WvsZl07uXACqrgEcffCWxJpQac/ekWi+ofn
4pbY+SJBJuiOgFxxbXlvlaQvsynm4I9drhZB2MrnT6v67+wulmq53YryridFp4NnpbgybsRKb5zs
8S3OhYQI1dPrgKfbYmVzD7oU6ffWaGchy38Dlie4VzjRx5lk8LVtCKAJs9WszAtqkdmlaTkTkTdu
cUNQQpf5KOUASW+d92ppY//lzSXceNbluYFFKP9V/OwXJ2yjzi0oI7jUE33YMoACFNFP6YFcLLCK
S/VhZGZe0jc8rNdjbQWA3/A2XdzI9wsgB94ybtZmzXizzr46LyWxwYcRlwfsTz4zmZr3FJdAW0CN
40z0Sdzg9uox3qRuPRoApmV3ZmI5SoSccr6PdGpt+mkIb5KqMvqGpb5swb914DEY7Lar5L36rqia
fSbcCudeVcZiFNmxKP5sLlR9LBrZym366eITJJfBgw8LgvuuJqgIzyroEHH/cQuQZRRXFVr75r0D
ZvFGu8q4VECY2dWWiUHK2BaKOUoUJAQDkoJxKhP6OHsAfkQ40OsBYYPweGLLfGTj7q3Nw2TM9xN8
U5MYgk4eiUo0qDVPM+xdX3mVR4A4c+740YQdMKyDUIdIjgK6YV32vF28C831BfgnGvNr0yrbSIE7
+etsIglUndD7NKy11+GyEgWBQnTmkb/nbLpJg7A1JdLqUWTEBY6nCFabG6L/ImQWOBeLin3ksMNQ
BdQWhFrwy0rIz9QN1cg7SgoAHEGxIICpTPfQYiF/u0NFZrtH/FxhPqQxYBEPwetYs9nod/BSc2mL
Bq1W6DDfNGuG5/4q+wOlsg/Cg7/fKYjDZ76VldA9DlrLu+UWgm+79L0IFB585IROSLBT7SRplpl+
OTq349MwL27hb5pPLxy2qPvrG9+jPInYfDXyvb9nPBC/O9cEJTP3FpJkbMgr+G0dVHqBZbv+EqH4
pKislw6V2fHb/8uOBNmWK07OBLRzDSkMMmrz40JUJI3wyLtZR52offIec+JZNqlRX2E2+WYcGxAC
sw6IJx6S8o61cgtVl/4wzhwatIbS0grmUOz2qVMA/Ep0cycLUnyQkvPnZIenfQJJy664nH+MnXk9
Drw4nj2RoQKhuH4JRGAd/taOIsV4kKCaNQptZdGTXuFQ6KE+2zkQzKkZurzy5EoMaLZBXZVB4pNb
tJe2TF30gE+uU+4jpL0w/sBwNyynkBzJPCMh+qFmcBDPtgaOO0OnLQX24GpFJ1VQOiZdKtX2r1jy
TVad6TwFVXkyZ9RTScvdPNMUT6I+03d5NhI7S8vnfFo48eTqnfdr7rWYB9AnIlCpDv8jjpSDMBzd
ZOtKzd27weR7hE1RHIU/fpx4MI3msY8eUF85b/11SDJXiKefDKsE5vAa/qXacmh2QPCN0b4kjU95
ZbIvuvO36dxJ0ER9JA4Iv065SnqRQ6T1EapM1a2WxBJAHvB3aeo1UNWS0Npz0VSGizJyDwCc87gd
43y2nM9Y1FuSV7E8X1PE2GsExyGzlQ/MakiE+kHWEp6SGnLxW2xh9aDU6ljeDZnKhAQe0Nb/FCsS
ifejNfn6QPrqIVU4r4za2uqMVDTD/jHn/ypq0zpvPubow15tAyXMypm3FjTBx1ygFPOm880WSMIJ
sBaxPdB4+7GdRClS/UjdnfWWd8BZkH+9iXvMBnKfSA1l5Rl2vHNRnYu/8hLsauqEShzTgntLRoS2
4Mqffo54lvHEZnxAto4NKfcSUgyhjtNbbRYSNtg6RcoSH40CQim3tDnuGWJ4juALXO+OjIhgSmZ6
fZcy6cxX4Sfi58ZhGMdn2eBwgWcvk+4UzuGT1dtzsKCUCyxI3bl5/7jpwfytj4s+9hOGYgL/dcTF
Iw26QsEw2BGqqyVStThsH3I+WiXuOtFWI3HRxvEL6Yiie0DRBrHuWFGNKM5eA+l9kvA69xSZQYrx
dN4gvSsg7b0zDrkGJoKkfSFbVfLFlOeKVshg9BL42KksbnE3c5IB30MtsAekbKO2xJU/jLnR0j6D
tt8CSM2+7G/me61hNE5OT2H5CjQF1ybPpytCtuApcMXVlPeSI9xvLzIxEQPvFEFurKMoHyjY1LNm
xrX8LmjhDJtq3bUgOdQi7QVZnvgYjYN5CKy1R1xKj0Qbgfvjl/FXZ77IRH5mvFeooTZNiTCGXfgl
+np57CGKnVBSeRXM0Ovo8AMm5nKU6Z+awsC86P0YRoncJcOYnhETjE2Nd95e8VzUX+i0A9fqEO8K
R/mKS3tPYAVvb6HmElvOquToCClQlk9jTOywbb/1QY1mAyeF79xc+QOH2LQrtJDTbVKrPGF830bW
81MKVPctojaX+qH/FisO90mVTvJfTH7Oz+GPlsLSLW4I58CzFPz1ZvnH+86Ndd4URkySzJMQOf8C
mYjbqNWc1KpekDzaD7ZB3Sh17Q6aTYs2FhhVPhPQCGjBWgnr1CmCt2WfMNV2zih8g+azVh9MIFFj
w+UKd2X8RpUhSKI2GyWuyYARye9WVw+BOaF5xxlBbYjWSW3nQwMMvXoLbDqfau28CAaAsz3f+cjN
cn0zSLj96Ika+xG8hGEpqf0bx8wHnB4dkZFwHaGN9B1+P/8nU+hLb5LOgFCJuuQ10n30X67EmWeS
Nwp42s9aep10AkhQ7EOyWYgM29T4MIEMp3NLILz2HZF/Lx30gcAK85bWRsGuPBv67psx749hd+B0
2Lms38uHD6qNji4BvTMfqEgBXDSv0LWAcI/8PxOdqbPBvrqUAmKAWdTQ8+AkWmHU+NHjWQgznxc+
5pSErJa01f83a7bQbbAIndC7yXvVDZRdwQGc3XtiS4rYslu9Eak20cfCGET95F8e+vXWVFxANkwV
13x6VK3fk5weyrXwst427UAKORy7EDmklz0/sc9v4cvMBvebEL0bk7p7bZ5FDIjBKcFYMo97gyPy
4His3yIFPJ5j4Aid8dWr6zJ36jzxqBTr7tqTsGGonAz5FnCccx0B/zUFdZwMnl2xHKKrnMdXSOKj
1oZ6gLAzS+UGUZs7OPfQZl3e60HNxmKg1WMXpNr5S0IvtARdIhbi0fKwuPvO0Z3OAe1HMBINVf6/
hacfeDtBBszmc82+RwRiObU7dmpOywo+F65Di5jpcKnBF0ESsR5o0K6c3kqMvXa8XHToNOjwATdM
gU4IvGOkhzCTqTM/296KjuUfDZAP1V+EULp4LRGTunun/TahkmeKw6Z3OV3FZltHdfFDdkp4SKmD
VoGUwnEAnLyYwX/hrmcia6wWELrGDx4yy5Ak83KZmG1XmPiwsx/uWaTTQ0jdimh6ovr2a7uuPLgh
Z/+jRvXthXv1IAt+l7ycR7iUFxHWVytnI9XQao+fi4HkSFqj0mhlNnv29xH21J61aOHmlUhglpUF
wI2wsAmQXwCqA5VkINqZQmWHMeIb14bBTIoOTNki7wY+Tuij4nNP4OQZoymjHlYWbCsERxrLzm5c
JuLuZjWWVrbTOjdMhFKxx+1zUcyZnwKavS0it8WcBQ+iYY1zVZXjquUTcRDZYsTvumXZDSEI4zW+
wzhAJ5N8ZW+5ckyvkRnH3IHmveOmVvWta01ZTmbiMTaT2kKi6GF+TxmDGfdQ/zmesZQM76r2pPOl
psQMRWuJo9vhy2HiKhWc+XDAyRIrVyihyY5pH0ELnb0DQnVsCWK6dwdVAPMbRnOVwGwoHw1oNZTU
602pkRDsdJ+rIDkhKvQRs1m+qMWs2goVuZjHBw1/QAWddy19jrT9HrpWxJ66lnSoodRmPzrB0yqA
yFM8iO7jvlMDudzFKmVJwneut0LJKoEZCfhdRjrppst7M0sJJkU89fnVa6yr44xE1yWD3FYC2fkD
suQgj4D8qLGVIM6aFNLwkYqCeHW58RIF7Tx9Ak5ZoRCMUXPdq6vH7Bsp1h1mzVfmeaaXpkcJDpVZ
bnocqzjbZSvIwYRRASMGK3ymBbA0w0IQ6DLIU7UStapCp+xfdw0x0bY8P9jp/NapN6ZnKrJs8Hg3
4u27w0G6AqRf+Lkxn0PbTC7r2WmQ7Px8c1dHtThVc8c46ttzpUfmDB9FuP0ggjsWhCk8MC9QMKzC
MT7bmfmsn+fl6WWkxFuBo+q+ZRCmc2iqm0SM5v4Jr9PieEPtZtGhgDvyLxYFGClRoEqe8gXhBeBD
R77qQpefsIlQfhsFoy9oE685RZs793j6/cy5phCrCp/Oc6r2NHbXK+8ZcT3+4ulPbnkrc7DMGwH8
ZXtc8EydbErzVgeoc19CHbpZW/KBmIJ5iGU18m4RwwM0nNr6P4RJB/Z7+Lk1J7OwSrNpCh6Rg/5R
E0bH+obgxj80dWrmbVA3wjkIwFDQvekZs31dfywlm5bxsukhchAyIuDIDIk3QzLCmdcaeY+Rp6nk
zOumIH+G5MxJ7/rOFThZY1onKCUv6pvTFfzRMd3RfR7ZzLtfygGrME2EIrWnNbhnYm8hRxv6lbhB
pH+ew9rVT2eMxhl6zGFtnswW3IpWfSaYcB6+B5ZhWlc0NmIQPMTn1J9iR8ST7mzN64uJNIsnfItt
dASamGOhZsTVcT23lV527MXOs99wPEX7NjL2h1gz4zu/7aVxjS/5Hi9CeBYVZF3NRVhV6makQqeB
lBndMcGDjT+R1Dlgg9Rh0sUqMAY6Fp1bKahj7Gwgt7N7D567/MUJczHX1HfPsV/1yltZUxqUTtTe
+2CIaJl6xndOe7nmfffvKP07HYJ5FMzcYT3bPzc5h8IURz72VUZ3gsx0Kg+71v/kJ17nd9KcxAJk
mm2ryQUj8sycPMkmNLqxWlaV3AqDF6x/eZYi+CO9nlOJwVF+sgg6WH99LQABq4rChPeR/3TL8/HG
jpw8Sh/mHOMQpZ2lKEzcsxQEv4kjdKF/9tpSFVRop7uYC+Bt9Dp+sosoEnZ6z3XFEY5JjHJzymwL
QOzV4WxDbHAz5/TvXbAx8mnidfiX3bW17ea+Fj9QI6XxeTCHQpdpHo9fK9MdpUMhTyDqvqyah3Bt
mwYZesh6ZW6mx3IVa0K85zzfdrErbA3DL/Ut5/r6HPFYwTshwgt/eQTCeIXtcEOkz9vn5N97jJH/
+XG9GoqVJpBy6HfHcV4JhAUNz49Ju16mjqdURwVs1rOzqGwpJzj3Pjo8Gr8S3dI4LzIVWAv478Sn
SDgChBsus98ZNeYUYOAmaceAtPt3pNoO7Ldxa/gFcbkIlxXzBYd79/LtpO6mIsEocf7P0Jm/PnNM
ccmfEzGfmmfZuHReSRIZQpYwMfq7sB4v55uhy1CgjUuCH+7YGhq7tkUrDdg5GvS2BsVW6CuL3YZI
sqgmsI8637lItQmgDA3GY+p5HM3fs8EdVlxhKRcJqbRBejzpVVZtd0oqSXeToDmfAd4w3Y/lLnHx
XP3GcmZE9xlLry8mxFLxRqWttCQcFxB28+zTOMQ10MsfbLZFBvmGm24nqIwOr9Ymx+qHtm61Z9aA
YxpDCHOQpCrjjeY/ONSqRUTEJhG4LJ38I4F9uN45VMVuwJSccgXvlwEoI9dLQta7ss0a8HVxSrPW
somUU7lDtYfsQVN6IzxR5mVy08TIpdpSXhp+ZUCvm8fH1EVxT3PC78pKzdMWf0LgZRk/qginwgtD
2MkN4CmI5ZBwc9c+k62jlbL4tUM9Sf5e5W672QaDY/hIMVE7Z6SHIAe2hc3AF6/PgOU25hGgPD/M
eLvqCh50zvsfk7cUzsLKGYdYCK1hUYUAbBkcoaZdUpf/RqVB4CUepwhCt+aBQw6tXLZk2e+DcS0b
DantxqUby/1TKwqv+eE+Pk/yLwBWLX13L9GY+d06LUFHrDJV3eeLRTtTSOw6XcHtc3oWz/vqnU7q
OF0SkfbspwFqqQ0YEPDVc+uYOmz/EMrx9okcx2jYfNNmwgHuLVQGbOGnb1/2PSFRSxsTGMHPgrvh
CakBw8Q6k3Zi2R6SQbNUGh9KMCQI8YQGfqAduy8FSeraNyR0fUMksdkH+0mHYjCTy98cvSmT8oMq
co65+GzRPb+e6+ch++nPxXN5CnzB75j+MIXPmcVxTjIQRMh2BFYyou3RbnI5r8lFEqLIv/Y+/3ko
aYEMQXLh2IXshZAyfE0KB7pFyVM5CqAHXPNLRsGI/DfN/cp2ASMz/4+TuCUi+E1HA7YnxPULHWkV
1Xp8yM0L9brCfyso3WadYSFSjdc0INtNadPqs/Bc/7O2zb/LNkA9qaSM3/5tHiPz2H3ywMBex2ji
H3ltqR9npo3/NQhmjWFG6hmP1Rcapi8FZ6wGJoC4DjNH6GXHpkYEKinSexhq+y7ccSN34gH/6EXx
Ua1+dzFJa2ud1jmTfP8cSeGVbrtB07EK2KKjFyR4X2KdLRRDzhuiH8WRJVM0mKKkK1mYWAO745v3
Y4fesQVloWEroR+MVkeP97bcQsQ7hxpkmVWke5rAF35it1R/903VYxzJ0siL0KS1i9XgYg4HdsSo
M/17zmQJE8WsJ59JhkNB1gTMZ64oIIODe/GQSFSVLc0GR9hlxC1zg57pZJyOCGeRkrrNv6uj94Or
dnymAPuHbPNZfLdD3IqiL1d71kCRMbzYr8EWah0bwETNuLgfQ+lZrFTrZFj+vnXs/y6RLu7r5kfv
BW7X/RQWfoUysK7jCj9G/VRT9iEWaeTtJr4PFI1bAEgbBZ9ldIP3Yq/tNZqgVH4JzLemWHZcwoNy
6iw0noYhVinsQRt84h9t7AtJO0M64I+TGsmxh2xdkW4tdNfXUV/zAE6N120Fyp4DH17hBVqm2nog
+fK3xAUKPWwgWw5SI4vbQmxi3qMqHP8zpKRAZACgKp4QI9Hx6VxHyaFbAsnVb/a31WQlfwPGjXXL
TPXFn/X5RHHqE/+VvOQJ4JU24MrcewrJV9nYVbpoHaFY2+FN9tjx23r+sTjN7aTQcxRX/o46hYEw
mljHItLIx/gC2/39uw313H/CiMdyNEvar00T9tOu6YAeP5ZwA22k2f0s5Y99E75YYOSGRq8iXhMF
DfBoKqu7jDs+vhsNKO2ZNoIqudPYjf2dCuN828u3Vr+dQlf0suQ6ejVqZRlWP7YXHxEH8nJgwT5B
4MYZuyzJ+AmHWclrW252wUPLT3d99GOWePu6G8YEY7Vt4x009ZhNXWIAuVUQwIK3oXjgHM5WXnLa
B1B7Hivmr+qrD9+0sfwyuwCXx8oSVEzgf4Ine4FMzmzrz75OUWLxBWKzdo8en+xtpgfI1wuDd2Vq
OTQ28PfHApqUaUuPnqjc4JiBNnReZpvZeiAS3lQgsJ38+sIoeZnsUCiK6Kz7QvGYtcRKCrwIROsM
iOdxsybt8L87Xaf/YyJtayjSjjLj15DN+IeZMkzO/0z19JDA/YHafM/bpveErwApCp6Agsfj5OH7
j9AUdgvggBIgfsVtSMykE+ZfvZyRyVQ6RGdpeoAtJb6RyUkzIuoZUL7pkbzm2vfFeDJr7zfThZHT
lQRRZmiEVnkV0P4XwdRg7HsNe56s5MctdXZcnpvTCGEn3qdwOCwsQ4Jg16puu8SrYx6dCXbKLDD1
/WXHf+PUtkleRbmqyf1GXIcAfO9JzRSHytk7WpK99jfP1QxiAhT3AexUk0HWrCg5q1RkNYbBKDM8
dUu4cnDH9nS6t+f7L2AFdvDlYlyni1MxB7ljCx1N61o5J4OJakBSVYbnGdO3VCBI9bihcMJkKc/f
F6A5LwXyybp+liDmmoDVK8g6tF6zl8+i9Xm4Y7pA731Vsc7pjcemwTIqgt7ebJZBxhgiI2lRMdC/
1rRYx4XKf+VuRUjehGsz9HPrf5VsdfKW9zECQ2EMMKZdhCm0PjHFjCUoDIcFDLGhjSVyKU3tjTVj
zxrkjgTNJWE3yDyf40LCX3UTnv/6Sk0SzQlrJvwUXDFyjt3EeT5mRqGLKf18uLpVveElGyb2vP07
FJMR+PiuB5GHK9oxFqoZ23QdN4qhbjYQuBP7SbCVLWwwhxO+z6OCa3YaIJZgutmIvfGClondZT0X
7bRF5ZPMpLM5wFJOFG1ENXOAD1mM4MJOvxnaihc6wOLSo7g2iDI6dYVfGInD5vOkAl19P94rfMf1
bPL1pnX19roESOF27rP7srfBxSPkxq6QoL4WnHl2PJrH/i+GXzfICowuRXbB1lg4V0P5NUVL6UKa
Qlr29oXrzkinVvdSQUE3a4iBkE5mg9nrbKeMm6OjtvOELsP01XI422EM7PZZhZlGl2Ka1lUY4Ozk
Owb6pu0Jh0cJnYiAtkAUIq1YVPJa17WyjmQ1///pUaZMMP/1BnbOvoNDaA9WXl5o1fhfwh3wB/RN
6Ypn5h3EmOP5tGpEFnnXZj9j+PHu3eQMcuTRu6tGxHQOBbCp76mIFdBOn/fRRqZSgSvDh6Ef3tBB
Aauww55Uohuqdu8UPUusMArNp+AEnJ6YHMnKzypWeDb7vcwSOLA6XWrSVRCFxAt954trzQsqO9ZN
/r8yaIfK4KvjTzeev6vI9rcs5RHs7T3tkGqEO1tFFiWqNxMbSodqVCKWUrtawWoKPZre2KNl9XEQ
NkU+2lVM7fuzzq2GQnqnPco1ugdPPtzujw/gtsDoCRmmPcjVx7s7u2BqiQxFgJiKCg/vVwwe9gVw
BWRI8OfRB5K2MLuu7U2OAyFZO0+MpVyvby4bCxrSVfhWHw9WCBWNLBFO6CHkqrw0UbVrg9CEma0O
8Pj9vjg2zPfWbyyVSviO5yVpBqze1yh+U4KCXP8yGemrWRBKMDiBQyWRNKxaoujNdBB3lylMaFKE
HSr9wd2aaIH0hm2dp6IjEUpUueX0b/AFGqOkKIorGasBHwpe3+BlWmkPVXllR1nEQ3GxR1VG3b50
54wv5Jtl3lW/tRsKx3DlsX9g/TQSTLs9iCHEZjFV6ywT4x1a25FRzVlntkLUVSlFr6xda42TrAuw
CqmumvvtOIqoFtAv3eXMAzYwXj9fKI9e8HwYF7GuDCCgHMrgc/0guM3oMP9f/a/Xg5tUL6dJQszR
/f6D6zmZkckgr5nmIp9FKrs94epSfwfO6wUtpk2IweiJlux1AlyBZEwo9rOcjjvw7KJGL6GZP6hF
l7IgbV4Q/5VGmy1v8v8nZ5wb0aqiPpRB2ceYp66I5IssomASpZs9QjozK04vCZ6M0woiX7EGuYCK
G3eMqaMJ5qzAQsWyivVSd2tm5soeigWBrU8Y0ZOYip0/Oq7Up5afQspLQEbDfGlnMc/JDS9v9vuk
E5FT+CQWNrOmDic+W8foeVhuIz8YYSn0iKbC8cZpVeM9SnbwT+WMm6jaoh+uX1oG63VINHeoMXpG
2ax7pyQaBfCa8rBWzbATaCAvtgEfCjB0yER/xVnCeaIKwppfYBJkCfI58LhLld39qF16+aV1Z8WG
lNOzK1sUIOYJzMp7VOLGvMfDLFUx5fLedkBNb6tKPX5EJ5LoJK3jxFf7ivmY365BhFFbc/xiXM0z
o5jCW5w/hkiI+qganmlrmAu0HSROcG7fcEdOw5JGVLWbMBpJ+4S3UCnKuUTtENBp8QkFLrTMPRH8
klqgMFLdlCRERIENov2ZT+FDm5eLG2tzhqIpNFr+jMYuTrH5NjO+MDg3auCwTVxj0i6A4WEPaRMV
y4dorTPflmnwsJ9YOH/LvYtyAlP9iVMwwa/UDGKfeYaghGpvTshIwAIl5UmN8l7gjGoSFIgP9M6D
cOtWYd8xLfhici3QMtlmr2+TuULFp/ogyBlUUXD1Yh6x7iLARsJbm6ucPiXGoCshkOfbCOCCX6qJ
Ql4dv1X9dFyjB3nruf3qGTkYm7IMMZ6RTgnX/F1kD/KsFFhRMNMxHSYiFVo6JHROKPC8leLlq4lp
Cx7H8YKM5NbeKiC57GggTQZRGjA7MiJIeTKt9E8YaeC9ByonZrsf9rxTWCurvpEXt2xPnmVWAHLj
3EmenoqL3C+CB33DIha/r3L4y7jpqnQ0cRZwPZzoaGf/9FAZnbKcge3HSEqfZmz5UQENuaMTEr83
DNgUea5vtE3Oizdm+OGaZ8e/sdesdZSQTKWErXJVVj6sjEwBd2owm78NUX7cpg6fu6sqy5pothMc
enl0OFOmUwaZCgwKRNJkP10ooRj9HJBoEdZQgIsmwba6N1llmf8ekk3VB1vQCV7u5H1qMjJHSo9u
p7MAGC86K4anHqUNYAhZUuXq2IcmyhneTUpSsve4hBLuIHUU8gcHHHLSohkS2dRlNhkvgkAoPjtE
baLtvJuaFsIyJ7SYWr96XB0dbKQWC0MG+c1GcPgs5fgWp3tvV01bDjcsbQk6C98IdkX2wwWvKwfD
7Fs07uuawS3wtks9yDiB44onxh47cjOYrqcmjW/IYJKh2O9SOZMYEO5fgYMDeZr0kiFx9iz6Jju+
2PSx+MhWgMJa3VK3EK/xFuP824yVjPkaovGW86NeVVby50OAJZyR32SKPtAMgSgXKRx3ftRlJm7G
gbJBmXEoBvFQj461X6f44gQm3I8gJf25hLv1LdAFi+H9nUA+Gzd2I4GU051xB8m3/x73yBVRE2F5
wJhMdXYFclDpXcSPJxp4tfuqJAg10if6gwxaZWtH8A3JvaR+NgBTg+eusrdTde3wibrBWM2vE1P5
8HVp6mh+CCp2sqgjFtEB3xq5Suapt3xWTGwdfWKTuSwfLorBmS5De9o3uqyxkUZVxuLyoyA4RiMN
J9jh4rHV8L1nDBJZwhodqzj9fNDHwMdOeXYCcvGt5IeaF7MENaD5GkqwMEKeG/PCn4pvmXHv39nt
5GsTsjVlcEDgWliJc6b2npFCb8cfY+yfJ+FZme7nunuez29nruXfJM0VSQHWfUS2JDF0ohY+Buif
55SHXJRS+85UKD4EvXoYQFI8Kw1SRl83pynNdnyYteNAeXZjfPF/RaQryCRKZtG+xdyK1I5rXLvc
URjgZRFNvpNydJnpk6QonPQicPtgGIrxoKH+PNmKvEMXWd9tgag3ABf0Amjq2iTfGuNxw0xUO/wP
uKgkGbq3meI1IBvQx5isbmD5YzHLIwn2EuZtnYI9bndnZWPNT6QiBF3OrMimItYcMaGEiAarpdna
DIDCEY9Ge5KD4jJ/UDgZ7EogdHYXnlKUSIB00jgWDIU/HvVQZ15+LGlQiUCb7RR6SGWPFdkoy0h4
opee7hjEm1PEM4ySP9N2XaeItnsLvlMdtKSQ17wvI+xRd9kRzlq5GUn2jdRLNSj0HBbTtlXGAtyW
uT+PgJOSFRHDs6Ysga5CcRoOAKJD7X64l6doqR0ZKnqkK5rLlvIYIT5k6SkYTCtNJSCJXG0ryC9T
xzcDTcGsZ8YdSpCjD18wiT6VwFIr0DSBurTlIDBSGdCJr7Vh2QPBTDXLmyEGAHys7VHe76Fj+XGV
bmy1PJZJrFD0Z2ZWsbqUWhDtt/ISpawNCM1Dr+tn5wbBhuVy7kxwaX1z/d8Krmhgp4M0EhXblU7m
rURCLG/+XsP+0KLK4n56T9D7fEPqss2BsBJhb7wrxOpev6u1EE3jRAsURaxuZtB+eiCrpuDc7D/w
ST79kWBwdQ22pVH02llRfQ3gquwgGkIP3wPSlTri1fkIl8GBEtVpQZ7NHDT1b6rjK/l7QffSplRT
ccuqMCqCiCFS7z8EQKi8T+nlK3Uy9RP6lOC9MIRjJM0ZPLJjCUsd1oKHM9+SYY8IEZplhTpwwEdl
7agvU1vmdPTN6OxS/YHL6zSlb8Tf+qzCdA3BCn1K0h0PrCCnXBopZnGX06sSiBb3keOdxfNXlVkj
2wjj+RJhkBmFLTXvtgxOC/qbU/qVVKzJUI7ywGEJQNiaUwaoCqZlfRpHHIYBhP4SnGlYw/NNLYYu
CIe1yOwriNb9pd5YjMU+GZtmg74LxVd8NRWGMKjCwr4U97dfTlQ+rJPnn+/EDchaLXOvbDVS1nYm
WU7GH0QRKndssveTgltRAIV10kDsVpBF5WOR49zCp+M/fufMUxBjtJstRxSCwQ8sEtDsRdQZrEak
jULbd5IRoe4IE5pwBQNX2n1DESY58Pg4lZBMmBWf9rqjs+3kTEolLveVulXgXQ9pZJjLB7bSCfSj
SdjmXby9M4opthW7g5LvsoYLQd/nTLxQ7RZDS0fziXOQv2Kehx69p9Gs9RdX5X1Pu4xYgUduc1aP
0Ssu1mfUoYjvC+iOZubwWtxm+EDxYnloO77jAA0A63895rWTsxF/QsCua/4ya2WGUtLCYeJesZZ9
cHHkRIQaU1UZb3P5fC++oYmSiJ9UWYeE4pjq7mPHpXdbLbGEi2HHT/Ah4Imqpnv+JCdLRDHxBe1c
se9Y2W0ZLBeFggqD9JFJyqOssMJn+ywRDcFXn3bPPJc8yKyaa5euq5UVqBwNvwnJlfRIoBCJ7g19
90K/11F8VAJP1XnyNXGvZ7kGtVYJPkME4hYrw1TBo8MyLXvZaxR4Wz/mL47rl/8gBo+z1CNbvzcg
YevwDSuyGoqT4tmRD9QNss10Bly+lPlI4bh76e1BmV2nAnBXjf9HcTUniXJgvPaR5mEI3wN8WTzl
+uRhWW4J6gUekfR0oLfT4TIgq28m9PVUgPiLiwMnzJ06300/qGvB/7+BPjr1MxLtfWaNPrG3rTCH
0OnB8kP7LgOJ4KTgYRI+ZaMt/DoTGgLU2qz/U25wk1x6p0Kymj0Oblc9gscaETdreNmoNJyu7wBQ
6a1j6lVvy3woEAUp0uQ+i+bf8OpzhYAcDNqsT/ulPF3L/PWKcK6YGX6cmHFJRqau4kr3GC8kFH3b
RgDMaRQJ1HS7egY3RllRFxWsaEQxh2YTu2GUq+nZfZcd0hgykd8jrDHDcJ/dIrMxHDcDIQYmpN4D
2r1X34nxn0uR4TINJkA+RrH5aV3tcMBS7QcxkDAfU3MuWVJ+rjIVD1ZDoCmdqhP3Vd+Wnn3UOaXC
2bDTNExYlrM/bzIsRI5DmoZIXNno4YDWBcuQZt+kIGAY8uZW4shNMrSJJktX/qymA50sJo/tPqil
QVIisKoPqFeLZv19FVEy55ACTdLqnnFixTJIHeVVRDZqzxNGO0Lel+TG94mqOvyxH2hOE4qf3K5O
Oukx1Cfb/WQ/7FtjHMWV/DUIP1yqOpXjBZAj5tAai8wbEriV9gJ17K9C2+tBLPkBGIPCWGfeA+qK
tucqdZhpBRBjIuvN7VAMdV24oT5OfYYp+IBxbHKwbrK9nJLd0OwFXC+Yb1EqnLkoYn0BGm6VLl5o
btQmxPvGmJL061QKySKpyIC3Y6aK/6C+k5uozL34oiWMd37EAdQ9WzzVzNP1rBTDdFL2ucKSOVpU
0x0+0HzaXopsgF6ItyI74PI37ljflEJNOukkh6dAH+/K27StVBAkvfNavrPT6+VNb1poMMdR9Yst
K2QpQ62ht+S4So1nQ5/pCVMOGznjmDxYoP1jDFTCr4D0UbgaZP8ZTLX7nYhc4t0/Fph8OP3mQpbV
3rG7DTfbfuWtrABYbS3KM26WGTQolBKAb5kSlkM6ThFgxeENFgmvjXpe/3iHRgvHUKyo8VqzPIKU
XTiAlZKu3vtCzXYpOiiu3fmXI4LZJ2U9A4+R/Q6hGUAJHHLhBbvxtJwzpG7K7WY6PtQ+8wPFAP4w
U3epUFUjKU9zqQ6/Whv/DxHzY/kLcmArg8lqvihZvLQatymCk/47NdgkGfZ5zdlRxjZHeT0c91AE
V85mtzocAT9ZPGenyyUaxfNmay1g21pLDu2qSTXLNwc/yhYuddohSZwz9x65LSdVRKpq0F6sqGxU
rET/Lgp0ulRBcjyFOZcUF3Ai6RaJzF8DpFsboqMej+monEN7dH7NPADkcRyFpKsYb9BBA8Dazj+4
q3W2IkDAlYJ6/tTo9D7PZQGomlHTelgqXueF7UC36cfz/xDxlO7OaTtt3z7LLG5kTBuTHTsNwmQu
bWjz+pcBMlIGB9w02+VGFVmI4y8XY7ZaJ5Tm9JjusIHmdYMoJ8U51jKfIRgm0eEqt/kgJ6lrKVIf
kM5N4wOGfd7fyFbS9RlbQJBBFgx2CBy1vyPDp1hLfGpZ0A2moyB+fnitjvOtgSu8+0Ngzgu+60IQ
5U35JhfcaLMksy9liE4r5jFduMiTgSdLHwmZO+7URtFb+vnDizvTq2vZ5IsxA/h9mc6Lc62v4tT2
qR4ugddtdP/nNXx/E5hNNLE66oOclTyU2AtKsg7Hxupqu30M8/aGbMRTjcuF3eh4H7GRmSPVw7kw
nB8hg0h4vA5tOAJ+jHGVMZ7CN5rohK2o+5pn4dhrRsrsQYQK06doEtsOfi+xMnp48yVt36X8At3C
uhpYZPHRG+N3s64fJckvVGScDPPmqRsVX1O3VohS5kud3ZVWF7540ehehC+Ku83Iq2l57wNiY/Fy
Qfj3WjVZtPTGLA1eBlIKh9qyrxEE8pkshTtTJ6nRC+L5zagclqDXTJe8v78m2XsqiTpGIQxVGLLd
GkKTiiyfxVSl2Xf+6hHtpbF4OL9zsV319FAOUQsPg+AurRpnf8D9Adyu5XOBv7bbC3lQBfFAsau7
vNLy3aHmYySA9kbSu5ExZIABxS2lRb2e7aFk22JS3DVouzpMif5Dh1YtzeEBXyanzeS3IDxl0PBn
UHZQt6lj/tyFUd/kNEP8/uC35lgKBe5KzZqffNuv9ZDOOiIXa+8hxb/0jKSTG351/Cuxux87hQuJ
QC2up1NK7KDt4b6y8vDw3+NdEZ0Xbjl7w9arXhljy6CunsU2ZfrZZQbcYxdTSnKvIUjLtIO2o77D
sZZLfqsCtSy8oZFD2R5cDNKWQeTQEMM3oPFz22nMf7jZYE/tczAlqqUJrL46TTjLIo38VprLjOc2
g2xOAMFYHrU5L765Z6FJv62e5RbPZyCpQbyrN64F18A6vwgEOjTRxaMUB008/TTwPQCTZKHtUKKY
9KI3THToE1eGVLINbZjmUjZZ2H3IgfrgbhQIfPFaXVo6dJmwgiiiUNM0ri/1lXMadak8SmxJUybN
g7QTnpa2kdxrdIjVm+TlzjFSz4POkg33LqyS2Zk3sUAgL3EYhcQ4J5v8t79z2SVkV3Wk5kjxFoBf
0tpTAzIPhG+NEnOZJvv58FHUzoBCe28aCU+Lb/4kyxWVBAvZ8uUEIz5NIb8970FXMN/DSvo4kVro
oFB1HyoxEFYtrgsJ7wwakKvHHeE0pRjyKJJVxpgOkHgWa2lfYje2Jfs129i3ZwOxaAfkMNg46S1c
Yl9F89QUBowI25dQSkdPNeanchQadEs0As8qUBLxk/FDCW9V7XL3Hbh4JB6sGyz2GqSXp9p1pqlf
zyMVdLf81b1gVBZ1zGu/1KwCULSEk3TzBmSuRWBviHXtDwcVJOMPKHQlGWyB95DF0ifXKu5ClMr5
SLwisqHsSvYVRCc+X+1mnLdg47ZBqltpIOY3+RHZ1ckOc3iLK6Bk2bJwEjXSuFhI6qE0XkUDjZjG
liwZxS5NuViv7TBEH2oOLfQ58H1icgRkiNgby2IpqpUkHjjQgfk4IrxwdrCMSU6tfkl/RXlkb+WX
WGzunfICuoUq8sck50Uvr2msv7jQO2Zjy5YazF+8edTKcHmYmbesi093JWuR925VwuUvJLm7m4eK
SpytNyNIJwTkV0aA4Z676wD/bfZerPFAOaVEtRykJ4w1gL0BTnVdszQpV1ZSjd5ucLX1VLa7ClY3
X/7+lGidKuZqbIsIe+owxWhMypaFjj2zlpJ4NkXfh9YrIq885oQxCFeL0WoFHc0whvvOVXHsPbLa
CJZ0L2hnff86zsVkV59tb9EfRBGZzPF6MS0oui/aaTW0DmLMmJB3WRU8pEj0zqo2W+BLP5BgSfOV
/3vHfA9qhPvWRTYXKMSZ9+ELXUuvpbCPHCAv2tj59B0sZ+W3aiLooYcFPxue2QT8zaS6NVWRXaBp
eRfBb9YRoI6PEMHYIc8ptv9XzcgWKRfh7oIEm7eYWl0Sb/2jcutGOIKelN1by9x3kCwxwZA8H4rl
EktotgDJ5vpyGapssFZKrIYCIl1T4WcPOHcVy2V7ZflKzNIndG54RKxXet6A3yws14hzSg57q05T
TjEwTcDwHpw0tRldPDyA7fJOb7WMRACTMpxQ5m47ST81J0LhHLnuudvF0hGWzKh7YJfOfeSsUclo
jkiymRLs2KYZXiT5cQPanMn3Funydp9zNgNGCm/qxV0nh4e4c4tQvFw59Xp9DJ3XWeWTLqHaF/jd
tQcu0B6+Mp7eojqxSLC6xLL3P/UoNsqaUIxECHVsTpe1pau6nqJ3E47tXtgcsvd4Tu7kzqxTSEcU
TvMBbSW/pMXnscLYhcl6Q4D5HpTBLLzPquu3UTim5hXwygnqDLu4gU/keOBAjJN0Q69S/fH6TzPf
sTrKHavz9MhNMt0c9NVBPgMXLENqec/k88Rrm4FUTrW2Y0J07alnaBW8aTM+JzJY4hJQ7jxgbNwl
cymK8FXDE9Rljg0rD6bmZe+sPLNduqCibSJLW2k2MOyEGGfJI9841XkF++S+sMJUR4rXpMl//Pa9
9aZyfWA7zSg1Gd+JQV+llEpScyXpH/viMcBFswTO6Gb9Knzs/0ff3cC6Gc3DJVhortGXzsPzjCu7
NSH2vpmRKAcNsAGBYpinF50RH3o5jn8l0Rkc40mTcilZLh1PvJ+XJ+3dascr2kKX9WPICZMfe4QM
BWLo5gj/tcKgjeskQdVlzzZ45+ZusgBV4ia2l9KV1JtWh1JAP1zN4p+NUiqdvMXN/DGwq/87cn5U
q7dUZ8EpBx7gHndq4cvDQ+xFN1EUQstxEZU3JdL34+ELOSXHqRJqYGDfly9bo11QdlgJbbiO3rfP
1BzfWrnm3WYpsEUPTlkDzHbI/s96bTcxKv6gooOrn2GWwXK3JqkKXPGoy+OJ6pRicicfZxFM1Fd+
3SD5m/DCo3vEn1jqnNgb5Wxz73Es3eOjtC7na+tdkYSKoWmbhZ0Z+9nQatxe9l4E76o9Z60lAnis
q5MqTlDySiit5Sc49SesIouXgniSpPhHbaZ0g/jGyvh70p0r7boUO3XIV+gpZrV7xujHA02RlS9q
6OqUENrvA5rS85OhXDgeg64obKxH7pDiwzIYY5DVLe0Zpmli62xEycD5AvaClJbN077tFC997ewu
Bn9giacCjAuQ2wydLZa1IgWtbiE+TLE/Ic7adDgE57wwHuN/vaw+ROWJqLUJUM/SRNZ9cqGalmPV
+SxLLeBPS1eugaNFWpYUS3owp+U1wsJ6GSlPhhBPLtJ5pGT/n5ZK1CPhtMkFyAK2YbmhVFuc9fgo
pV6srrzOZO43ZvuYbAHcF9eOWj2JlzlwzQYvyC9S6jbV80IQX1O39slYzw4he1TBgiQSf/ZFREgT
0P6bOkDuEaGpvw0+yWRU0+o4sqaFiLz0EERZfaZhM61RiPkHk9G2lxe7zQ+enDSDVf0icfdQIwoA
fNfTwmnjrbgowGIWlsqLlXnvPT43M/OnlC9WwqgbRpDYX+dms5A3UdWs3j1u+eUQ9ovL33iZKaMY
KHXcnwLR96NfzMyyuVwdTuJt63oBifLlcaUYPdHFYlVfR/yUE2oNwv8o5K5Wsjf5WlJzf0jwAR7W
VTSHX1NbzpLD1lU/wxbBfcVGITw06STabZkuL94o4jnL3WUiwhKKR/hTdrSi8q/8AZson8o6f/OP
QS6BlRLp+tXjXBGltP230MWWbZGo9NIqpWc4oliZvQTsQuo3d/i3yPZnKEkTL1TqwjuLCxbLWZJH
V49iuFHZOhye4hxvpCK6+gPZvfw3acqKeNoCH5MkpK7IEy0zw4uNFs14rdaQ04gBYXL8+pR9vlOI
rEbsr6kwp1zOtcyz+IR+HLnYQkNWQQQS+K/jUFcW4QzYQgcZ7SJPjxqcY4gdzysMZYRMSJaA0kxV
zfNGAmI8XY0ncyLTEqmRb7PdXCmCiRUFzazFNQmz0RvyFoI8rpkVEsH+QqpHtoAGuFFnzBGhKQ/I
O/zaUZft1qXOl4QBnDbH3H/VHOGhGDwfDF4Qf7j/OqPH9bSWTz+YfyyzBrO9wTvu5DNUzwVrzEbn
Sp/Bt6DtWJg80t93cUg4295kejdyFuxo+4zziJr3kPTCjp6FSnNnxLJ0e2YPTHLE0GXCrFTd+BRk
kdYz4DmWGfhKRQkEy4et/VXcg8Joiab1IvDA+byRLiRw8PK/sIQY4GA3kYycX40kKGcRtEgimNEv
xlATXqb9sMHmKfXDg8t3FuISsNlAfSwxymIF0/bP3hCZIyoLGIWNk9lRJRApWtM8LfGkDWYpjQfw
HGuxuYSY05pzUk5o0gDrkjYEkBUgNe+/ZD4mVKqjgXbmyUXqxozFiE7y5a0NKsiAA0poOFfe0dvz
dsAGg0rLcy68sqFt5U2mI4zCmgzz6vWT4GBJ1Bg1mZRMUCWve+wLYrK5wT047KCXGOI9DKFBN0ph
hMq5mSyJxksOx5E54aw0jHPmsxu6dhwbdvfbuYHohX0fNgpMeOEbAj3XOXEONTzkg/QlKWw/OWgx
MJ4UDu594sKqPHE5xGYxk5WqhFjyVozxqYuOL6P+MF2Xfn0CQ8TNeYhLDOwE7SY4HWFV37gijMJ0
PiDlou4n1ABrkftYwm6RI+SCKH2oBmRGoTloTF6Tdbnifsry3rDr59hN5KQvgadrbJdgew88xErF
OzX8vdi1PUaE1EYRdiwd6H0/tAHf6b+QJooBC1A/Y1Ldk7cEZL225qAmqqm3UyC27vm4/fq7sGiH
HwadkIo/qqRluZtXIKGTK84CP3dm9NrVpVEgheiN084Ac8fOz2MvnZL5OIdSscItQ5i0F7hH0D5a
k4eA/Lcsg8sLp5A1HoKR1B2VB9T1wCbIZyTH0ycwk6b9Omcrv8UyAn8zmIpbs9T78PO8WFvnujuT
kOh1DGmHkov0JVP+8GN8PTbSP+iY7+uUoGHJqL4yEMey5/52q99KAJw0ns08dv4c8bOO5biP+Hsd
bKSi6ffkqs8sENGMmLENej5i9TEEqfj8Ua7xG0M/K+/Kv1u85Niya0KjGKhYl2Trzppw0Zx8Y+/8
y128tc4MWeweDNh18q9gcPL93owVISdxndXm0jIgjbdDyqVNOA7wXCyH7CPdl/EaXPe0LvQjdxtg
r7x4PrSDY8XWR3Gz8NlmtDvN8pweZgvGy7SGMPSqjn2bUbQgacWUZ3fz7cybXgMlyY5AyBs1eU56
p7PLLG4/XEgSxCtZCfRuDagx6gnPE8NPrT8EXmk8zeywtJ7jLhwixsU8ImTmKbVRZzRnVSC6F9Pw
TnFNF8bUUJKJtLm/88uLlOYW0XLEZ9cziTSE/ZkO2w8iK+8A3zu4CnV2pMn8QMN0aoR8yO/sfip9
VjXEW1dyDH4qbIRPTgE+ws7tdabnPVK0pddiz2IlwLWh7TV+vE1EJZANg5fY4KEDpBZ+1830Mder
j3Qt/OFuq+a7FjOP9aVW0IaRRGWD191AIvHTG+S8P/C+y/gM1nSv5Cuk2G+PkbXZIlMYquBxVK7c
ox1Rowq0Wwr0kS8Ov8ab3JB9ysI9kx/TQRlIF3XlQRnHnat8YUVv2cPX2635vla9LQN5FD+UKH4S
ezhFdIUAeYqgvwCIJ28uv/ToZcAmU6IVhh44OiIj4FKW4evOzv3kEeQ5AOoxlhz0xcgSeYcJ9+R4
JdirHd4ju3gyBGOvdBtn8Bk+rSa2HWSX0tiQRZWSc028w5MfWMuxm2W5HuJkan/NfT0t5CRpgTTR
Fdp8HOURe0muOwjmDx506IN7mIs/z8IXIozzo1pv2osHGikTCU4PI2Vi4+e8HyG+cP11QUgOHk2c
KwQJPoD8hiu9mjO6+7SwwMH+1w4+2ABTiodAfEUFVeDADKj5o085jSEaF5DyFoEqO4VNSBDxtTcA
WCSFTSKG/ryF5dJW036AT7Q0ueTyj5JD1AHdevvzTkc88E/ocJOSeBTjvkfQui5uyJ2IE86dlFkE
esV8uoAAD6GfYqWo6Pofoa/AM2uDYTzDgF4G2Dc1WLPbir6vjR9CeQD4aeauzKFEIBgCPJX6Exzp
jep+n1h94Bhz55M/G6jni1WBmBb63tneqjYtDpw2WRopAlVDJdMWMwsu8WIYvjIQ46Wx0focY/pK
bCrsHi96AYhYhSeTlAvJQ/MVjZ/yJssmklYeXOKlhxwn5SKWQ9Slpu1olypbVBj5RhP0ikRHF40c
2fxDtFD98JJX5ec0up/uXVicw43x1GXMpNvM+806q4Eh3S7LdjxVSJu0d9NB22AyDZveydelDHRc
2D4p8LQMBan7mv+padDtaubCCFJI999YFFd5pBkkRUvHtv+oyqbcfYbLJVY92oRf+byONk/874B1
L5rhdtwgVfeCsl3jK4SqY3I+tJ1F3kM6f3ty1vr2pDL9aUcY1XcNAiOcwMFI6RR2iOOqDxW6LJZ4
XGlMN4k3Q5wu4hhj9w9xIAaEtuKU4f98xyCT6CSPbM0laMGwWpmvDSWFc0OGoJyfisb4kT2MOf3N
hJxkUiP/l4ZuArvY7cPkGwl1AlC+zLdEwDpytODoRcKrzi2CpEBdsLrFzyn7Z9E8mhxkrAhMmqKK
sNwgUYC0hwGK1bHJhO6pwMdWv7lV6PvlVlv3g49OztRBd4TnAKLc51Mm/kTIyxOtVbwkGMH1GvlP
EtusenYaLB0GRRa3VTpyEJAvuSi59ESf6Z8tkD7Z7s6fymiMsA+6MQfIm03Za+2+12H22AiIMpwx
VgysdV1TYoub0olMXbfhk8xpjt4p7588FYbDZm29S80iJgczAzQY1LYiv6mqlD+NIbp+QTq+R1Mi
zPNvAtDk0uvyF2B5v58XjnemcVGgNKc0qgHDO8aGDgelId4de/FH6u6HBVzemcxYqjb7R+48SGOy
pMBwstq5RGToLLx/DPNaqJxZ88rgci+MVEXi3KQzx9AgwmaQrVgurFkI9BZ221nU/LesQ27AOGYl
CoLalLn28TC+HSVetapWca8q53KytMLHtivj9ExmFtVk6lTmo7i1gJTCKMEPFo785uRTlvAap1v8
BW4xj3q84WojkAV3+6vui0mKpMU+x0MPG5SWd7fbjAw0JMCsSypL4GTrfox4I1m965grXcsxgJU2
wnoFPsbWKndrdd8/M3E9Ul2TJt4m5PK5SigAhukg9dLlK3nXv/qYGCQhKWnDr0KGVnnRyfhDCbqw
yFbnyI/f6k1p3uQH7uGMyfua6Z/ccvyPkYmZKwz4+29IjJgvHbzS03aKUwTZeh7tB45hObTpR6G9
d0BgHQ1tbAjiaTNrez20KFffyJmW/p96JsX9XIxJNsOKZDJfszOGXC0xTvT/P70C7b9Godowbyxo
15Dg/QQe5nd3UHNiWf+oOrPbYcGKuGozq72CToHLSgvkgtOXYkdTlVyRhTBhQ7/CRPOHUzG1aGoE
/rcnJYKFHkGBRnfr9pez6F9l7WuwTPbr2Yj15iKzZnqRlbsPeJ54VNATomAr7UBy/o+HankkNTA8
2KDI7ltWQqYIuKpoauNz5ZTSKJaJxU3dKa3MKpR64iaYsnOKAE5+13grv3LMoa/ucFW1LsK2I1qt
QMcfg9MLW5PsYlic2Pr6yu3YZ+UcgP05u9c6sW8Z4xRek3WQd2fD0+/12qgR9Y/Q/UOdFVzh0aTt
svCPMkzseriehnJ4msmO9C8rcLESj1Z0EQ01UZut5qIXnX3+Co1u5wbTZzxBLmjFYqbpTdBGWmud
//cd+FTSI/gjzVA6sf46Zb3MBFLLj9vIVI000Pbcxc1blBWnbqwFBj8GOt8DJGRP30vLvxTCcKtQ
pot5Z4uKNvQ9U/6+1MjVzJzr+Kh57dUuVoPvNwdca1mgSY2pxN1TYfpMfK1w4tG1r6s+WhY61nT2
OhzNkAkO9fnBlD2LJ5mrEDQ2QQquyhXBQCQrLu2YE5yI4TpoDAejFH7zbgKYHfJbGm7lvSrveUbs
uO3yBKxymwr6kHTQG/fKZ412loKgzGdMa08Zo6/Z28a9Cd/C3Bbf3FKmyP//JIBNRgVi7RftwdR0
yzxLg30mQ6V3eJaGoqULAo5znO5W932+/2bFObU5RiSiuhz9sS+BnDima5J0uOcLBihJKLKAItna
vdnVDUCxw8hJSKJl8eXaGoeNIZiKcX5fBTxlcq5qU641Yu0xWR9I3QlsUKX1EDKZ6dN/XzhwsKUc
Ui8Kk21Nhs3bWDJh34ajhzSwbKyF+SW5Xj6tNsiqzt7RafI19HYfG8IQOyflY+pt5ht/GrZzyqcj
GQxwQhLwFyZml1rjhdWrQznbH61IEnrd9C5RsoGJERRkLRvLw0De83NRO7ZVyFzljhBtGFPhqj/J
TNF/hv3HWOEK0QiNdnlDhxY8HRcfRLNSrXmblJBak9T4JLjV8+OzU1KLSxssGq8Q83A9cn0aGERN
hT9CfKs4l32bCDUXDC8TaCCpm1JoMEaITgX7pTO3fNzdyYLMEdDDrkuVE9MfNaqZwPfz1SDRoEwv
tUc6HH93kYygIyMVCvPMelVsV6xpZurWy1CDb9ASNZxMJxla+vjw4HtF052mfMPL/7r80hKgdu9H
jV0u16pWCUWSAjKYvRkEIQhwVClmSoLGqH54aOGzMyCE3XFGxXJ0TxTc9DSSQbccwYqpRdFFpoEd
hLNm8Cu8xnMacoI2hCfOSBzw8QoxK6Wwo5hYIF7RyvqynrAkY7Pz0GVeIqvvYZ1UQVdok4nFG7C4
fvlRkd84StYjaEvaYAz9DqIGCd3fcSCCmoIbAYwxwY2VoDdTjM5me6O1eyEhVxR6ptmjkk1ztbJj
FZWZlXsGPPgNnRtzVyKnHgI2/sCEeQS0srREky8ymqg0s+Fn1ZH5YZsQjdNf1Ia+VwUD2veJRHRq
pgxB88eRhIII8/iSlJ3iQRxbpXAmTnSOJdHcsot1mglGibvhpFSqvHkUgYrhoP5WYzyMvGGPgeGL
CxcRGLVcrZJaMfzlctdXZDtNa8xgaXRTqPJLThKGbGJxL8WtO3JpQA9DKEIJ/ioTTTZf2cdX4LcQ
KRUXCtD3mp/BY4rc9SbWkMtMTUpA5NTl9vct0VMQDXOm/pNlLDECsUvQ1OoRCRhcaH2cZf2fNJ8/
ulmde+vSturPpZ4Tz4iEo/GmkJF0JyskJPVoRceCpJ660NGi7wElmWK3PJWrXlECkxbhyyDyaNZX
PUluyCJcz9H8L0FQwTEyC/qUaGZky7FKdUzDynpIzA4/DWb4m5pEDF/dYriROdaeRUzObPPwXcNS
9VLUnq9RnpLQzTNGxQZBzPwhVgpIChAVZW0r0op1Uc2u5nxevePdBKIRml44nV9C089LGk5ECbtg
t2oiFIf7DUCqGqGbNL68JyxSoae5VIBXqZwq+OLTbZfOqF/CIo+XrPLa6cKFC1OgFkNpFUfxm3Sr
VJdmKRTeQaq4gFOPNhgrgzBrCIsnq3IYbJ3F1wp72xtV5FqDbOCYMKF/qh0gnh3FN/cvOvl8hZJf
O69RfkebCG/Olzn6/GPyErttCYWxFLacFhfCAz2SqE2VhUKfe6IUWCgX92ZljlUQCvSWQWlDKmN1
1saPrhQKrJff/xtp9pRXts9Qkfa+7IcovNCedhzHzuZjhGRw4ODFfxKk4SfCCU+1hQypLuLJy9y6
diCNsLhaRerVcWjPrlzIt803iaMeZf2YlNzu9EjOuVPXE240MHa5dxLpQ6wU1EvFtp5MdlOr8Ucg
NzteW9YqFiQJf0Xa1nRu8YNJz/PLMatGVkMlFaybbVYORMxZD9UAkOKLgQdDeAjzbn30hLeW2nrf
q3NrzUyK5n/SRiLsjxuIZP3CpBShQXlJSoQhueeO2BOxPhhlqrd78L3KikFHy22qRoa4S35yq/n0
NrebUAzhr2rSNKY1S6Cdq6mfdB2LuNPjDM/YdhcCMbHXR+/owiYcatdf3NTNDDkm9/xEGNNm0iz3
mQ0zc1By1v5YnYaZnUlBCo6ke7v/apjrrn9yTYpW/IO5L5IW4CsRGcORYP/LJCw+SGZcIXfk0iLn
Un60DInkjn6BJx9Rvzb/BqWv39ImCtETB+waKSVVxS9mCerFQ/4o/8DgvyPB8lMAlXsYhm3h8Lzu
ZY7RBuxySaZ/6pUJCeX2Fm3KM8+54CSxjtlZkpjetOYuJUZtX9pLzepkSadQm7/VgRcOT6B1ixrk
oni38WTo3pch//D29NHHA+tVb6tkr/+3PpsEYGxefmMK3Qj5E98PulGD2ylKjUKPilDTUhTqsAwJ
h1sQkdph1pt5DtwVFx+PgxEERTn3S/qNuhSrySIDdPKoOPyzdgrtwlNRtsEw16x4hziKkWwLyOeE
aa07cHml8ZNU2Q2JiI51lw1CRsk31yVZ9SFF87CwAHq6rIy8+LeeXIOg67GHU0mMu0sECxx98+UO
3eVhScrfVnfG1DQrYqfaM8jiBjj60Mu1OR1ClM3DDSAvYp45QKCym9xCx7b3fOnh9A5J+QLN0gCO
sLQ0mNhXOcRVMAY8Kp/hwLGDGAlVjaobqt8djPSMlVXfav9eySeu8i8SpmTkhIkcobq9QygmzODT
ypWGfCktExojQooNv78NbhJo1I/koHk1sRpnpaGDj2KbE6ur3liNj2qOJUO0lfLKlSwWsWEZUe5u
UXLN0XcMB469t/npZOzKrX1zYRRjQJOmNPaotoanF98BuPwfIwXqYCzusB/Gpg9QdeEc55zJUYCn
42u36bxDEtZIHFsStCrMnD6ehxn9nb+uw6TPCgmE4SyJDsjvywrV3Kp2Ua2c2oHBbF4KjW7Kc67X
VOSslAK5Y5CD6gHj2Q7t1jwrWnZFZz5Lg4TdBi4zslGx/ByZexH5OVLkPsvRdALKO+7OOERYCpf3
f6gtmRk8O7lQMnj9APSKxto4/etNhHtHWn6Ld7YAZ0hIZFmKO9FcfBDN0xR+ciGWhpQjVpc9U4qW
dvgnSgYce963fLABTfcJ8DaHJoUFZ0LezfMNUJUCMsWwPU1y8cDbwff2Kh3olyazP+b8NUJewQ88
NXWv3JYMMpAXoEroK65UWjUVPVu7prprMq3VGULOLdDM3XccIjUD77t2l9HalGTv9u0Nn1PruF8e
xpHveh8Toj8mqMfqgxXSL3efbH7yppgIE2rQV0grmbIOrPCKr7nuGOtf6wevOw5Bc/xap3JjPXle
kAILqak0GwOueW3K0Iuw/JScImSL8/p2dfrbkSfCCnQtgNOnvzPxATZdfDxfTVQ0EegzEsxKVVF6
OquPizQmOgWCck9fsFgL3aZNeOFKduXLNl10VwOjc5L7RAJd7yZCqU0vtJ8pFLTesCY8n6ub4Zmx
/R19lRaoTT/NO8ugTgYkl5P0u9dL6vnNbKYcRCPX9DyZ6u0s8RUJnaQ6uTBm+E1fvbv7mghVaC9m
Y2LXRl1R0au9GpLTfALDdwmuT1kOJg/98kXnY1dkn7+upxjWPKgDxcjmMhhjdjj0x8nUfA88U+sM
JL6ZQUZlJt0UlyJAlXKX5O7oCbm7ud9kVAtfyKbglWFDNlanARQnUt7h7WbSj/HEDjOkK8OgpqNI
f4t+3C7kVpYFN0zRVZJJkubnpUEGv4Z91ZkWGem+9aHwmgO2SQh0yzIKQk5S6Q/5kwIX7KjtnKBN
iyBpowvASn2ng2z0MMByDQJ83V9p5ZTSJxYHMDdWfg0go1xi17FPx/OabWqdQev4i1CrLPO2fZnf
B3WaN7QiGiR9hiIH6mUdV0ccs2qTicfNsWY0emd/5s7qoCzw+czVjYjfoXvyON1PB7bwQhUaVEkL
sh2l9aAlywS9BfmuWDfNA3iWgXAECpB9h2C+y28vvVaIqJVfbDDWDlVPDfStUz9oMmK4o6M1mdTM
Kl8nyIq0qzbdsMTkMxWsIFsMUMWzap0j0jZtgVdxIwdwO/7GHTFi6oWcJ+otEpd074MX01jabr2h
IlVY8kGvu0lLnsyHswYkDFGBs0afdAna1mB0OsSeNTQRB/QmRFuOsrGIpXFRxOF1Y1gxi81msyGv
7y/gVbVy34w8wK8W3m/k1+TxXA0TnQQDzkeBL2VpqYc5Hc0vpUffY/ZOyZeTPg+DFlAG+iNeO6CO
QJrBr8cDcwuosj5Yw9i4+8jzjnvXJXhZWTltQdLGeBLQFt+92jcs91RKg/KTxAZnyo9kAJieza1y
YWSriNcAHG4Pa8EUbrkZrN1pvfETnvXbB+1aAyEHgZB5nOQDQBM4iN/N5BhdKYXhk6U1FJYDYuLL
HWQOjbgTQLPgBDCiF98rPD6pzLKI0VYTzRFlzse7Rez3OMzZnUkem7ZPwupNBBoHxpQuuQ9sIZfk
GCxb0vTlFK5LrbRS6FNZpUijcYQSiZXf4ren0AFdY2NQDeYqemg2gyBfK3dJRsWwlsP0ZVXpTGSP
bLcwLEIOSsWzxdHzIzU8oEesFOHi9RLv77oTC6x5DafjZvKmVtL0UVtZJRUbjxyYdhclhGDQHGaC
EHSAXLtLBtyBhUv0SCqLJyvcwxg1pZJ6tp7tJMnPVO0T0GCb+JMuVvqccmDCXSlTYQDgMgTPk6up
ovXX9jpCmMpeS6SimrOcKP9dDGk8WohcNk0a52uAexZT6XXTXprb7nwEY+eMqvaU5ZRJOyl3Jxdt
aitUn7jOpYUV7FQMkqkPm+UW9KFB1rqophcsVatF+FpAP+thLsWZWWpddh1m9n1nNady7+dK7QQY
CBRLW1mnMS1cCMX5wMqqbvMH/FUon1uEQmLdvAQh8d2t2wQGROIx8N0dJOrgFbM3sl2Wq3pFVL06
RAJ8gK72SqazYXxXoe4SkXtJiIb54Zh1U8OGgVdwSZHLYXT31dltVdF6yJNvb/tAayaSzG2Ch3wW
FyMyOeLmJXLS+jyBG7i/KkdiFnBIFEVxPas96PiNVgqL6T4W249zncRwEQXvQTxn8DBhWwP8VtO3
AZfhsLD70pOgmzlE4Uws45J5miRnRMIldCDZ7M8Ma4AC8MpgPlndQflbyYW37U0ZYPPqhoN60m7h
t6fZ+LU7EhA1toehIdzIeaZ8D8BpqSpVfB/964EaAKwBH73Oo7rCF8b/fU+mKpcjJ3/CS8TI3e0C
WSdP80rzTiNjhv5Pmb1EVqNsiCJ6fQuvOdGs1qunNIWvR38m50qbbExD9HPzCCafkVnFdiZobYr7
Bw9MUiAolJ7XnghuhO8C+zqPPTOYN8N1EZ8Rt5wxjnEmXm0oTx4/rewq/mLVK3qqVdBa03kMRuwb
ZyFPghrGulEv4v+Z5iLze2YNWd4c2E2y8BaFw9pjonMxK9z9u0g351Z81+Tt6M7BqlJ5mRKd9eP1
2Fixxhx+FLPY2A1D7Gpg+JcItMzpuUAuwa2MM5AcI1bvC3H6AIThKw7r3YTXxyz3maXqCum3Fn67
IdJ7F9VDLbtjqm1vFhrbYceqbWTBArkiw+avr5k+r4qjWOYoNiODZmfWso16iEbJHM81oDIEm32t
Sz7d5u6COz0y9sZGr804Vp9B0cXSqWzRd6QMyrQJvxcKsDg9IBRljnLn1ia8qZiPoeTOHl7p+Yhf
wojWJmriXmMm3ZuUOmwjH26MQAWWA1fW4EvtcdTsRxRkRlREhIkb3eg2mn0/g8bP4w6UwiFzydby
CyBrtyK9HdyBFg/Hqs92VjMplsJyt1OGKzp0gEWYrA8JDlOEZKQFRGxtbaiQkUOy4iygHnNbteSC
ClXp5zuatfJ17R4AfinIEGpQjwZ7/S9rdDYyjZqSxoa5UuNmjUCcyUGW/+yOu8e61qAN12gnxYxV
8bTAvRbXoocrSvIQ9MNQSdziPUMJ+GzNH1j/V6hyxHW3qEuA5ZMdh9F1h6rishL43fAh3kgaX19r
D9nGdEvphSIiEQafbw+r/6qQvFRruFmJ2ZwwIaLCU0FRmrTECUWa+mLPjxCaAqayk13YvbEIL0LA
kggQtKZeu58LND/38HM+VpNcv19XTkkIBiBUK8PGNx1/HmEng/i1TDq/y+VrL1dSklQiIIRRuZrY
AnNuFys0OXDzrVE1TlsQbA4WzW7HOkhS4afPFxT2goMUPNBfKLm260Kwp/uDY/sIJD7N7TTKs7Lz
5D+XnsFG+OowYz9hrMcxGDwsBPAynutY+7HoPQ3shCm7apeP5BYUDU5D9YdAUkv2AfXbXzB574Kr
+eHNOsO6WQYv7k0pxpivvmhu8C7Y6HlKkrHsnSmj0SPfkJl7gnCZ0HDI8PPljQ26rGJEWBxUq4bV
0w0uc+k2Y49gbJxaOISmDx+OTdFSbMhZYd4FTXpa6MIdK3HcmP4Rm7TDMztJd1vaKVSIOGXFX5qy
LxdZV/Lm9St8I+0LUKA5nbIq2PBFLsqFWRxF/ByZT/32KTkBVn4h/ulKfiqZfKaIuPWXRX2KycjI
PVasugla+bvDruphcAx7jSfnhytvxTWnJBfxnAV3Jg8BCTqhMmZhE8rZ4PMBi2GqSgwJtndHpMhG
VNes92v3Qee0/Yyv00dCKFmteGt2mHtaNAxmAE7g8wB5IKRLBK+duITniTOKFLKRmwuU4U4D85Mz
qJUltbs9zUF/LoT3tSz6Ke9VB/y1mHqO054eQDKwHWaW1wQ09QEsp9GDFLyfp/iHlnJ0eLpSse7e
QGqYikAPMnE3wQvE697jhEkgQ6gc74ed4O7rNL7Yq3zKKNRFqrkGv96D1VfedfVBUqQO061BAFXW
ZBhmqiqdcaKcdXoclG5a+mNeq15xvE3sY87yn5dVYVzQ0hh7b6EWgqQPfXmAa29EvocVYr3ksn0o
N+GpiiuAA9I4oM0/uPQzJaL9/kFnSwi91OM0tAZrRQHGiHhw/OLP3YdnDdUp1adlz5bdloR5Q2sw
mgv+gji+H2ZYFPs/0aCclfyCaJLcBGXJoOOPnpWNf+5gxROQixaIcPmZwvyYz6SYJ90N9qmaiep6
LL/G1R+YDutQ0ELWvBronDiQon+0qqWWsj81ZLMCYi3nWLLt2u28lbE79SWewYWj4GEX2Yt1eY+2
SLYsrQneLmalKKOw+BO1VKxqUeqCeqoQKFdsjwslV3vXM2FX+YobjBoKZXewD0HpAgub54ISCoE7
SXyXwdFolV/kIihX5UphiENKbsIwuB14bxfVHL20+c9VFtyb0U7YQJ/GEzmuEeXQEK5GhiloLQTz
lD3Xl2nARruTgCiT9eugvEz58iza9tVKR917jeXJM+PjCq9sSiIOK7oJD1YfkHHAjCyDlQlf2xdn
Ocmu+LNvbHVYQNCuFzR62cGritRuBU75qlDLVCNl02UDZMQGMuJ0TK/5+/rXA95EwCjSLgndft9B
Q20aQsNsqC0oEulBdA02HdneeyqIazWtyl23eeHx2RC0PrYDF2A6/2WFSIbefUPH2K2wqIEAmrJK
8a8bW5xSAKUuNLyOsn5k1HEKk80IoFhQMSwBQ5SMKsIxeFqMfm775zcZeZ1JYTe1Jk1TQT4Zy9wN
f4kfy6sAcxYBcV5qa3bUrRKbXF1UTq7G7uwrgkK8h6wPkH8W0qtjEyvFJuygt3Q6qczoLshGVPo4
/YWClNCFzjBmDyVE56Z/KxehkczB7PggdSQbHKHBdwxj0owAePOfj4tZlJJYD59I/mqvXKQBT7Ic
mhEe2ujUjnD7EyjwLP7dv4CLyA5kTqguKZhKrHeCW8gP2KwsNleKAKBtV9pXbCH2RkdWwERfNoV9
jD2sVokRMe9eTXUBEqmQZdkY1m6j/OK5uR9UvwmWPItQr7gAtGxPUpsQdgyftjL4VCcRWrVi10dX
OXjaJ9ETAj5wLbH4NgD2Qf2K99tYAAfdSAvKRm+ZIxnCthcxZUOYeiaqlNxk0ibTa458f5V2GLUn
onjmbWmRGVEcIGrawCcCB/qMMAxhQRmkQRHDBdyZpupdo2kyVMKzZvGuPV63PgTbLEgmmwdzw6Uh
j4spKJ+7w8b5rGrnbskUKpnMUjpo+AtZsjoRmLWfN8b1in0JKgUgPPX9PIuz/0lhd8OxgcBAOIgT
RMVuVntMWP8xwD5lUSZmvUpxap6/Aj0ty2UmkomQ6uw0L2vDxxk0/xjbXJAK+ZtqqoEj3iCEivCg
GzBxVywT9Fw4BbZuaS7oiMqeo/xTUnR3av9KCEjLcoc6g/uK7VHjKGH9V5lgmSsEfUzSSUA9Hc89
qq5TtiI6Seh9QLOIDxrPgndY2PEF9K2VVB+iRcPmt4LaClK/uh6St63jsU1CyPlkaUB9nomubgYA
gbi/dsmh5UEElwhVD2DURHy9PM2hXd3VJXAu6ZmncyKBNcZ1dZZEX9ym0EqldRdbU8AM3DJXBq4B
zsyRGF1T0AO2c/mFb98NCWav9myqAWN0drsLDGYDAFpzznIzg78lNEOb7SB2G16W2AjjkjEVAGVI
HVWWeLHC26Q7d12sDC+/MNkxIo2v/1BGQXbunwF8sWruM4kbfzFsCD/hNvVzCeCwfeJdoihc31Tv
BJTJiDZKbGkcOCA08DDBSMhCAF/yx/lqnL5aeUT3Z/0oJO0R52r+iwZ0mX7uBfiFobS2wyyK+9HA
CDDrAEKToTYPjnTh0u6thnC0Nkmx9fmvPhKRgJvauY+76qlONcKgUEhR5mUY49K/dw7BLD/SSjH7
lM15KGa2MDOVuVKFUVoI0IgFHWN+dNNF5SK87pyxYopVnOdX0t5/E+SkQ4A8E6syjlph7KJ/Q5Cn
pc8LkE9g5UZ1nnJIGLDbDT/Tw5POS8YIPYdPteETxETWkiOtB9qp7QlAKO4j0hbwsZDeqa1GazTf
M+fLWWDGpi95sgUPvoWpEpLfHszX5wQxzRK5Qn0nrSynczT82s8Dqh2XK9F02+MRdMEoYGtfVmRm
mk3caIayQtON4kxP1iBznQMPbT2D/nLUtetrnYYDFdEvdqf3P5oEB7G/yw1w+ECQL+v7OKvmk+AR
sXztk1FOmVv24vcKwICbX8K+UIhQcrKj2nC/u5xpxOKOPbM+6Dzpl1n/RzNbTfW8YKQx+mtV3+16
f6TsUs/ka1pKgNhtaNmk1aqKrKoDC4iyrQT0Akcpe9sbmCvJJJRYxgqFciTcC2D9ZjxCS58esXTl
bo64KieYuwQt2wgSCvXCf/gGUiBdNyELeZyA7D6DKbmi3VcyVSwuyj3Dkc5RZEaaN++rmulpEnfF
XbPcJAa4mef7MaBa6sy9EHQDdEM7vPUBkGc6HV0KlfRm3qrEggBB9+85Y/aKIqmt23tCQvXcMkYN
O8LMvWpOqeumMaO6lJFYO1dGuDR67CYJCCzR/Z0lA7cfjm6HPvzNfsXPukrkK37gRofeqNxe1Mgk
gt3bpRfO8qIRxZcXbzngzjlebqdnOW/6Bntw4P1I+jUxEMCVk8lSbkGsODf2+hKz2k2m/IdKIm8p
3Bm59u53bzfdrMJwGh6PneQ7Q8R5C8WNTqmqFLaWDdehXYaz4eJ8h4raSfoCcVmi5DtKnpQ8Sa3f
V2fHj0wFnm2l/+XzIu1/HvZGJqzDr7aQXgeuI/a9+ZNjN5qnvODK7sO3ZkxpcS/QZvnHBT0bTpdi
BivRwxGt4EfxtsmUcduwsL54JACbZoQEEgw/P8JWqpDZNB25BRV8U2A5srQHz/62rLG94NVFBGeT
9DdH+xubYsg/giIOEvBZNc/351qeb6CiQkW6SvtjcXMnhkRK+8eD7QC3Fhwr4XjiTDYBxsA+10jf
zjhw3RoNqPUJ46nzqhhvUmvFQMqxEud8ogUdq7zEuTJkSf/Do1aYmnsLyaASBHlhfg9z1p2UbDu8
gAq1D+5uBqu7JbfemRfCk5bKBiMgbPF9llbYK09tV67q/5mclfifdQGbc7P8WYGlbnOaT3m7+vBG
keWuhHbKKCblt7UjCnbiKCMiUJGHlmvOGHv452UNmSOfSXBHeX9L3KD++zeFa/O5Fg8KRpRg2R0r
Avf2aqDU4fy6bzLdsKxEd/mx5YYRgGUeg9Az3scqyJ/mxwLjKUyxcNEbhAv0SAypzl8mm/5mqH3B
zC02cnca/VOk6mmcUGIz5eq1NCuq+uBnnP7sbUi8aFrkuATpMHSa3e1kFX8ETI2jPhrzIUMn3Fb2
E7aDqEW/p+3gAXLEe5UkgVh2wc9nUsZMzP0AyXnDuNS7Ln/9Sfv+eZ82guBAiBopajWDvOsmln1g
ieLztuW2Uj0x44boJMUEtHehXdPTvPUHO/CFNncmiRoJA+Fi6MGjrOQjcE0CCilXyzAdIp2L07Db
SMDhYD0OkZ/GkjGKi2UO+ZwebbT+g56zlcOZMJSIweD3VcnexdCjjxATSbA3tiRu6U9IgpKBEARZ
z4Wdd7GqLuYC59Isfm15vgsAKyaUQr+IjNorSGjpKgwD324L3MInMpqh+KUGKsg3wXXaL2CtTMxp
sTIOIedhJ8fY8keBP2Q/2wPyCJllnSKq8xaJb4DGnAGMnRRihS7qY51Q9sduMPHKO02IcyHnZ/jr
6rbjWvS6tp0PMUJIqgSOK1gWz6SKJV4I10QagK4CSIR9kNEBp19IZnpW8MZ7hUgEUM/jQeMAvtEy
meQM6FvJjaDhC+bjMQJNwg2Vkk+UeE4sWsesigbmqxqGAWG+hbK3MIaX1ssvX70jKXWCO9zChFGr
4PG3PxftQ0FonHzbGaILaAzlyIcbREp6gYPhzm+1Yc1K6Ndn2TkFVsi2+RIwVgf9irbQro4o3ISf
AgT6ljKNLjbnoBHhXo2XFNSw9WEkEtOl/KLUPrNXWPlfR0RD/76DLOA8geZ1iTfBJd8aS+R33TUY
8iT2XewXyr6NS3k1bFO0/8XJtg+w6LmfYiu/WbdqJm5MA6P3MOK1L3laaxxD+ltpatB+De9X4IyC
tjtbnhNPH6Rayq/SYQiW5QheNDkOw6wtqaIHboE/ZnOT0Xlki9PYI2tD6a4H0igSdeY75la09MZF
+ZYZY/O9GVOG4tconUexjb/EOfZM3KaQULrTlBFNtUqX7E6E/DLfiDRL4dxvfQmIHKjbtXTRHBrX
zI6wB7csklLJv4H/BGLIrzyXZ2KvOjeGWju1pJR4pJiXef8LcRFu20qvd5ygnYZteRUlAQhvjwtE
kBwZHeL9wVvscr7jaXxtLpc11rI5Cw6UBvPGWmeyzOdpIMThDFVVZLKugwU/V4+AxGHSB+gPqfol
i5nKeqIRUz4H0mXSuFLwONMtcidzdIBiflgWKXttWlEGSGr8b4a46FnVWx8AXPnPDplHa/us2Fkn
03OWDuYx+yO/WCNbroSKHTuj5bL9EmLUdfjkPZz2CB7i0tg6sfY3fV5pp2SQbHcUPgw7XrsNprWR
NU+NzpXatK3KkYcLNAuJGLpVfNvZds0cPnV5yNzt5FI8E3RyvkjDo/VUzNKHhSU0mKLt59pDccAP
Nfy8i0owJQ6MxM3G8UTbf0yFq2NPA4lqv6Aw34gbe+GDV5PZ3/A/phnYW63DcIHtuPPJJLsKiq2d
CJgldJ3LxFyjQnkakBAQdP0XHdbRgO2oN7COkW3obxAtI47BabmLKUpZ0oQWAZwpz7QDR9H3oH1a
Tzyr4sP/QxKPEKvH/XHPgE+Rt6TYRC2KTngriVci6GgyDh0/BxtBS9ZZLhWKr3PQcCteB+L/2lwI
8SreoO+zJb3mDoOkHyEVIcs2wUqjGsuCquZwPqFBMn5tJcNuihanpSy81J5a2MAHQ39dGV4jYKS7
+SSx02qpvDkqjesKYFoIgbWr8xD9MY9NSr7GR5uv/L6p8Wby2EAK9RtNxp9O48VbIsaoa6DvXN+V
r66S9jhdxjzWyfloBpMqMT3rm1aLzNg27WId4R4t9smornS1Qu3OEG/PiyZHDznEs4xxcNUcMm+j
3obT31NGwt+qp7Xgb7rffdgBnzFLN7iymjcHeHBYj1vHWEEQGU0JjpEetgdgdnvc0mpNraa8Z+Dg
tGuuHTBmyaXWnOgQ3Z+rHHmMw2UBZz/zRSeBkwq04oEZCclcmkFqWOz3pWgUmIf88c91WVuZaZvU
0QEzcQLv8Dgkm0X+Mq1chsCfNZT0AgQnely0xGJ9Shm9MTXO/+J0RmwxmgbDSaXiXPpITbOGeogM
zkbmTcfRkhHF3NHUaN107ERl2oMN8ngXQ7Yn7wDzCRwWnMOiX9UM2JzhQyAPypY2+7u2/q8LuGM7
M3HczLL7kj2kyEXZlinnMEIpk2IhwjpyD3a6r3DlFRqPpN4RKyfflqRHqTrpJ/ex+LPKBxwnD0ay
44Gkfq1PvEGsxlcxtEqN0Imvlm1a/gdszuimJD92JFfm9cUgDX3ef7Y7V5c2PtWFNfSba67zlJe+
vgQMtKxx2ciDFgouRPGD48aziuMZQvW3QS03x3paeHMlqiIT51bgEV85s4jYyC8TmaWSj1Uu0wAA
R6NL1XdZvkUj/2/mWUD/dzEpqNOE1Y+P1VeDTO/7Al1TuFSNhGIGm7IBsq9CrPQma3GyPMnDGUu4
D3VS+3z/8Q5Jf9V1XpWCEmexECafZ4Sd9kWRHeHdSt3cDwIg/zCAaVwofS0RaKsL1dUEwlkyHowL
VrHTDfrxrZ+tLTfvviaS414MKyb/jR8l4I8eDFAEeaDWc7s0UsyQyKZVy0OAC+V6FO5RD6zo+3dU
x96Bazq/+1hyC8DDB9LSGVA7p7UZrp1DWUJyGw2sOwb+lGv2qB1Ihc3iC0fj70UUTKLsASj7klMB
wraTaeIaD7LjZ65ZVHd4aM2YU27s5JUB1S7gfzp75r3/27qqLKNvc+j8rfqJxX4ekrcHMUVgnHVT
iMFJTz5ArfkSOVafRBhbqwXGlVJiFARAwjQGOb0OySYtfJhELpNjGx+Ax4DAYUqYq6eqk1zhy6H/
iR2WWFdKEuQ3vlosKZUO61fVXwG046AFM0Oc4KuEm0c71TwONrHSvO2hY9D/HAh6Es1f9F6U+BWF
ASNQdcsjlH4jF798EiKpbnbF8FHdIj2VCe27OMs1xsC7PugWAy5cK9qNw3y0JMYWpX6TfhjdCGZj
UbeaTHiDHk0BxIp/dnRyKcKaObHkfxkRTDOkCAOmXLACgp/d5L3Gqnvqn11vjmbn8jrJlZmYVjrp
7hB/43J63IBuqEJIVg/1w5zZWOcrKdi78IbiTPVC0M215iCpFNff52vIhQloZUA1EvJ+tSPTzytT
gAVKPw6OKpbdF9rW9isWrisoaClf8XHH18vcBfP734edjuIgV0Kqvc6GOkWyLCUqu/K9XEicX8Yv
F1er/2LLb7KNiZDJVja50OuaSxchhY4O3+avQPlmhYzxDfbWODBJBNU2Lhh3Mjh9WNiPbHCDfGhl
mmzbOoTJNE6m6A6f95eE3deFJL59GyCo9volfCh7WCNJgWmgbV0G7nGG1QdHP352EyQXdriqTqAE
tcF5HQIZCgLg6BiCfjLLwS111CpvZvt+XWvTFULihiDvF1cU8GJoGA3+Zi87eqn0vryu5sVS2Svx
NkrHIXpvloRQRWFOZV4Xcs8DqyR1xhcmdqj5j4rgxWhCNyQux7YamhgKs9SXLELuN87Qm/JBLaRl
YwTh7TfeF6Sq7MhzhC4sAV5FI5pjYhgu/edkYlzsG83eAzBWB+zbPpC55bfLrR+aNKK50CBOoq+Z
iHrGhkKCi6CfQfmD0rZvCYlsX4zjr7TDuCeemVtEoWKI3jitF2CeDuVmF5UXYFJVib+yjvQSI3hr
/GqbLXVvbI1/n3Bmxx5uRM2ylGpP+tnzqvFn9zHN20M3uVLbtIsJfrowcdyCdTgPVNU8VHLp0Oju
/37S8OW48SfUXkYKVvGnVWcQjzeBCcBXb+zbazyIa3A8dLd7S6U+KG+Wn4KxhdgQhHn1Lgoc7w73
m/kMKnSIl3gRlYB0SJy2llukG6lJIpaia9qH7dTuPpWsnOGAd7HsVSpMpZClNAlQQcPvtOuXgufq
FnG7voNLZe4IxPnZDTL5mXAFdH9rbP/VVrBcw6KmaoFdVIkGmRsftkEJ2NR+3N0pIwtA+wkwTgw/
O3td0q2El7KeE0a6w2juIXi+iFOtdXyO11N7dpdXxc1sepuHTwRkR55Fc/9mFcPW7sUlf35xe0YF
EOmQpHx6ePfNEL/ikNDF1HYwDOg6AQ6FTnsQCFaTow5quw68wfsWgumy682mM9yyp2usjHPA3RR6
pLkIeLQv89+RFOoq67iradMAd5IRS1gAZAvAAMmlJhyNMWDBOVUH+WzDwecOoDsD88IFJCyageV/
0+fMnUt6/3HZdlHNoN2/HrZUWmdN9+V08Ax1zzZOZYTakAdUD+CUz0BGqb8gzAmb0T8YC6YTUJX3
73b4LxT43u0ydgFjxnzUdqd4Z/BslkKW8fcEC3rfffaaofYpqpOspGteS89lBYADVpSjBNrZuuVB
TJLjmWYTSDma4app66NKtzctWjiveZSW4hDgGpexIdHs+cLuPMno9qyDgLYndFmzeXx3e3gcX4Ze
3RRPjbNG+4lRcCjyLW0W9XpahVoSPNCCBkEsnEwN/v24Nr1tNG0LvWDp1V8Zf3Vzv69YYmSGcKty
kVaQ4HPBzj/nQT4wX2NYKcVfsS/1icffzxEWZ2QZ8pyEt2T0Uc2z8JuGvNGu5UTi87JBnQQybylr
Oc1jjaRpbBtEDJ0MgvC/OE3uVt2zzQRoFaZ1xkVaSengxpTmN0d+8wLj2Y4+cr2xQHNSXgwcd7M6
6UQia15BSh+L6RbcpP/0FEEvPEulE3wa076FwqkHTPOIgiJpj+/z1/hJx2wks7pcCr3n6b2Cryee
2Gp6v5A9vs4nf3ozIFpeLn42vvhhyUOI6sDPxD5qdrsywHesUizWdIwATQgeXu/IrHNfIbY4EMVZ
ECdt0ndFCsGFTmK6G/SQIBBaeJLNL5LidhRt0ExU3w23YsuhsafaxRRY0TVnRcuM5KP2Ox9yXuzm
FDTGr+eI6qoB5A8TYSY2UYfQtwfB1fa+9DK0ph8sGNYYUQNEGytu9SDh2sGpae0cXvDUTvTZO4eM
8ecsqzwaRs+o61ePYUNTNkoqFfjhK1ROSJaMSUeP3MvSPAIpCezCfMWU0Nf/A7Ag3qq49IofbYUL
By4wzZ8ubf71d2dcvqmZlGWDVc3/mMnZnSw1NoQxzx/+ayFxiv3FeMJgws66UTCniTfafixz52wT
SqxX+YSCBrdwZOzEjnfOLTDEAv4IWtICA9Tu8Xt6CJJ/kz1W7MhEpqHrc2sSwBoetXBQybTxh/qj
dniY4hCQdmN837/acKnd2rohWb6+KeMaXTHhOGw+FxqqNy5w1XPrtSnzpe1nsfxh5NKfI1KcsI3c
VH8BeT4skxrmoV9xntJzmJgOTPmYJFsIJYFNA+vvcJrikXVOYu1r51Z1KUfSfBBAC8eMH614F0KJ
1ZRtuOQWG3mKzpEu1tLvaG6OrZt5bCU5FDa9c24QBJh4fBDIa7dNatYDvIwsVwV0EbPD9JN6XBx4
sTkR+hMj62rPKd5hJuhybse6QIEFDqteYFpUV8saxl9U+2mfiUFWU49S4ZUs6FSKZ8bprCV6lHAA
7KTHrWfVfR+AEZUK143vJk3Zi+YGYZaXxsdrsepaJ/jp72WFN1mAfnnyKSGf+ZYYEJvU302wOcNb
NFLdX0yAZal/7tImn1rQqwXWLXqLnAmsWPauvg2Ay/hHKN/TYioc7cWdLtq8vKt/Mg5lCIE2GQjv
GvohzpcacjzS4jbdDBT6jSnq3GjC1Tlo5zWRs9o0uOfvdr3lz5uda56b4G5LH0t5dAd+40TK1Fgf
9WoImAEoj5tV9LBXqH1HA6dQj9G0GlQCNfCfyfpDTPpCWDpTqgZn5D673smhqg1g23ZVhU2zVmQQ
Ikw3hcu2n9G9D3pSZkHLbwS/WITR1UjuyE8JEMRYTK8/rmGFXPo+ac0Yhn86TCYj/m+BFafA2RnR
ciW8PiltgFw09r6pd7phq4S+vYUMLWVfs2t62SakjgWw3GYGvKtMjUPrNWpa04yHdZS2MdDdvF1u
Iwqnm6jisYOIjKK1yagDCWzyRrR4X2FaK3vbEe3DTECdykYlwNlwSQMH21Hz/rm2mgoBJ6+ImNbv
FJb2pKcCc2kruSPDj1Eik/1SKlLrzawSXrcN33y2sESnsoncCG7PtZld+yTj1vao6TEaKgpJffZ2
SQsphPJjeptJe2Cx4noN8mETw2L0iMsLQyCXkH4CuRfp3Ov/adoEkOPapj4YrlNRl8yfBHVAQYqt
MHv9UvN7Rm6sMswA056C84QF/1Oi4loXt6VU82V+sY727QCrJAurlWef6rgKtZJycTrukJaCLnA1
IMfQt02R17y2/sPLpd3+e3HlS4kNTKmjcT9dvWc4eXMxMrti0MUNkGwvkBwpMxjVif/itTpSOA8e
olu+jgnJYy0wg8/TrdrRuYTWN2y/2CYKzZJ1sdsHQn1fhVuK0GA9rIahtVEYjSMwabrnVbG+ovmE
ZVyd45ENfSYeMdDc+xRG9MiHjS2NE3/yaFJCcqjnqoYKB3rgtOeCNM1UqFVjno+ModdEza+XhvLL
FR5wEJsvPHPlBfE6z/yC5nLUnXQQlySDX/1sx6W5o2xYp5R5RBraBRjIgGh08t/7+DfZlzahwRI6
fFXxFy5kNtKS/2y07JvZepazzyySlRHcU0lSoc6ANfR81EeOtkGEuyRt9f0EzsV3Y8ne6fYnl51s
JkfNdCiOTLj3agq4KOgJRUxYQZyYaAR9bXoJULkvHsDj8ZtX+VYL+eFjKzjLH/vCp4lybqwP3uDH
Q6Zc+I+2ShabPLk8YY+xq3OYnqGsw9EpKpcTqkRLCT8awCSHFwuYm8dlG/lKDn3nqyuzdptAa8gO
3HxKcRZ0zYeCccuSiMaVb1668kJTKS/lt2PqWNJWiz04QabFrZeUewgHrTwDtyFXH2tREaMv9Pi1
/xk+6wNVbP4MwVwzEzrtAj+JCZKtar1IpTDvvIGNhaYMLD29ho0Zshx5F4PTOn0aXgkP1u+cvxhW
irehTAxstLleupczBT4vt2pAHddNDiXSHz5TjMoZ6uTOgZHzQOmudRP6BcPd0uZuV4xIlN4cSYHM
pRiP7oqe2uO1XqFX/oYF4ncNeHao5YFdEk6bHS8XdmH0II/l2EC3KIXD9dOJKcfmyT4rar7S/OtQ
wyR6zog97OVhLeW/XFSqbex2Qpgb7UjnHc7S6z/94pIw3JOGGnvEgFPjtqkJQjMocaPj6Pt3ZYEv
Idwyn2uzBiclLM/a6PhmTrks0Q/RtYsObfh9huMwbjmTEzrMxgQ4qzfKoEFq6Uqn7akUhVrm+ZGF
eIa2iSCW+VoHzU3q393a8k/sGhENVxxaB4oBGP9JqA986oASJp3ZRtMhjiJAG3w8nTRuBFgN6eg6
8OFG9tsmFAhV4/bEm6VH8+NxyxAbAHmjWjUw4yKmgpXxR5oWC4jFFTbFLhpErzq3T3M+u1OByf4H
5kk5kV12M1dfGwy8+GRVBVOE0N5e7GTulyTmLoyu4yteNJ60/8pi001tBwWf2XNoqTu21B6g3kdw
0XwRG/+Y/1B7pQzsYLVzYBcR5DmxdF3WgmXFvN1MxCofQtVihhQuVaBdcXWplwyOXO/W3oRwDqn5
rdgMsVWtMuxyHZfZLd00m7bgeNzGER2YfZtZCugwXgCuM0MQfu1yQ+TApyRcgLKhnUS/LQ8buOto
85umn1qkuS7/rul+ysO1zPaTmg/i6oJWJbISFmn0R/eIcKgin4cFTYafrNsD+DGR4qIOy8JtOXGv
60SXf2PozSgHHFrvlMscHpFfY8hnf2VKwt5OGJT6mBNefSY2Ne9HwFhFyOA65rl0r9QmPDKK8gmc
xOhCXNLws8vGKDHlRisnBG/XL1KvsbevoA3bNDs7bXPin1D8K7AgTPlyNUloRSsBstsn7VOKbpM9
hRrZ3fVcpmMcjansE9yfWAnZG1rHzx6K/QO1lgaopUS3GV9wr5+P56WHRWDvsIExKDjeDyrSZmc2
nLILeBaS6H0ohEemC/IEkF5EQo9gi0w5KhS0/hv7y57fTmPoQ0tbg4OAtKLFSZhs5mRDKw2XtIKO
27JMaU37AAuPZJLcO8bBdr57QGReQTrHDQSqmrurZjg2KBfoKeOnCsoILGdssPxKUFeO0WrGOOZJ
4kUudo0Aoz52lp0vqIvODHaEk+rPwLw/8j0LyZLUL5Z5rWK8bZA9GjNRl8usZ19IuQV07X3pqIBK
WZ0VLP6elQT9CYjLFVz50xx+vi38m8uI5Pr3dO3F96KpLcBJ+CRj9j8vg0In2P2qqTMMKt40vpXt
tluRn1HIA/nv+NXfBEa4Xv8sO1nSjrh/oOzJqJ2YCdlhiaC0yUQMaF1l6tko10p8Vh9II+FDJbqK
C/BI4JNr+ye286TGUbfaXO4K3Caw4t7NbFJsbQFJXvN5SseaXju42u7nHe3dXn4CiVnWMiwYI1gi
YUEi8aAduw+VP7xedmIqaKhXPZ/xymm+0vg1afLzvxDD6qsR9+o/zdO8HXkxKszAjY3ECioXIP5m
cAjYmo/mpQkt69i17gWR2RiZHFbSrKfnlVkGH//oYDceMvPHUfr3Bx42/B+DGSRCy9np+67Fr5j5
PpBIXV8M0TJFPhZPvFpM79BbmKXCjvEsNwi6FKPuYA7/lEdW0HskAKNiAaV/i2oiqQ2bFWHOP5vQ
JjoGv5A2sc0zu7V+wqo9qWoA0qTtX+ZNbqg4nm7fhIx1vi96y1uPwE8B81shjL1EcdtdzfTCzCfG
GnLq+NL0HdgxgnaGduXFmqv8fs610WvhbOW6MQwlFRLZ6RgMW4KPaER/uBMa7RPKb3NGvECb5acG
BnJgzP3OKgLTWL9XTdrJfBAXPiKlOyb+x1MUHQQ3uwgaTNWWpwEVzAqlP5OePYrAcI7uUGZgt6Bb
OOKtQPflnFn4A+i8eQVqa76YZPcmTg6CqhQ7LKFKUbpyiLxZPByS8tlZWanBCluXfemg68eg2Hoa
DgQJ5HQPTDWtf0IdhgZL95jXJW8IuVfJHw5guTr8cKJzrTBgitGrQh/fz8hhbYEnBJ4Je68QmDER
O4ARs/tihzWjoq7fCdsAQH5P6+f1GDenNhlk2V8azSNMxHPq+R6/7LvSOpEzW3yoeLmiL8aodgDu
1ldzGAANFsTedJKOwMJHiq9+ci7zrL5NbmOG8P6g8zksi97/mBM4k1+a52TVIyDYyBYqaVPkHRGf
b1TbQr2nhZ2iEygLbjfNfekIdEa95hxwkP5Ks5sJZnOIKlzLNTQ5Kac/ZJ7bKnMLfITgG+AghYUD
ZclIhzxEqFJSSaEDLtIKRvQyLp0daK5jjh+5h9K47B2TcvB6ud6H72yHxCmxgTU1OemGOBC/U8mc
ocd6LzTxHjj0pEzCcvL/j1J3J9bpUUSkSJWyuu1/CVH3ygIwY4ZSMd4KBgb5VqSXL9Xza8pJ1xfJ
iXh6pwqrjeutD66C/sJMSjuS9JvKtfYstzoUngpf7TK8t3fQtOi0I88Kw6zQsILwpJQNR3Y8fJzd
bitZqMC1+V+dpmaJ5NfDcOaTdBv1XcEleEN/DuKt5JDZBSLcmXUS0JU1dipkrqlSziYBtqgoIVCY
HCwmGoD1iQ+hD5j3Cfh7d1xNVmndQoTgtuWjpShpbrl+TE096dhfm/SVW8eUCwYxotgxn6GlbnPg
lVTtWkjlPppdmE9sDX9j5Aeio0ruQ6X9cxHbQvIiozSu/rcq+CmnjWrsHdo6eYh+T9SCIpf069dr
pTGaWB0bN4aHHhhPqp8DUDCSPTf9t+sNHD3gIFdigvmIztZsjPjFDh0JxJ/3jlzMG9KIktZu5pP/
9fo391RVY7SEb04hcn2lT+R13eA1qOFNv+tM14oFQN5LdsscG9Ie7DO6FfcNwKw+RrFJjVXNuQG1
C8ylgb6u2H3N9MZmtRL4j5NAtelQXyyrnND4tw4Wo+a+1dYr3DFaowcGANInCkTItRX1qLKLgqEz
JodaAZd3+35Lw4oDTsG/0lPsM35R1HWHD5AgjEICQ4PcLVeKRVM018+wie97MZFa/CilapbwNZG/
bOHLFVgiV/vtYP4JjJCcF4N02oVouptILr+BRKwXZzS86+hncf8CwRznZlQfBfNOXw6HAY8Lrnrt
+W3XxEt68cqvBsnn2adjTx9LonvgFJUeYIK8M+OwJD58A9ozp9Pxuu7AfqfJf+AG47Q7gneqEpCW
szh8Z09eak7U9uOrI7m01mmnU3pVBs9E6akx/8jPma26p9weSv/0w5tYubLZb0y8z1oQsrJNvkm2
jSBftb3g6agU8k04BP4U+xk2BOCI3pESr/2LsTP0RqgCBX5KVSXUShAWvYXAzVjf0eDWFFPSfHek
adA/LeuODoaM9Bf2emj4fFtmhwTyU2uY80GUFpFjBJSwxheYlX3IQUG/vC0g12L7pYNOdH8V1pnl
fjsgGQYTDSGRLoSbG0iP1lj73RC4ZYywMKfEvJAbuI+ILex286mrsAtbHOtTMlexVanHR2n+h3ih
g/U4KVCtlTnYIWe8/uGtL5b0bZVQQ/vQx7JygdpnMfK6atydX6D4h7xELmEO/JckGxnbMGqEEJGQ
iDiA60CSKR3GLfEvHdhOYlQev9wxMkgfKmjTxa8xtVsTbQnpwG6akYd427e7f3dPEfOR3HWDXJ5O
f84wUzZGZ+H7okzWwkVJvGSyWtUnuiMf1TutKr0h3XfurYMhWr+cFZ471NV1LQx7k4cqTDBhFAcu
KuBMBngkkfT1Cyq1NwXh9mmArHZ56tORZ8q8Cp3CvHKg45lP0nPFHS/6vyWWmmAZCMVG+pDcIeOC
4fGotPU9NAIlL5+b9ZDvtJ9Wx1Ygw4qy5YpCHNrIis19MFn2F7JQ60/vM+cTcIj2SR5ac4dpsczs
Nc/SQFvOXoeoPiy4Rbo/AiGqZ/zN8swDf/C4PTMGGrQ7CioCfPQxFCLWE+trJ3RWFPCDih4B3H8Y
Yl/q0sHCi/6wb60j2UWXZ6eKO2mqmyK+tBWRLqnOzjihTBhLljgO673RtcPjY6P4xI2VHRHGtmO9
ndrpvZ4yTGYVQuPgldn8Z6HNp78NojLTJXGHh0Lu6rd8dEkfAjkofxlOQKhPVLOV6EmKykSyJNHp
zopKgZCjCkU8Qh/pKHExC3yjZ6hQeX0pxOnVpDV8BdLZYxnCB1eilH1koltAPbDXZYi44X8MATCV
fcQQ77ir072KDzoncjLfevV52u8FPTY1BjL7BTBeYIbz9KyMjKbzBFPPC/utBxqu46Km8DHSoJnM
pxlG2/IMSu776eu1HY6ydUTe9/orzt7kz80GItw0imr28gpI9zoAxY9QjZOveJyXiKPnccLbLl8H
YR8WG2CAONzoJKHftoGHaFPlhcqnTPOqze+VIxY2hi8daiiUsD8BGbEYcmHT290St/rqrhyqtI9X
refQLsy49O11B9iCGPw3HyClaL03w9b7PBeBRBJcqqOC/ZdiTo+/4Stvoc1DRXOeAXSw9rP8Udnj
03ZoaynoVBFYROyW25aT4e0xH5HBeOh/pLvsL6zyEESbbvgrwptNySl0d7k5T/tDxci7EDXXZWX3
0Q/G3wEKITEsgrKW8dAX0uVM0ULItsD52CzSAd1LiuDVg1/sCTEGhvdeBoGlNEY3WKx+orxO8p8h
fh4g2tSCtY0WoKQQufhvnWM8F73PXfOSFcGquuWbtQRkaP7tuuN5xVYicvxiWn2TMc4Y/kDc5EXO
Ar+CiAnQVBlNwJVAqOmd53cr8sLaB/VbONEwGgH3vWC42RQgxlQMS4fj3vbbf21kbDtd7FBXtgzx
xQRKQBzlRaCCNNqgFuN2ZpOX3AZbWTr96Q7t/p0zyIbbCmW8xVhImf5xufX4UeM6bWmSEQpF3yMw
J8ngPyjzz8qi86yJUBPzmSa+791dNWO+B519hUJ8haded6ifDir7gkwGK5A9q7z63qXSLTacKpf6
f1rnnuonkrxWo1i9nbr0NGUSSci7kAGtXbzVyhBeH0vJSGNWCjw+7K5uou9A127AWgc7U0aAgX5H
4TUYuMb+lRhfkyr+nIlwxWMKIx8W1urJM5x100/b2cKp0sPIYi4tJhAAES6I5DVdMyBlt+5GZHZ8
L2myDUUmUWtOSb/dbSKp/1Xygx45BymqAyfHQM1M/LEEiuaTBChYhd8pCFfZVuLtuCyER5x94RIq
9/kTUjLDwIIOEzmoN7kr7z30YAZEv3F2PHJvul5YcCjP3f6piOfbICxV1Te9OM8zQu+7hLMNuMd1
B4VZS3lY/4XxNVhRoozwV6JogvCXFUXxlYA7yhSP4MJeN/wzfdQzthFVHmGPcRT81vjk4U+zT+C6
+DabCBCaPnAHBRO4bWZyh9fYBKqqNiHAVOt1B64ZBVcfPXAYkmJgkUCaQ3g9DiM/AeTe/I7yeuzW
eZNiWv4jM98ap5hTasKr9eS7EkknIUPBJEyH4avh24kE8y00Eu2ZW1Pgmc9ebOvtmQediFzx2d/2
MllKrZL7rngKfnQHtCRKEG6wECpBI7LtRRuFdp9HXBiP13e6deJrcYkD2jeorOhGmyfo5KPfSYGO
G0B+8QS3Qg4CkDsyiSUQb80bzCEPxTUMz4CjJE5jYuWLetzJyki0GOq2W9rigLamKX+oYqidt5jr
gublPn+P1MbiSa8Bxq/KhMGQy1r/emPsfowMI8IDSG7DiK1NgDiks4SzJW76F+1kiD0n4EdV/9Ua
xiVffwkjurqjxTQRJ198yDNL8YsaGVQJJZdhES1IK3oPwRwqdy68OPOHAzDg56vsGw0A17GPj29j
yiOaQkp8CU/nbbFwoaV2mpacZQDfY0wOY2ScTUW3t66HfCVX9OACdkeMeGRaAzOJgCk6UH+TE2XH
bjCaxkHvQKk5lFOfTCw6FIpLSbtNqIqwxshcIiFXeuV+1YSdOI3yby3MRK9mLdt04miUqyffdK+L
v0MY6S8EOjrTMYjGdCMFxjAuCmzp7/KGJpFeeMqe+9/j2hLvK3ffo0MU3cpsqYlU+JrjkV2mUp/n
GOfP3pTj6ias636lEOXTkxNlxeoxOGnH76vqaBeZWGCUjpycjHp5QdCacW7pqnCIhYtj89XQrBIu
jEaNnIno/kfzgkG0vh9NQYq7nZRPyVUTthQaqAV78Vj57SiBV2JD2CU4umtBiEL3gsSb8G5G/86J
JVpAwdc/dGcPj18N1ThRvABdAPlCoJjniwBEafpelFlDP3aaZgh1LIXkNkpEgLBY1Gc5jGtcWCEd
t7s7r4CDzenB0XfSYVWrpxs1Y+aYS2Jp0+22T7ss450MYQF3NKjBWy1SqU5iKJLmLST+P3btkczW
OYGolDe51ocf7/plOlYaJBgfGAMBlDpIjhKVYqmn6XGU1tjT4R4BM/7J1n+qWpW5GDe6FpOpYYaO
sBuPZXoy/lC3I3a7sl/kmbIZ16pFKB5z88rU4ui++/C/ZZKST/aDspy2sIvXzHeGh5vk/x3bZYee
iocEdlSnWoHIZlYno8UHIbcbV9/Itok1hP0KXChqMN1WiDk6qS7GoSSENk5343h1QKyAvuq/Dgoq
eNNeZu0HD1mfxwD0437TAslegMs/jdiPo9OIULYstdEjGXgFwYvhhsXsd2Irq9uKiRLCUUsgPh3F
uaZzLU07L3gxneuPjiYAX7ZsmsWUl/tWFlJCLYe2qg1jI6qy8e8shZYi1Hmq9ntOSrifchThdjXJ
T3g1uAYG8KQJQ9v/iXSi1YStm9TkoTBhgd3bm/ld1qblJ94vijCY7PZWnRzyQyb4zRF5z1rfYsoD
u1+pPUga+CHlzvn6C/+Z9NKLEQBXy1DNlMB6gLJ5DwTQHEtY3zsIpIwJeg/hh2tJiUL38yhVh/WU
/cePr9ySZ7aQgbtfCxQVjLSjN2VbeQr8odZXsywuyGT4uHcDTEWE3T0vmR9be/yBFTLPuUbe4QBr
JD5vhP6ZxHJpcqnb4X9F/vxSHBsErco6waY00BgDKzCOnxThiAKLtgXNOJrLjV6wRHhYknTDs0AB
Tq69a9jtCp3jhRb7GdrMGQ1H2YYRctvaBuesJax//CiQR7NEuH0l28Rlr+LbbRu8d5ENmHsoHDwz
ynOJUW+dbZyyTkxCGbHJoJmveV0Yn086rL0eHfL2upRnifro28ktXis3OfGsrkU6WFeg/G3C5GN+
2tWOnfwKZ/05PS3X5fOGQwXkYnLdScrVLGUqYRrg5sdZWVqURF1k2npg+vLv7u4OEWhCpEeXinZZ
0iFXLb102bJtlI+YzdCncRE2TRqK5Bc9v0jL0apbAIeGdqC9NR2qsFEs8jQrPevvYYrnL6xG3QBd
CgdADqFGPA5eCdzicFeBu1RXnfYr1PYbunN+/vQXWjwerTPih5k55/4nuAIr1MMT1XdUg+NhcPkq
8vBK1J9weEyGXqja0XZM1ERpu0VibVXJsNwJVa3MPx5TGtVuNQvfBKEXtZG/ZHc75OlEZVPpaMz7
bXd5ui83qsekQ9cRKxGO+7jAr8p8aKEx/ln9AjRUK2UVmSMA9OwnsXw6/1NhHTuj5Z1BQ/1HwR+B
g36TSP9NKi2pa8gRjw2n6VTFkC5b4MbepVr2j3Y+xULQd0t9I/wggu2dAJcjN1xNPXxoOftzEuue
ANvX1f9lJRtj3LrvA1K3O9ONcz83B1FBQIntxyLtwbFuSH+BX1e8cEWICYSdFuPvHgtwUiTGq+ey
vOxZDlfYa7mdJzxzA17ltB5kUx4xzitbV9+jPVDXh7jP2tcVkU8cIlT/ePtoVL/NuBQFIeh8siXa
AxTWA7w9lZjhBrJxQUUwqjrQJCIc/vvVdcYgRtRtZsDA/PBThx07wTtVsz0QkZzPGoi871ye8cMj
HImhZlXoRcYnGAvh4lES+1iG1IkQ8toarigoSUZb9gbZcUXgo3MkRU41hV+Ojt2lAX1wMObFF0kR
Wa0v+IOn6iqQ4TExinv78uSganz+8BNNle8SX8T++E4LssLIEStXEU/djlYNN8zSyXX625btQPyv
hfOi+MtMC4vXavOZ8yNoJPlcKvBUWI1Go32MQPZtLij4818ZiQI2RFnriOXdXyR/LAgYxA6S7CiW
++rsrCjSYBzrKU3rRXjaY21hDnBJV8ZrbnEBi/Ulb9q8HOo+D2mB9r8rdONh0lJF3UGN7BmSFw1f
cQidmjj8VjCAxhc8wGSUKRBSj0wxT0+WUpybQ1Scp21UPtmqTu3OyTyIfn9SeicKR5PSmusOBuzp
7nqrSvxZPm/JOnGLX02hwGYt6GF3xdoU09nRnlb/rzDyNfncc2Xdwm1pC2rtapNCWjD/T7B8CF8s
iRGScJiP3ue74JGPbMViBkaV3+HLiJ+M2Jle69Zc3VKKclOftBrg/PBpsqnlIm3amXUStzZ7ViyT
lM4jsgSXnMlX3Amvw34h1gULz+p0quEuOZI4U5NfRfNrZS5DYU1bDCpWryu4k8OrijzpyEPQkrN4
G27gek1OYczZYa+29PBkNn43NeA46ss2KNeYZHBDesNQkntg3N96UJs9DP3vRoZl8qfSyQtHXLMP
7y59pF0kkSJZ3FKrolsI2pYhgTtsaB1RiZS8Wvb24ogR1IHDxlJpadejtPZub/8N+Yred8zkH6vR
ONiODqxpjm0+G4bwqeXiTZ+CXgEK3xt0O4YLN0y/GzOXRAAsjM/5QqB16s32Pfnlmquuol+/BPj4
m31+Ku+9FdhM89vGshFezbJm7bNHzAZXNfxEf7xNHzdqFM58Gt32T60Z9PhBoXrsgwJsTySDPYF5
5AjevMVt3tkfrMrlVb0UFt6H5kDCntMLRH9cDA8vmNsknJcRALtiGrkz3nNCfiG/Rsbm7HOqsBj6
1o3VWGgCW+KiMxDe6NTk2kF0IWk5aKIxnZC32/ZItqnjAAEQfBM3cdqNnbm1E4YB4M9+xg8fCpka
NtCDXCDnBw9ViAw6zF03uJ0WAaY1PTHdZfb75v4V5ymjtBdewSVgSz13Q3/iMqIfaSl5NHZrzhHW
3jlt7sqdCJUwAf0r7kBOzwosmEa95Iga/fQmCF3Jit1fbAjpPIj+qeD5uglHdzf6elE4OQV+R2Fr
WiNj1JiUwK8P9q7VpDtSa1Vufz6ar2Au7YxRq22q29wNrZYKohoz2P6uH2ppcJ08ZC6LMqOGocPz
3cRsE8Wm39YdW1kXGdKTiCIbwmdOBENClh6eGbj7HBp4wiWBgWtQksFQM2p1wPV6Oev/EkR030pP
zUkDJ0Z/4fFuI5gB03h535LzoDkpOTNKqTj3YCjT5v/FV0SJxb5qjmbFll8nrr+AhH5D9GCwHxm3
UP7NCqcbJEuJYeeSnAos3mmqCEzoH3mj8EtnuZH1enqgAYBFc5h0LtDIXcKfOHDHQAODiz5yXhls
Pil6fE74fzuTP8Mq6GVcqt6A3ohWvhRMnyEululCTdCOamRi6PmnGwBBOsBsEHcYXgBeovZxKWhb
wZ0HEtIV0iyaP0lbtgtYpF9XIGbKW/oyi1MH2YteqLQqmbW51eEh8edp05KYzUg8U6ZoPFc3jhiQ
7p6gUkBJooKVJ6TCyOUYJI4Gg8fPZg4uiUZ3M1OGqff3nyqltD/snzQHtj2gB67jbXp5nwgUjEGb
8rVHV8fCE5N0gIcx7OrpHd9eh7ZfGfWNIeeexMEVeYfhTndTg/dyHrzVY22RVBZokqnSBDeih3UP
LdZbE2qRuPoqgnDJrOadZ28EJ5+FH6zRKtnUPiWZmRwcQs1uMCxKgBQBf47aABkLcROGI2ifb4O/
/0UX6NVPinti/w23eaOb2N9/TA/LS91GNrFRQLTOfG3KF5dD7K4A2kHU1qu6vS8sykCZ/U0rlaqm
ZDQUeKSTL6lEH/Sg6buWUYT9PyfgUGLdAlYIAPMCCb7lQmwyem29AS0Fmi6Irgn6TZ/1Govvl6M9
B47tL6jg40mg40OOEO4SUhO73sH0gC3xyxAYYR06/pu+Hn1WJjdmahnaHAmjfjmd/MvSYv277MAb
E4ioh1yJWcAZrZ+0G6od4zkzx8/Ke5uwD/DIRSWhwIUGDETjhhGJIXb13gpk2C7WwXZFJBWKueJT
LGvlQdBCz9RPfqH0yZ5TFNaQkFYkCG5CyFIXE62DD39NTzu7akiBrnH7o3YfRIEiqmGXb2/1jOQN
wntV4z0ae1reOoTtckRjWwEOAjmLy5ZPcw1gj/2Hi03fjC3J+2peaF4+IFSMHGTprNNZ82cdLrfp
BNtb3O60XD4DSKqX13z2WXxBFO6XDwghck8ypbx+yn78SaaSa/062y+X1R43+++PCAeXbBjmcWsM
M+s1jBW8APCtM8X4TIgK0Yeo63CHDfaoHu7jxlyVeqDvTmQUl/2lLY/Hom7vH1/AYR3weEXL1wji
EpdqdxtbcTqA95CsuHnKJP69JSRyGfvTT2H31Z1JY2HrgEZwSvR/M9euQq0hbYLykQEyzgd872ON
AJg9lc1azLi+8WwmwPaiWO8UW8eOvJjSL4LRXTEK350Ll7MmMBbmgjluWNuxC21ClFoCaR1kryCx
8TZsDRoC3BpCeFDhfvezwydMNdpgo98n7AtoRS9jbkWnCZFZTKNGlk0zwD95kbnf/aRGrnCUVGvg
ZbYW7OkdjrXc56iGmr8rQu2YhZ7uesqOdyD7AruDErmk8M3j/qgF9OHs4WUff/SPSPnwA9PbPoGZ
A8ygk18duEjkKMsemLenFeeUQQvrsuPIA3tq4jKyU3SM14RBxZkLN0cxo1echv8tEmhZ3cTFI/Ck
2YW6Ja0dnUzXH99wyLHOu+r3ykyn4TNg3/GhjyhxC0X8rBtaKmbqIzQSYe1a4ZoGIEcw2t/2PBCW
2rjWl51i5gzkpP+rOv1SqSXo5nybhGUW8Iq/IDKAee4N2DYIjhJnx3haB6QYVLa1Cfwuw52Bo7fI
Gsbg86WMlQ7HzjnmN91XQe/vQb+5uERwI4PVBf5UkbYvRdVsvUgt7bwGY3k3868VcSC0BbSJH5+S
qsbu/GulxBeEghMIeYs8mZn39B09I7lRHCgWt3ceURjaNvbQy2bL8KUocJwUBYL9vsN+nfutSvVg
LB9iTHJ3+DDz0uZHYtYKEjOUgIrxvqKq4wf0hTdeuFouwJ0eF0RfhpD+D+wLaBKpbnADWTVCXAFX
iUElQhC5oAzk1tm7s0oHra5Z4duVarq9IUynpS9h8EtqNR7FxZGjA/wdfI9lyuc2AnNCF2ufoARq
afuDiBr2SA3Z+Hu7rNNvoChod/Q7WP9DVH/oM9VvTcEWknc/2sW7OVNZum+NLyjENaFj9wICHDrv
O014DARJE/vdoWeXIk/8qq2BJVwRkZixae1HAH+7Gov+U9yied1/4hH+t30HznVhG+26GknjFRj6
uoIKuXcoOCnp4r0naOZSdSXMkxz2+/YdhrmYJJ3/Wkku5WOASqYNa6aBGz/3BcULXu+ujmvPAMlm
dUM8aRD+cO0xMOe9Ay1kwYHITJLz4629kHvqPePnkznte1a/YVci0QJfATVrHOqJ6jbavcjSEmXC
27gtPvo4TmuOLeRLrkVf31sQDWrr2KAGO67i7icTCTIMNAMEf+VSo18UI6Ht5cmaonyTg5j+Fy/R
Od1R7bEmWCHxUfnGAJdqc4E1Go156e7mfHam7yAJsLlh9ndmO1ka1VzmgIw2ZbFw3UALuQo8v/0f
eX7XEclc3z7K6I4dIha52KVcPEX25B0dbpszAKzSymJU5nwfYQyEZJQPc7XnEGqMvok/gysjsOr1
8dxPnFMiFUdrBhVKkZW1TIQ+kXWrKQM2zwJ5ZdN+AQn9dOwewPCGRImLJ6zPkoIuJqT9vWqmrolw
mRlH2BxFqMm3z2nZbkDrgnx+3Ec66/Iw4nkX9fKmbzikbu69LkC0FE2BUzrNt/NY2jDarFF6mls8
94TjpcIfQYxMeCGAujzwc7HIhpT7yclC8RdQ7CzjadMhfpjCPuAY1htD6pjMN6sWadqxunu7WCSd
ZuPD1jy6T9I5JMD6dO31skQ9q0O4Tpgz1NLGEgWkLsk2GL15kx8CArwyLyqSZY5WySfhV2d2J7zy
GnDPsm79fFifqQNFqIidpQlHL9+82/gD23RClC5Kd319S3GkR3VlyyWGKMwKRa12D7vrM4NO2uoJ
l8F0l2b09850yn57jcEcOQnDKlrsXWCYIE+jY3o/3TvECPOHqVjXa9K3slBx2zMkpycrBIao/qFm
XGcLofDg9/GUROVIpdj6Lvff/0GR+fWsUluKEmHClLuunZFCq/Mu3DMPl+JhwKjVxewcVGZvzO9F
JZtQAnqcTWTIDo62xFgMxNHdRbEaCM+6JG6t8ghtoeLH6JsQ9lv5HR5UVxueBQ+8TiG9qUSgWV5M
kJCuWu/lF9n0W5X8CVVT75pWzti7ln2LR6GqdYruD84tAOBfOCeP75DegZUGlqVI6VcMr/yG7TX3
QbYRyRhYHQtZAlY5q2pr6TyvB7h2aA/AwdZafUx2iSDibD9nAWeG2RmadKVJCU6tMpna+p2oX0M0
O7LQFF36U0FR7tJDH2thT1AGHxn+PlIkW6G9S2QMNkFLMlKUl/gaJGWOnWdhOaLnfisG011ZKfa5
jv9PKT3N6NVo6mrT9aRrW6e7uDQPXkkCx1fSwXQQtDf9uU/Y8te/yJx94+O8gibcK3Y4UvkB2ylP
YkxNXqM9Hnv7664SHmlHRmUk6y8x22CuDgqQbZg9ONPUpVuXaYue58Zy/wm/lfuiIWDlecJIddr5
2cII4VnXSnDyp6llc/GraZgsXyj8x8t62KqSV6meOV244HSwpfC7vb9HoxRGXWi1MVLvvE51k90f
/XRki6zvY1EUZpHaff/aOWs6QA0c4V0RSEX4kOmoQzoxM8CMpmBz3q/NCmjxcYJUI/+gdFM/cqiq
t+31HCccFpBJZXNxUV9Cxt00rRw9G8esekAhqEU9DoLKlrHcYGHqIL/kh0+q/E0EEGVHuDqUrFu4
NnDOOgo2SqxpPTLaYEDmeav5/nUnvFt/hyaB5Vgml+EF3Tep5sk/5JFFCY3Y43C7ObjDDPPUze3M
AEA2IURl9JhxORI4ZQ/ySri4vfjjmedbQKu/ymkF4MIsAB+9k1VVRsnLOY8sKJEqLG6Ap6QDMTSS
jemlwzCp0Y5/cPt0kVyqlboWQc0OJa1MFplUkPY6nL7K62aOPLn0fXcJwcLeH601EJ4xhy1KEl3l
Z8bwH3av+o8HSOg/CSLNtWianqRGlpwbvp8esspsyO11qRWZNimisdkFtJUJDq74opQuzXUwq2p9
alQCE/oe5S/w4e5X8ec48d0O+FhJcCz3wdtKGWGYhDnvOqDFvLOd9eOjeJP8jZwPGA4ABuqVliPq
voR4KrQyGB0Fmf/y5daQqGHeiPOD4UFYpqt2o5i2yhqaVcvibVeYgPt8Odd+omp84spHaO9CDK6V
ke7THEU2wQAvC5RSfD1lzghqbyLd1DHH/YDTdZS3/5cOxEL8X3FgrJYtrxPjHPyv1WBDg8a9OYJd
mKuSO4CI80VaJnPhXXPUikbkDskcWu0TcJYwgVOuEM7RsApXjcU/mF3xcVH9C1rSJ2HyVP1/1xUJ
9C+M6bm+WSCaLwNqNTWsJMAyCMDAj6WUGJ/kpwpF7BBu8RV+qUPm4+xDH/TFpWU8rAQTGCzOrKAw
t9MtleSkacclqFt0Liswfe1nWhSf7lmcwzggviC3W/zTJNV/vWpHFjwg+RSowpO2fBM/slcINky4
YnJ80VvQzAbeCQd/kYu0St2XOyfyhMXGtBXcCnq96K4oYjwa6XnSBhrWUW95IfZAYLE0KDUey79o
UMNDJdpNQht8Al0xGxApgU9jaFiMsKf2+7LIm+OvwT6SYXkHwN+ARoHsWsfOw673S7F5rU5hysgi
7D6LebsCPRBDOL7Sovp5ZEhT1NUEK348ifiXRMpTZ2UDaI6i+nXFvTWw70NA6LBGv+Y2R89t8XmJ
1kbL4kEXXW6aYMZhVdOmIAJlJ6LTgzQrVYuBMKv4jnA3UBlSASZs6qzQHT3y4NyVKgKNnXWDwPzJ
uuDIv/zgTox3B9IwgcRk8pcTDSsMMxsAmCDesY1o1qi9FwIK3RABgHYve1WoZN01akJoi2mxoBGs
aXhmhTscIHmBC9HWQvxrxtzSK0y9UIpzdqTpCsC3QYEpVVnPDF4k/mTDQizsVCEp35QT2zujSvLl
zVfGRNm3ZAbVdq5wooXweCSVDCAuCSC1aWJ4Xt9tm6J0eMy+Q4F4+cnLj+E66sGXFW8dF7Q3dy+n
2603guzxDgQxWjU8Xv5nrkbQeXvLdQi07boo/GRDHpXhIHkOYRYUED2PvfiCuifhlC9i0GCBVF/e
NC0xNlw4HZhN0KZ27ZT+8pVTRghU1mlQGxDaDxHtqP4WXlxGUniyRoZhkkU1DKqP5GTSdOSsGicy
sIGEhUbXBgxuagCyuvqT3zCXUkJqy3bDlHEl4dMSocqyzaXzho4rC+Nj50yiDgcR4DTEpv9kRt6B
mE+leT14/S338dzRXbyL9XsBETFbkcn1/aoXycg5oEvk7zKdbpkio3fFv3vGCB82MMH7yPeXs973
UoKdQDm2eY4Md5ak7NAPIb9/KUQyPz8gklVhqh3E16g9XMFE3TpNTMDdHEcWU8+I3USQWsD0soAX
/Y2TFGvKcjBe66rKqYK77YZfdd1SM8cw91N8veOTE+Qf1gOG4hSTpB78PaN2WsakBaouUENQ//si
hVHgW2kz+opuDfVh8A3d3JOsSzqgHX/dGNXbNZ7znHwK1Lc0HADB0my6n5ADVS52ZSPzc85PpwlS
vnTlNk3a2pgZkxovW3dfZiz39O/qrAYzpkztIDJgcR9aJ8dxv/VCMad1qG2Jl5DDXmsCqCdZyzhQ
FfMcYnlGD8gKQC5kwttBev+H2TkZ6aFr5iY3WUWc2vbv40nh1XOCTGZY9kmHgMzVxzzPNFlZFv9P
wzVVVxDouMamR1QZLG0M1I9jPgU8NTheCpCDtuAjpEVTbjp29fQwJmBWLDY3SsUXxk4OTPnwlV3x
P79KcbxltljaJCIXnyelkFWwj2lPYkHxNnZOEM5vx66tr3kdxMnW2HqTVaWMm2PCm2Vvdht2KPZ8
cy50I38zFGiTINlfUuJXSBrvq0WxbxJYW4IoiXwp9Con54XBtDCXniYvcj5OmPVBD8IhPTpdKptw
DIXoUYlYU6tK2lnI1GalyWUeitH/MRwVhaPkmc/gDv+0yhzapsMfCJWBGeO8umJzcj6CmwEKNuDy
EVaGKbdC7UIQm9sC1RX7ZXU2Suu2JUJecJ1BH73As4Pzlu4RWF0/Wxr5/rcvVDYMBRQ1UVLA88Kb
N+7PEN8QPTzzyWAiy10SKGxM8u19tkh3f2AcKDnhPQlsCPxLDKE9AN3FjXmdkTDa1BMsA6dFeuJM
WGYR7aD511o///RihCez3HyylGedShB0OxuVCjlh7oWpZ3AK9r3RPMGrPo+QGGO/jZN5X+rgndBb
h/ciWNCa8A8ysIky4e/KqrnU5B5fLWuOrH1WHwbF78RuTHc8dPrJMT9yBvIAPlmz5TflAgVyWdXa
icqoN4EuByYuAO4j2HL7bqoWVMMF9+o/KXDVghsVu2syuAen+jUPzJAihspNoWGTzilkPefOVeD6
FwQoQsa7nIqTAC1jnrVyhQYadhvR5clTCYKTe4D3fA990dGvCgPz8KLxZjR0gJU0grylm9jf3pu+
pZRV1+iHxW1SqqIucrLAqKTRfUqCtTonTaFsHPHKD4GQlw8pXHphj1agRyDXlAsDB2CTFwZPOMOl
OIyWyfPVVIPAEGV4QjYKK6tkz/xk9reGLpROo8AUPJs8BWWW5F+K3XSMh+1NqNFtP6xBxFgp2Die
iSitY1tMOIYlvAs4QGR4q3q1ZavZPI2G+iV0a4+9YZ+i8dh7i2fRwvPaGAl/y456o/l0LpwqvC3G
OjWHblh9R3/JQ1IhDgd9s+8KV6ExlL00whA71TZ1mtT7lYexTBa3oEYjEWPCOeJNmYIK59/LD4CA
HihT1tD++Ku9lGi1q6AitbCELsHPnDYz4JkY+cu1heqOVsak69jMSY5Pemo7dAQrpVuQFB9/aDgi
fyuIFX+TFxg+BmhPfVaVhud66bFPECj0tinxzgOYQXeFnGudcUigh2CYmQuXcuMwBvlha3MRGbE/
HeH4FaKpZeVIJPrK1Xv0BdGH1L+HsW+JrF2EMcEa/G2EsNTrAXNdFHCKNIpYdukuhvIrGoBTQm2g
DdmaBQC1qOCeC1vyeoYOMVBLjcNWGVhxObSDAjAlUy8+CM2nHfI3arlu/ZYiTmyQo21hJT2OETmP
DDB2XnZnZ4JDFm5VAYDw2nKYH6iS3WVggN3skwVlBCL6acP9mZaClJVcbVyVnfZZ4SyATWkCTsf8
CWSlnckc1hGI2ZYe/8pILOZ0mY7eC9dGuhvS2AeFl2aI64RVhNyfu8mX3evyrrixjkMryieCMtSB
6uxRVahmUN+o7TnnBMWrwAdN47hbFUX+DGuTxNYfAUIQiTbizx3uSiKVugNRNKU0IwA4zSRwZLA4
LKeXGUneyg4lx5PUf7lt+2+5PbQrpVOE5nV3P1cfmg/NDgXGjJw2Uxf0ntRzoqu4lXfemCMvaJBZ
+nSF8SLrXRspfdDVAx4tINxL07VoOb+KiWZ2ecNimH4wCuKtLBwTCq7A7H5sGXiwHx0xJKS+RAFG
hb5+IedhlY+wtVvaCgAAkp3w3pwtJZOITcitogyMwEbNUksZ1jLhpoCuQu87A/e56l3MsKZc1uEX
8XIZxhLoW3uYjOQXUPVU0E3HV0nGAUhbjUfBGkCQ5uS9w5p7wIM9Jlzcr9BGQsjjVUQuocB8ybw2
g5bRhlmhPl8mKqhP2xgi6VZdBmNRLQYomO24CsjX+9t96UnoX5O9QDkuoW13Qy/0w1yCAuxHwljG
5UQ0R+O1VGOlGOu0fanZ4l5b6HYJcimjN3FKFbdUXE7al/ayjjFY2sApt35qLjl6AhAVCIn5hhFd
zGg5Ki6HNqHypKY/Fi8hr9t/kd9lzgXOWgERdO8XlRnJAUuQeT0OABoXhWTC4SfmSKc+odcCmzhD
ejbiKn2OqGCGxgvOaUSMlYPlaoDKMNlWCiDy1v+VmwwQSu6OvMolOF9OI+9Q0S4Ke1NHA8rrVWWK
yY1Qx1t5EFzplARjrhVfII9aaSe9wHjtgk4EJnDRrelUoII+QaZ/isc75s6KTI1VwdnZDUODWcfO
sxvNuja/scmgc5rO4hDdeP01yFd0jpxOpxj6YCfhvZ7wRYQigrUes9Zz4tVsPGXW0IkHoYU70mFk
BLE3QaZYL5gFZOJSmJPjGAfpoaCpgJk4CaFZ5YW8ZYj6CwQAS/uDss6mDy+XSBZz9ypjMw5J5/91
nTNBLbkNzhSM1i1M93pazaUaG4MZ652JU2rmHA2jjiZAjtVuvxJ5XUgBlrw8ZJPxqIIySHsckoRn
FOfRzmUPzlNm43RMaQBLihVOiQz9VlikjOsTHEhxX8N4jgQNViN7Q+7S9N/VclzTP4ziP2i4Wg9M
keoeU4PqBkhpeztedSCUHf4rdP/kcD9MsvJFaTPhgu5nbPXCBFpmqp0mlAmgH3iUI7MDPyWeTbI1
aOlEsy0CN0hQ/q6QXZWKofUTNWe5gUk153WIMIJcF6vm30obd2JjAqlVyeEuPCeHnlTbqzS6Vjhi
YY8HuUsjGQb3rJIMUHSsa72o4Qca2NjP3v9nGtbLKaI3Ond9Q5KjwVRaSdty4gI4uC/0W4zeZxKd
55DqCmnOK/CJ0x7kLr0KNBR5VZGyZz2A2uFUlLuVsj626Phm/BwSdA/QfGpsl1r0bSslxwojJ4o2
3c1j4jkMP1Mt5QmeaF6iM34iM8prBhy+QAExo8VVpBRucKdWVDjVUNjo/qS/oSlGLRG+qEVHkvth
eGzBIRUO1oPt4klwKvRCKtesKjU3b5F88kE9ZF1cCfBmc53iPmgco0GDVo7tb92IN8iGzJayCP9N
zQFkC/POUL3cK/0sRz+6uYNNGpA/FtK/ov3qECZtwIxsF7wNcpQ2bmveRyAvfbTi05hc9XgTnciD
Q+17PM+2A+0gbelUA/zADJ0DmLGXPjtGCesNvZ3XBYvnbWVi6hlkm94nXEXAKd1h0g6Gh1pNm9Ly
WCt69VQoKN7KjsYb9rwqFljfwwlr8fzNlOVD7JML1vf/qoC0Dm59xb7Ux6z0eCig93yPmIXYxHuj
lZr9adarh+4IBcOo02LHn/FXvNcc3IUp6Fg2eOywIq3c65ZKBMySVpbBLLqZT9rueIcKg6OI0bsK
8ZMuZrCRlpma58SrCGpXGWccOzksdu6rwt02bsUDrnCKsQdrcXJMJZ3T5b2ghCnNBAICdWXuiAwY
lPIq1tPSXXzTJQZQF07zMtkb0gkj7HFCM7ViLMHWiX1LVGvtExcP5g+6CTiv07hCPwEKOln+qKf+
Mj+sPzi+1HmigIQvvyV+bz718CcgR7UplgIxplMm32CQvAxnwLo/9ouZ5zujSCJmfGVPoSBbOSzl
NF39yaRo3o0gCsrL1WiZN4kM7ujrCioV0V3EoTeEpB/h5ahZI2hdPZg3C1VM4I5L1VCdQU2ve5X+
Axv9DPa1iHsM2RiSe+wTCIAyNQHJ8MKlTYq4H+Zp0PX1dLbnodolt3dY0w+V/zXcTIkhTrS1vW2U
aAVUUMgUpSNDdRWtlZsL9wOr5qtfw2OSImMArA5xJIUlHEgXcIQY+9QLh83HI4Mm9RVWy8l6dE5K
Rst0E0XgDxVFd2DMOjFJ3pAbloXGOL26Pz/hoerywhcru5TtWBUkfTJNyxg7Cszh/vQ3SpdXj9E5
0r4F2xFP1qmyDghMjffJpKrgM3yz6vTRKo78Lf/Ev/8zauqPN8x2S1fVkCtaZ9wNNLjDsW3JTpki
0vuz3DZ38xRTOtmj15xDcDjjWBSy/jZ/f4jvxcohPVgvsAPZMv73z6w/eUI+/0NC8AjQSeaF8ks+
bQ11LQk+xx6ah08nxB/FplIkEhLYw4iMvLz8BtJONTqGU7X+zLcvDLX8RurrYWyGqj1u0EzsWrzf
qKh926Bps41LWaYYKHbp2YJ62CiFF9PThiD8anOWswON2w62FiUyFqGBV0BrQF9lgrZr/ywq+QNW
Rz+BcafGKyDBMhCKlx3F94DmAmAofjpkCR03BfxS6E6Q+6LCxO/yavoHm6RKjriUSi3PIgZPRh7g
tXSAObJs/eW5tQJ0yb4vNiE9Lm9UhPIVYC9oUzJdx+pD72spHnUWWAKhyoG624dmxSJUrb/3TQMZ
C4qzExJh5YaGzQZXeNCSTRCq2NimUvLHg5nGFEFsD6HJhpfi+nnnt4yHObOjZQ+qtMXuYC3ty6Z8
Uy5IQJWBqcxREaaRSQA2zOMgdsKXLmD1NAB6laYDpbnX9rHNHwWR200TQvgFvfU96vWfFVSqu3VW
WBz3cq/VROuXG8VjO+a9YxYBxWcgzc5o3TKoACIWwT5+4iopwJvXxDw1YJkmJnxNB9j/pZuKMYaM
OWMjH7hLkgZl/oA5s4yoSItwxWQGwtdp8zAY71Qgc0l8y8b4abi7Gfefr7JnJEpTZmlZ+IqSVYLY
7EgRAdKZWIEfCZO9h43K9Qq/6kFErsStC6AYtV6aCKcuuD5DhVU+EeltUt6oeTtHZjoeWGLU0qCF
pSIEkGkIIM5bOSbL9FT7S/aMAj6C7sZix6aG95aE7+dnlTa67Fz8Hue6e4XMwzZmlrr+rmZ5SF0g
+9qlKp773lKABQd75aadtPoKOYia9+6DH7gX73evQpi9T70XO8caahZaSPlmkYESYRpzVasedZg/
O6kgzuboB5zFrCfUc3DzGqHS/V2Sif/7epgBs1coLF52D37uRoUL6yW2TR6Dd330qKKw3L1g5mfC
7QhA9PLu4qpYnTCf3H4SC6klzq1N0vgY4qZeM62xSObgIkJEFqMFYr2TjTEj5/yrrBrlCwENWRRz
qmF5jmuJNX84cdRzRLPIVaaeqoEeETceSFyedWdbrhGijt6FwpD1N3u2lQ6/Jg23MoTgs+4rzRde
q0YAemMHTazLWfQXsFkU6OVYUMOvQxMrZ5CjjAolntS4MMPCaFlvtte0X+BMfZmbgYazYL9K43G2
HlyS9wHb/ivplE6+ZSPx/R/MkrFb6s1ueom3Mdi+kYjTVm4NUjNt4AdjTCi0BksCs3X/iNkJw7j1
VI3Lh4SNJ49eiB3QSx8893lrYyPm/E1DBB/kut1jA/6FA7vmXlmNJcGIstNl7PVDREgxsYTE7co+
6yb1stucznglEw7yfMGI7dtLe+LSGnghkkqvWVYb81wP+IZOPhpQl40EsTDTmbOZaUPf6nCVxd4W
8ayqCGnfWRR2wgG3IyImAQ29lDXhdnOVAoC8SYbm88WdmuG3w/HQjVepD33gsK15W0Ir0yWMv/DX
Tg22lvxQe05YKr27+XKgozBxn9EsW8beOabYl9hio0sHWJL7zfTNOZelcOm9j8GEL8okWR3PaBJU
AKIjzraEn/B1ds8LGZ3Ru4tKxjvRDK5ME8SUPo/tc/V9uux9iQyvXq1uQPtD2JBjwPLwBW44JPeN
wbs93YSa3Kn1lFWvFP0Eor7636MeNngZx2BKFHuUvPSC4vffhaZjPkgqd0Ahtv3AVmLiUy4KO/Sp
0gb3UZvVu+3aVmFi7LxYu7Z91tuy8yUPRuuIHgok5m23yTVf6fgieJOWBoitZcwMNikCNCk1xMRy
AFvGsVjkyP/HU/1F3dgVHY5W5gpymVuUvoh7ntGstsFsyCiCHhFBtezyBm/qNHGZ4iiqTsIqys2u
cNKlvDQE5g3HLuSx+os6HMneRHe6GyWFwcALt9XTkyT/cIL7VRygMQWUdBpRFfb6nQ/aX6g2eOO3
meNnUWTzWlqwrfhqwTX+MUMlOgrN8DoKqOU79gIjttF9brQoe7no5J9zfUZGaS2UcBuc+9TY8Jqb
mOizSCg8SuEpFTr4GxXkaqC/4aZbd0pCPPYMvxlW5hnbGQZtOrOehO7E7KepWTJij+LjLqmrefrC
f0+FeN6Ms6dZbTeiqvNHFV5snL8bkEeFBEWCeq/iqh+4SE8NDHtsxpgZXv7hIj5Q4v6CCwvVTrcO
froGJxoLfvGwbvwE6rkLsiQT6x+cEV7tgpdyuBH036jBE/s+ITrxvjmEp7LszxKsS8+x2o9Jfkd8
yiAodSALqHW95A8uWK+2YDPcazC3Kc/Gf70iuZvNNTHGOiKnqjFioEwTmmuP9E8h51mNAzDF5dWy
YRq+dFwKbyFzlkAeaF8ah8gKpL4KQMuRMy649IkTh95iskIajqo2AsTy3jMz6P7EfdDcFpxUVBah
xQcSEwnPMMsTRI+H6fetLtXRA7bOBoYVgv+fns8+xJ1oBx5a/9EzGZI5cW19qQMNZ7GSubIuuLCW
vMoP4w/XsfpUDfjNDNu0m7xK6b1dy/R+Yy7iIZXHN4PptXKSzZqKIgz0ok78jE1K8FyKHxo8opU2
dOJymZk0woXoZQdHtNv9gxuVYKrYKv3TW7tvk01rSqgIJdWE2m82zgdbj2HGlsWDBcSG00Kh/4w+
kts2a+daMRUc6/Rpe7i0EQlAxdMZOyJJShf+osCNOailCsT3QBf3t/5SeQ835dSPxX3IHuuMlfiN
5GZDk0ccwaxWQPph0RzPwoa1eyEp8oQtTj+P2HJMBlvPNa39faC8wMQIY6ZDbWkbNFnl7uUzgdP2
MOGdkG3yZes4XSXzYQSJ06cIzc5/Z7nBS7piatzd73HmW5nrmIP0buTBeHqMPY6vJSku01PEpAWj
QA5hzN2agm81MO93lJAp0uG6RXBw9BjaFoncE8WgBwJhvUbCUZHqquApcUqpQmnR2wezIIngOMLx
P2ctZTI3j8zNb4TxMmkXzrdoqu8BtZ4brvSJqtlI9oTcaOnQlPLWN2uAhv1XC+mXLv2Z17O1XteD
Oz5V7EbBnxdEdJ8KpLpaigzJCfsCAEDBQ2MzH8xuUQzoXi8Tv0Wv3SBFtYHV+KnzyWj3BOWgFSjT
XoOSkTMKwO1GIQ4jfJhPLP2brV4d90j6d1KUKtTZHgShYKPqKz1JZWRfopCB3zwUV1Poe10asMRP
+lR9wvIZANUfqnoUnQtptZBP54aCgFE+DGyfTrSxg2bWafiD/CcllWvZ3bnU+BINysH4lMpyIL9D
Q/UyF6MTdsicdvj6OP+xXFSB4fmfe+4SwMdM+K+QwBr31TsyhLKIKkAMnCQcsGuD1jRBxSaorHwg
hrPZ2KlcCOpDMpoxGr332pFplBet7VAbxSu9jcgkCxUoxYFOhF7vCbWa5LkvUMUMd3lSH0v13K/h
A2CDtxiyh3TKZA1E6UgXs8LUSLHq7KjVvKiNfrnJnEELSHTqPwIk9ngLWrgzjO5RMJxXKLCuW0OR
HcrA5RrG/cvHzGRLvTtrZXIbVNi7RlyWNSstsfcFeKhLmBlSxdSq4fJ40TA7DCwcblcQS7T6f4Lb
A6X99FsX+gnz9WH7KvDy3b9BynfC2nnnQi9Lqkvj+zWBBe/+Tm1e5KTzD1Wu0gLP3scOkwRDZOAq
964XP6Z76SGUi4gqeAeSe2Vm2ECEwOc38T01CpOxUVfAjPOcWIRjPPEX0ArBhX9T+O1e5a4LfKjI
FAwxEkWwKjBLmcM0ImAiFq8kXfH3iqiEiykIYAbW8QgVoNBFOB6d3MYYQ/ZdvDl/22ec6Lnjp3Se
hpG7TdxBsDZ76cGK3yubbF+2tkI72CmNxuMXF1uSmt54WgQ2U2PsQDEC7LdYH4SCwFZsxtZdSW18
T5+bD6cqqMJOC6LKuYDh7wwS1Bx7iaNmMLAQOLeXSopWarmCsANGo1vAJ3ZE1QI8iwfmEGmyDAFw
t0Ha7Q85nWsGVCWXkxsS6/uCQEwywmbLgl6zIYDF5SfTFR1NfR7Fy1hcPP0kJ8JQ6oCtcUWjkcK6
CtWIe6aZ8RJA0ZrXG/kLGEGF0jcakTSxcDCJYAaCZTkuu9pAHA/mJjTAZGDpA8AnTjweL+G96YiN
CS3H8cXYN6YGhM0m5AbB+F7xrTrhCCNJo24uVLYauk5smTt3YT2TUrPrCEun3uZx7KncTh413Ere
Aty1DOd6N2PbU7L6G7WQ7x/n9xjGt8jDgnDWT9O8tKYK9IZN00pV1eQkHqFl1N2a+m7Mh9jjnGf9
dZorastD4+euDrXpPdt6jGuyaqgfDC2Ywffk/1BeXAuRO+dLqGBadMOFH/GZfdaq+yJEuvHpTjwA
EF5D7Ae1Ep913y6/BsRS/wuWo9ScKw0mkHZjo+KlgFbKM4xCWNgtLQA995hGt3PYhBsxoMDUU8er
dws7kFNHMs2n1awX03Z0vpPzf3MZPgvMZUY3x2VzM+/oaUL5jZ3jfAaFDy0lXMHRQfg6o8amOQfx
U5fNIkrWn+3irUvZJQaEneVRzTMAPklyhbyiPuEv3fIPxXM2+Mu8cW1VPdOa/xnPfP3laYSbVmNA
tE04Sa8hTGCXn0i2r/S3fZyEtIQsdE4ldGPDiCpr+9jn2DHh7gQ/Ot+dwI759yatWgsZfsH3syo/
CHrOqoaGbA6eDRMgqVD3TU6jFoFqvOYpoQW7nvNDP2HtjikI/u14WOdps36uk626fW7C61GIG7Sm
36/DZm7guGjaCbj775osZWDKLgngj5HsCPTc4wPM/x7JnI/S5U9DaWXFrZY5dBikeEtG58jfO9/P
ePPaXjxQU8D6oKXJXzBPKfrAUc2CvTL2D86cKP7H2wPvL9yxUFvvoH4Mkbiuh4qOOugC1KrnvQBd
8NjTjDV686y96GEN7SIi5nRUVPscl3LRMt49Sazhoz0uCTz6+WJkQgmohK7ULSGQNCK+q+/3BePO
0nxQbybGZVEyczPnIHpUkMg7sbAslFq+Zuv0Spbh8pJlrabj3pGYzhcelOVnHUp7jU/juTVkTMng
VkCEO7K5A4HODFvD+Y9kcVSgSoJCFyGh92FjTW6pTRyleUnEh3H+lqOhojt6ixvkGy4as3mzMj3x
xZXNQoIcNLrmuz83nCCz0PAP59XjSKRnZEcuu0jKqDZvimxTURzZMsawXuEBAbZpuptoKDxTCTEF
6Yns0Z6zPcGsnHYCNV9z1dPsSpntuHoN2XVToy7Mw0ttQGfeg/uWMEVgx4NXUcYSwpL+L8ee3mTx
gutsYjclvQr9cCts2l2JM33n/kW6Or3/RpHLVH7nahoRhx99F6iaAQB0eacLDoozpxJ1F3aJbciA
Tzr3N2uErYNf0I35SDg0Dud7+LK1wHGU2iT26BUFfQGs/T2aPBkJGg30EF9MNnFlZHZXOgF0c2Pt
Qz55QGWp8Mwxb/i/TRbYy3ATqU6vageiJWh4EV0Aw1IDvXyWAKuzKrMXM13JllsXAH5f+qKJnPsX
CFHaJEF21ff1etx+9eNNmlzZPQhqqsnOWU+bBGZm5GFb4snz9HPzOvkc879f46Ig05g+zcIkezqe
WTDkMAeDnkpcy1e0muARLk8k/pKWrG/FivLO7xxieO5+erHEDQzmADL30DMjjiqnF1/Kqmtue2gl
PQs2vBy8D3161145F9Kj1/BXfhg3PK8a/evOCr+Y+O3KiYC2XJ5Pz5zVaG50Y5rogxlMHQ3qk9Jx
iS7GE/495TXB1I5sOWKd9cRoGXzMisuWZOVO90Jshm5A4NoncWvW/GjgPkRDwT4/gsd353OCbYka
DfKKzOOvJB36S0K4M/2RaSQZsJOJsG/pY39XxS82jsNcvHjBXnhPP/yOZvYT+p/E+haKckSSxWJt
LearExjc5YFi0CKQJ0fkyjees5HvlXrWQynmin+FEaGzGpCCm0z2EexKe6cdciBxMUMZ9L7eZNBE
2rnSqi0j3mXhxaoQx9OFPZgMUfaJqDX4RyXFuPmGsGDzneJHp1vXXd9ZxLauPgG1MgRc0FH/tP1G
ixwoYg4z1JPj1ItiuHo8R5URelkN7jpzj1McD7pSYMwbBkRjDClGVKLkw0QznGmhKaafuAqjv+7T
Zx6p4fnlf/vWPaeioIF6CmwswERXTZEuLWuNhZcp6XOElyw826vr/6K6cvH8D9UWfgJpjicDlFzv
HYdIM36PI1RTBmsgst2xUA5YRsHF9lfNMUlzl1fjrBGwquPjdlCvglInoDcVuiDNBUDHkWyFVFzv
kYFPTGUklxLdECYfvt6chtB/4aHcCD5Ki5ebtzLQKF126bJG8fgWo6WkINalJdfcVq5svsNjVbvc
bZIFLZyvf/B10EDzodE+aqEAQfKXso61beB0iwwk7ojpPYfcscu1Xz06vq0EERFRkmPGEmmPEbc0
cdSZyFxCJHwTP5NPSq0KVoRCFrDKu+2ZvbD7gXplp1hOhWIfw7LJAs4s1FrqzmMxIrhWb+WNe1zF
6bCVP0p+aM1ZOepFb7mU5n2Hk3RvKXKwVydWPIHENJp8khLUtAvgYRsC3zPjdGIUhUZrnBVUKiVf
qvZ/BAZT7/EjT+TQlJPntyqd8wMjXhjmG/IuX0bXOeKWFaTdHYyzBv0FT4IT8xTl8/Gke1KRmZtz
ZCT1wZ+EOAcVqv0PNUyKziFg1JQCPIXD+KG+/F/cbmfb0cfCQ5oZDFUm30sZ0+T0MZTttp4FXNS5
EmtbpHrz2M33dG4LsPbRjF4DFPt/cWmZLQo1XTY9yTHFgewP4LU93R0J8KRR9a1oZlzFLnI7DDHa
ghkDLJv4vdZ6LM/06fVLRIxS59NLRYzFFNKTezXXgX+0My+XmrxD52T21S/VH/7kqMK+FAoMrLCS
uzrq6e1x0xWBoziyTHq/cWOcXD1pYljmnZYXJiZFGgDV5cv4haC7J+WJTZNNcrEp9MMl6UOquk9H
LPwWAU+PNQxHFPwwvo2p0ivuJ4QbWWRJsylTZEj7hykPlTrE9pQIZ0qVlyjut+s0Lv0rwKjd7iw9
S57CfhWbntBWOCyskKfPLLpj1l3TjNxuBuX1BPEAUVw9dAQf550TDtLdT1kBWW1Ymxoky62fjiUA
p6jx8V9oL0NavYAiYmBOfd8tK9rJH2ctZtqBdIiy3ADSFzeOlGhGtD5Z4cWo6BbojPDRpPQ99W5i
S62jpD3L9ZuvBrKljs9qk1H6DcBRlAAlGz9yk+ldKrjVFHHWwClx2UFH95QAPQYBg6S//IR693KZ
StVQ94ru0imu2Yb9Ul5vBAxcqpEsut205zzFoMJ+3BSmloR/dVoARqkfPNbTQGYGYTPsiS5GLas3
B2okpqJMhadbA733HPjOFUjHkWZvNRsoJWVTU659ig511N3oYlTpsy4Z91uIzRScEnFY/qtboYzI
zWr87e2KvusJBZ+Zz5oWC0BshC507pen17cQ5tI0lEXpVzW5FDcs1OlN/XtJcmHAPfG/LA6BpZB6
iKhk1Wu/mg9xBYNHGIY5Ycf44JsdBnELvZoVQmztZPLOYgBACfdbNpvVzhyHu8ytxQ04N/O/zhGc
u8QOuQgJ7a2wGLivQEecuKKLpBOVgtR58HN+WCX+hTA08eOjN7vl2Lu5Ko/f9HEZlNlAXPO8XGJz
0cC1DdsPW2KV9O62+3T3tlZa0/rdHTZsgh9LtEwr3aQr8OrBtrNfzSOzSt17RegoWVDxpTgFSQgc
upxGQaxo28/+8runr9bTEBddfwgtGCqYFbvOrYZ+Sbqjl0m5lCghOWWgyE6rEqVrjZF4jmRWB1ux
x18dYjS/bwOknPqB42KnTByfK15wwHD7Z6RUQjN2DxtFz8Zxlo6rl9OH0S56BqHhDTpBziRqDlsq
XvGspTEAoYs+ncee6SLcIyhnMs4LnetBNjaKV31oeQaHrc9V4ROVm622akpjG6RXhRbwu+CAOouV
UjLuWi03Giz4lFeehnIh8pT13poQejQbymGcZQAtBVD32yRSMKTumvkWZD3b5jdAQMMQYTV9hOSF
k5eNf4MWqLyXVtizc01r3vFOFUWMCqF+hQMO2YAaGrS4qsA3YArpJZEhxqsxyOSRYrtxaeHp1x35
RrvvbAfBVRp5Z4Rym4BGLK+Ddj3rR3qtc7eF2OPR+GuyJamKiUe314SfCCdQQMY/DUd+yXa3/CuC
EKhYWlFdqBI7nFrnB73UwJF6vz4Pr1G1q64HuTzk+YWY1HbuV+FbcxjLIK7LoZmHJ2IdsHI5YUdD
t+SdIHhG4mjf2Z5KGiGu0vHvyc3gPXzQN1eIOG0OwZMWYbvveyiDTr4MiNCG4SHhMhrKHkWW5LPR
TGh0C8UTTslkxhTASAlwvx/3RyghjUf+7dhl/TKXKyo82MK4h0BgS/j28uDVT4fDcGqotp0VamCS
ueaStur8MdzN7aaLraMOPd7NbycpA1VSZjTQBRvbvxcjKmMYdNedJOnADoZU93AluwlX7QL5DyB3
bubYMfYZG8qdabigkRpN8rj7YiDph+mrZyVF3qd0aAmpYHR+xJsJQ+4WOepxOJnJc6i0FH9oDrlk
Y4+5TUdTbX6+ioWh5gxDepQ3UdXoW0VWy8prNp4cCCWaWmsnktx1lmfLk8B82YgBrhNYUkP2jo+Z
eOt5Wue59vSuV8qqS459wFKvrFBW4yGWeLS9AJ8Q5jjRQLCSuXFgq5z8NcZTTX0dPvQy4QLPpeet
Ww7UWJ+U+q8OYsK1JerbiAPiY9okehbhWYpn2ybPX6qGx+60oY68vNsKgypjhVjo5rRfwDlSXQSR
DgT9DIj9NnVRhHyIEIYZyY894F7IwQmwt4XxvL6ro3/An01yofViedhd4gi8snGaVHJBlc5ZfXLK
zOHrNzrqx6HobG1pOcL1dFeQZQo+QiZ+ekXNUpAz3+S9ecn8sEGcPqC++S51ZvvCx2jVluroMGVX
haSO4e5/W7Jalwfxxq310fXrQriWnnkBupkjl/mJikU/ByCf9QcxTtSs+XR8WXgFMSzW4C5+XqGt
47ilTBzR/buDklyKfWz/5d9mHcm6d9waprSehIiylA56E6r8e3ctOytl3V8wwdvhcWKREW9F7xqg
VAqNZg0nZmXHYwCOGEsuf5gH3eVG6gPXmaMcqPBKDaBSYp8HIk6V8Et7I3hna80VSVtTZbIQVJ3d
HjFURZ8eyTHbEVscpEixx/cWR469Bjj28sGchv3bP3SNSOonUTJq5IeAXtmimhcsToAIwPhAsOx1
oLTCWT+TvcKhatX0GjFgECtlKEh2wAblW0FOvwPQ+vuD71LHkMjCgdNSTVst3rGt8Nv7OgBrezcD
Kox3DaRC1Hvx3EsZj79QOwyW/4eAAO9TQkMkk+S9PnJXRbcliQBMTLW7Zod7RYXlDqAe0SwaiuBl
qcGztEq2XFIityT5MdGVz5h6FNgF+PUNH9mIxeRObdic4iXVidy/HcDZX/4AJCFVpddN8p3hlAVL
r83ZZa3oqyEuffwSERkgIzN5205bwPD3e7D01QOLtTS+X4tZaSR6fPZRcESJ26ly7kmIyDC3s+JX
HhxPtWTX4oSLP+4aheBXGILOq1V5g1O1nS1qcx69anJiXL0PRccD52zKgVIAVgQ3qytRBgWcRBv7
m20kQPcpcYiVJMkFOiJdScB1p9Jq2xi138NGcsGvQoodmZyVd7XBR2WPWn+oVXOZvSW2hqj6/klR
WWsBKnNM+P1tPvAH3vhfxCNxeapwuQmEULEiTvHgmXABsGFcp2Esz8GqDL8P9ju9dogTBE2aT+wC
oGWEZV6rlVXyGOc24NexKu4igNxJGca/t6/EBDB/0EvEePfQbI2fLM10cRTdcAwI0kdqYS2WEJtG
kT3kAz2CKyPzZmvZ/QmnjTzWUeKPyHTBdfa6hO8vyBXnCjQxSGZlJrON4tPbfurl4MyvVVRiYuAF
LCdBEJ4xYiBiODqWh4P+HdPuOYfruUc9xt3HtS2+vcBX0dFYFRqQQef0EI4XlL4CZ6jJXCrAkUFP
cXUSMbwjTyHlnYGy/sgzQyU+KFg7ZKgLcv/k2MffsgNDakoQ3nfwkXGj3iEZNQLLFGEN+H563/0w
2cUbXdWoO6u9bIIuXUbLMa8VPgU3twHEpWGjV9bRf6MlyuZ40jmL4f1aPATTtL31hMYOt5eXvu5r
YLvbRDebTWexq0EUHL8ysDp8yLJ5VUfF/0y0rxdRRnBFBHDGChsCVnf68C2xwd1WYg/zvnN4ty9g
USKpQXni4xxBaH+RsdP8uacd1/wFFGnwiYdknwJnrM/l63ye4EO5Y2W3a26UgZYPPhCaopdiSXP6
htrwcZoWt9f8y6x7m/SSJNPGeitO580SB55IpwP/SBikqL9eTw1uJJVWHw0/DBku4rNnTZ6+96mH
aTb5eYwlfLHymVuh96v2sRM/xWnCSlLnWKHaRv71YZqaiO5eVE0TF3jqEX/MmQgvYbrhjQYIKywU
pMt8FdDnx9W5mhTm1gFZCoAVZWwr2vYtlwYmR1EsksIxiJlPHWB5cXN6ZXC+l+Z8cOm+rXgkJkKc
kaYBh5HuWaBbdBK0r4vO8c/opsISIHG2KJm2qnSiGJZaVs7YpJ/vfImobtTjyVEGUdD6JRjCcohm
+3op7JJNrdU/ScFN48ltVIrkawSPShq16n7c1bq4dgLAtv0XKq2YocoPLJ7azdgDAvBXgPFf+Vmc
QzC/GJVFbQoOCjHTNLPb0sZNV4WrqNl11CIW5jg0WrJ4ABqsfG8qJf2bUvvtIOIiYynmte1JlGIE
m+WpuorXr+EFKzYPfF+9K4BFgDXvmI7x9N09OoME8hDTOJuard/M4P1yv1b4uDdQr9GIsf3bY77q
NciMZx7bkZt6GyZH4hzCGNvU2tXaWDEtQIUmX7Q/1doyHaVpACdXznL5YkNmnnPvfcshSbxUqcrX
a9UaA5AHAUQA2wvqFvRQIpGToC/AHqJENdE+aAjUIHMGuwv4XfJK8ahG3Xa3zjaw/J7GTI/wR0wc
jca2TJAVhKGbl/I/Z7zmek6CtOyBPfxDnDda0tg9xuT2CZ1ptO51QllnuLDT/Z6RP+axlLw5ua5R
qW1E0GqOi6j1uN6wdoezHzxEq1Fs2SX42rVvUEG+kBo/Ff+13NwJwVw43b+4RX9Wj6kNnQwx5PwG
iftJPz1uhoAVArsBTGlZQc23q/6DvawVJZMCm3fgKiDZN4ODOuiFar3KrvXacSPebQ0gCRhbtavb
J+rg8BP9tjDcvS9SMyM6WMP53xSd9YKqw1yQ4qK9c4uS/3SbbYAXWEB8c30+ZGdMcRUTcP3/kbxH
efjfwYPKNHDWWcO0Gr9xInBdTpeiLnGbaOx5YyUBS+WohE97vNd3uMQHQBpbC3yQpecgWB0gUuew
mTfLrPqrfBXx+iwQhx799CAtOjILzGB6W1JXYi0NN6eK1FWTLJImHRBQsByVyN1WXcVVMWrIJTjW
tQA/sI1MDgPeR9kuLJSanyfVP05grppvAxh7dRVBw4ta9tz2qoBH/AHQmikb413KKaWM5Ykq57JK
hMZrVY2olnQamsL/o3H44GWNYRPduMfmwTpyufkmi/sfCVTtzMbhCFrpDJnfgw9Xb3FtPUR0ZdMd
Fg/oAMHc5+TjAG+0dA9ZJ3Ey1AA6P9VM8G9mYWGH3z40z0TIjcj+OOQPwokhs1/ezAj9sfN1V9Qt
8TN/yy3fxBcrSymw4tDjUqlrhshIUlDVkvawbFuVIMaC0AdKDAm/Z6dERBqHIZws5aC/sX74xZCc
nDv447bh4ShEM1EwOuMmtNiIB/F+bPIXTPKW6TeZNIp8wY51yskeAYhJ79AksCM7/IMbzdURrIxh
U+wHVMsi7bY3NK+MHMXofXvM4tbKalsQ1mnXDXHdl2PwqkQUORBCawinyYJMvZ1GtBvgKLNepo61
/Fm5W8bQZ5KqWuzSTPqvnMge1ehHot1+8WZJLdze37vol4RNeyHLzkUXxpkRIPdO2fIlQqnIl+a4
3pjyGfeYs6iYyy3wzItsYk0VcuvaIhfGus/eP8vfYuu+kKVMNvVaXcaf3HuHkMLXnW/3ZK0gD7xP
8/JLlmI+52lUsEKtOZcxPA09lhGhYDHAfUd6Pl+6eQ/1bSifcWJmoDvnvI7Qt0Wu+8tyJq1691oT
pRSDrnr/F5nK/j/lcCYxf3mWcTxrUZXhuS9Zg5C1bcHhB0OBMOLtoeBpFhGzhYllo9h0Hswq1eSf
fjag8wD2ComFuRzo+c7hm5rLm1yWIWYwKTnhWZ4Y41cwIFkrUqcArcJdOqIbgBTCxvVgc33Bq3V2
3mY1JklMffbG9mZE6aSaBTmQCebaM8+SrS0gdMTEeg8USHrwf7VWI6KeekuezSXFZEuMRrh+wc9b
q1QsH/6JyZeBIW+QhbZsUntX7VRpjmYzOwIVux81Wlf+ZMn/XhA7YlaVvE3NS4xvsQNuE6LLTAeC
8jBTHg9GO+hGJ13+ZJJns/x3LnyLVqx70eY/LbJ8VSHSFKrhPcfUTWfJVV5XF3lr8tIavkJx4vvF
uVuUhduRw88UxAOw5wIqtEHbBJX3OOdPiZ9HQyTXRChs3tPK9o2QfSvqcevrJVpK1j/7lEv0ekCr
8Iw2te59cWzDIKhDzDnYpTaPMSOjzhi4v61fqjTRNJkAaKe3SI/EhLDmOcnUP6g0fSF5DxBX1uTX
HnL8YADUVCt+wbOfJ+esOndoeM4UMCq/tVHQE7+GqJyfzFepjQlSGTbQvybIDPoVRfR6B4Gld3H+
5Gznd0cOoys1YpN8Z7BT6/FLNEibusxpVqIUhBC2Tpvc/49ZWTlgkxhOvqxEGz3+R2p8pOuqGXwG
KKS5w9hGRFyFMKXxwtGaWPnQcuWav1+WTQNM1dvFGfYiXF+2sxHjuMtBp1CCkO7Vy1gmc8hTXaYH
NR2xRfcHLSTCrIkIiCCGvXdAbaEhJ/MOjCKffcf51OZMZeK6HSW5SbZxRn7/EbKB1DydyJy4/xmQ
HjI3G9frFhopNJgI2F4zqL/jGiA/DSIGR7iUJXA9X/WFDYwaAStWhXGfwMOifRlnY77h+PJCgeOT
yqOAr0vxe6gLyFFG9kRE5eYz0WCHZq34BWnqLQG8jNmse0mpoqX5X612wYElBFW2enTddkzQ4vVY
gAG9QpMcH7D163yP/Pv+ucvcaopGFjACqq0DZpUhMvX1UygNPxOUDKpXxnlAEAkGjxlxiQfoFPs3
L/aDxifTmNlqXG0sgWLAwL3e6VB4K3K3aYCHpXyOECpaOFYCGf8iUZ6cfEnXWdPnm/9FsKB1CxJn
gMY5VzPWoqO/rcdD/EXBdEqwlfO+kZE5VWwaW85G+HmhY79n4Qe6Tk7y3QQAGcpq7laPfqhWBGFu
WgmVM1zbMk2lNxsTp7xFHYvNv7vlQ4sGWy+40rE5ZMkmsW7t6YQKzMSr2C+Xdtu9W9qQhbsoxX2r
4oB6r9Co6/R2bzg8G8bY60LNvOWsHoN6rhP8Y2e0jiKAmeNUTGkRrxM2NkPHfhI03S6JzThCRBXY
/zsGRqgHWaA63EM4At0ClZyH9YdlIEymmzHqhQo1o3Ivca8yhzsngjPJYY6e1nXPwC0gQZ/5L8CU
MaZ1jpMMWpT0Aj/uittRi19q22c4NnbMpqAckYVe51NKhudn62vW9m1Ac6LV93iN9kSk+/rvIYdb
S3lG0l6T3lmgAvcay5F9tmdhyU+FHm0PUuDHolFPZVZ6XUn9dALqr/7XfkfjqkiCjIRvaY3V58Qa
oPROQtEWGbZgwFqzNLP+1nCTf2+qcMJhYuXNzqgUIpSu5xnmyVZe24vaJU6dvXFzeo74KhQJxeSh
7akJZP0ZLfZWt82zxL/V2pAolWI7ldOeu8Q6AUGbOSb7vm6lxHhjkqrQyi087e1fTjgkQwqI/6X1
X13O+GzyKY4xBCySxagUHhuDWteZtiZ3zIexrcx5gmLktA1Lu12eaUfIdVuoKenPiAPOVldOXmAy
H7t3Kp7zLPAzDgmtWiyyKDnt87ZCZrLpmN6CMt8Velgev8JJM3DA1ePL3t5mIedjAzb+ACodn2ga
rVrW5x5BpS8OOwFS92pZtmpxzEfJhXBBYJDwzCIvzhBhQotxuUb4aP+Q3ydRSY6Q/KmoKD3yH7VL
FlBdqiC7GvTkKLky7smVRxLLr34Rv1wTG7CA7M6r4P39BPN0cdboY4kuyuCiDgehlKIEYJmwRo5+
5sw/q/SYZhiEEk+k4YYI7agMaPv8hYCo1qYO6JRTYRLczLyHTWw2DREDDVGjaNSLzNXX92gqL+C5
tBJbH2To7FytURZPi6AsVIMyPIIo5Gbw4lVb6EAxg8EaTc2KeMVj+VfVSjQLfKiwFVy7I5C5/S4S
zD3jlafVazIX4cPFVLqxXMi6mrL0iP8ii9aABTwDaylsBV7TdVXdhkPc2oQ0oY2ERNiDeYJMixj7
AMwuMeo7gJ7Omvm9e2ZKmtQregIeOVH7ZUmt7t0bfZ1BCntkWq4ivXxPr31qG9Waim1Kci5cd6JM
vQhmNlK1rFl2NehtJ6EWzoLr2X+X55I06muuTeDNK23l9DlJjtQuIaHHqlNwLguH5FglT7nEgFcc
eocIXv/8Z03nIss5CxiOg6j+2iyWiQX0j0bU8zw/dab4fXzs6oS57HyFPW7uO9zoEXenA8iOwT4w
Jiy0KjHs7j2tlEA8HLl1sln+lXqMKGoTFIdDd4IWbA336bMENaJvdTbQBtKhPyIuPZgMp9BmbTyv
OvND5vcj3ilSSeRpgWcFx5Z2FFcYsfcKG1iCrBVTRozcHnbNGdAEVx4TVCtwc0Lv3O4Tv8kq7Bpj
RvxYte7kH+E9EJNZle5Iuq5PQ9HJ7guFDVGI3GCmTcTtd9mHduxsC1MFYJfL6pIKPYm6MdttAxz1
Zl2OzrxJafr5uJ3qBo5ERnb8E+bsfONPWe9T/0shWtCFFqWIzrhsKkrAhJQKMh7S/u0/+u3lj3oG
0eqoeA175Lg0EU/Xg/31pO7qaovTyuj+C2cIOrju2BMtmTaOARfSQ0yvkxbHONBLWvaPk/0885c/
PAT6ji8IzYGiuR+C8rEX9ap9M7QzqIMAfKfZ1bhcVIohgcuTTAvE5SrwN6DopARNrvNgocp7P/ZU
GNUsBpW93Ho4RJkkp4HIPjvdnSh8MN43OuxFGkhFElJVCAhDELj4HSIc+gqBZC6weYpJgf4QS2v8
S7HWOFW+xsHL01koy+q9obnpsWeXV5qRPXMRfFepcaOvuI6lQqy1UFttJ2Vckak9PjMq5A7g3pTD
y07/jkiq1+e/tTWWxhIvVS102fTXUQGtFPrXds7Tp/+CCZtvWx2yOmNtWASwXqV+cfy7Un05jnmQ
dr+pe6Ax3A+vhMxWGLb2MpzSJSnvdvhxWanLK1qlGQqZLmLiiirPfWE+bSuHvpBS0JfVrBYHwPS4
XGA6rniagu0JPb9C8qb/5RYV9uWi+4PqmdYezXXAaeXEgE+ZRGX0ODmrd7nOk3AhUTN92B4+amdz
ghPxedLSMQEsGgObA0p9H0DbeH/e0HZXuqXakZJ1ApQZoKv60UyWSngGpLUQvKktuEmZhGyoGlJb
k4tdlhB/3PRRb/4fCJ5v3/D8N/9KyQTLZ3bxLXD0f0JL/wPqDrKCYkfl4FjvrGDW0grNhimii9DR
03L7zPU2KhBNVt3jHdrymoydt9v5JbGEb3nG9eBMmZBcIdCjrcQYuf0zOEu768vmHU+4nxlHtkMc
kuA9LVaMXXMamI+1jGwzPenomf2Am2WD+KdqB8GrWX2Yu3ksr/jMEqqRVkC5gz5dYKuzAZk7JNtA
Fp10nByLUHS+1zydrSdQIF3N+tjGLAOKtb6qKStzB5oM4DuHIwHLiaw9riWbnOLDtWR8UxPDDNeR
+l2et9lL1IXLnsAuZotpkQJfFdgr7/tSg/+Z9d2cCQqFrwE9dkVbmhan60jFjxHu7WCqWjf7s73E
msAAiqLKgFTbhnicJwZZSB0MXLAY7tIqMKz4AH5KVvec5IUIG+na7WGJ4Swdmedmlk+trkYfTUo9
ygKQSNqU259GOT2aCbGDPL9i//KS5jBPFnNLcy8Y/iy6756GQZU9nbdW8DB2HA3xHnw5fOxlH2Vf
nGbUZdM82KZv8pajDbMVXwYag5coczmzcfG8ncsIKCxQj7rVHH/ZlrDKzmWnUjnzRrh5f50aXUTF
u/BglslR5B6b5UXQhqZE/mpks4HlEBp/XUOvbC32YWXDxHMk6J1HADQLdKyp1fvrrOJ3L792ECwy
Ro3R/xCfb02xymqP5cbJw38cD4A4g+87HGXTCj363KUG+URgQZ/dJ0slrj80I6/QcvVvPfyfbFip
uZyTi0qbRepQ9nD+cJbZTwGRCavE49W68GdwZ2+ReGETdMf45Hp5XIJdKpJ7kP42Q8zetI3Uy/RL
sq90yAbJf6kMzvWsqo9N5w8ogysNeXcNeIZJTgTY4LLp6gTufFvMKJImw7G894TLr/dwDSfaQgk6
ojOBzEVYXAXnwXvfum/M0Djbu2EyWiQ0It9bz2KK3wIrKCC+bIuZkiJeKHYxaK9Q9y6BuCPzS3A1
gefP622ApjjT/zDn+XQZdJ+drTZLezB/7DHm2x1n7KkoeVe8ff70eUe0MnDj+keAXsgilq6pigMF
rGhy0wsSjLhOUiZ7CoWKXDsV+rTWMdsvmiDszqp3KjyVC9rZ9gYQ1vX5ShXbbwOrIBR6ubEjRUqO
K5ryoDE1nQ9vNAAgzKnM9pb1UyJUOTARZP8DncX14u2lOHkZOg1nHB6dUDuPkFTO6H0/jnakVPN6
EK/vOeaqg3KZqwrSKfNuRu7F9UOI2dhEN7/F4su2zpZ8YTDgIfnbTAOmn9L66I5jc4X8OHZPt1Ba
4mPqKLXI1PUW9bqGvcaLMHbG5kcmOB60TRdOzSp5PygMCVjnRBP0YuLuCAimxWQCG9sjWwBNMiCb
dyUBZ5UzH+TM8GQob2Y0WZao7/ICTTilR77RHUAnsjrvsYWPWDvUztV7SkokyjRkIiu5bVWhCGZ4
dVy6GX23l3S2m5Jcar7KbPvCrUjzWbW19xBuXhiFbz9OhzuPx7Xfv597nUHNumdXoZw02Q5CfU1z
x4n6jwlVglwoGSJgvLv8JJom1vNTWoYG8AFUDNu87l3St1LVt20V/Ke4MsIAflgPvA3p8RA72Bwk
Cjy5pj62QoV2x+pdNezGceREaJzMjfGE+A95ed3Uxk797tFY+/2wclRcuIIi5tEkFPsrPWnJVsCO
pvyxuJZhRbDlCt+63xsbGKyKT7KNrqpcJ9qyulB1qqjakhDBf2DPV8d7dhSQe1coFQTDO6nGEqur
69kDxovHI2uXL4Y5qVdDIwhlSUyTzS57ARwKptVnUrtjJoBkwHPsAUyJbjeW3pHpr82DTblD7sUt
g07ZC6+FWI+CXQB3UZc7n9FGKq0l3GtdUUIyAv0rJL4/Z/g5NoZOrRr9eI0UX3+brc7giKmlxqxQ
43zSPTicO+u5Am4wmjq4EIMpfNu7KTm8rgnpWMsFhydS8EaAFfWo56DMn2pK0tNhzqdDJE65rZeS
avmoR8g8fNG0AbY7G4dB3u3cAfVkZMlGn02YxiVUQIXTMPyBMdngR3pPLFt6R1/hkvDkCSNCHN5x
WevDwZjCLa8D0cxlx73bzOcXKRUtJcEbp66+RcyBkio3KNjCrlNOTM8mWTs/nnHOxwjt3TE9UAMB
z4wLjWNR4iKTbV6KkJBrv01qWygKVca4kwDlhHeVgijWFncYsRsuFBG2DQMGmjxpog3HFntBRLvb
Bv5GgwR9cL9BdxBeWPptfvQvQSBhFWOTVMUaqamJ71QDSzamI06EsGLQ1ZC4IeaLya8lnFRPKASV
ebrtAnaDoeRCPwMW4PKZuwmjnvXudjxWXU+3kzh06O1pYBi4AcTxFnWNukeZ3DgvznC7EvXtqSUT
5S3gFhB7oKCWMmbMbLTEjGBmjsxstpJ9qHpQq0DcwYfXQwLi8xtT4M5VtsjQHEveLDYr9SeYuGWl
XrZ6ZQt7biV+onIC9BBE2MJ4deVDjApOYIVz8Uk6KTKHAO+qkt43tyilafVKKgB9Ov2nUuJ2TlQF
5H0O7ZuinXXW0KaObl6ofCEKRAFYQKiHoOqoNAFQvmYkapK82jrGFY6byH+F7Jg4vYpSkiJiV2EN
ZNVLja+t3GOKXLieqA66vwqCMJr9eNyO7KlEwniW6i+V5OfOz6nLKK04zJQwk2yrwEtGQ1MVcC9O
fDZwxUHM5Rt0ptalUi5Jf0cryXpQJsQ40TWhmZmnzNcBQnVHEKynOdGUcIBAuRA5wItGbDTuF4g5
gkvZxEzOHzvU9Xq8qCYTMaGGf+OXRZAvRTOrS/XNx6bFPST+sWgJ3nNRJeEGVKiNZqFuBJ8AQ5cE
8slaD7kkjX8fq/9BTv1ZpOWnuvnfH2whsAKgCgv8GIMxM/Y1D5m/tvVV8jQxXa3NbYh/RJ03B/25
DntTeymmZnAy8T4HnM6kTFy0ykwaE15noBj2x89FE4wEAfrMvLd31Qz6eWnV+i/gXbXefN/Ka28z
o90AOYegVAIFvWG2mhOHNeAk7Gw0UytZqQvmLjoMevaNEFHdGDXYhXcCnxcbUZ10LUoqJALYH+oI
pYB44sACavdupFB4u0EJyowEY9OBP0cPy5uTKPNU/rX8m9UEFV66AlzsO1MGXpHohGmehhynkyDT
swsOt9B/xmHb8Gjq+8J5q3UN7t0twXN25M8/NxF96/7J3NaFKGtmr/K7FoebRFCRnr7dl1S7DxD7
fnlJNfomZFie8WhNKc0MhMRwscElxy+v722kYr68gMx73u+d8xo6qVfkkihXixQZv+kMYkApEnP2
g/Fv4G9cYnNVIl8WTYMAdn81F5BUPDObcf51zlbSMnqLjW6DfJUaJ9UZav4H8506n4jzmrGC2yrZ
fv+6eSQobuXZfuo88Lbn0xsEXyahJevgpF332n9++cyY2ono2JWKSSBEVZMGIKD6qG43KL9J3gg6
ckQE3MPtMewltMLmN+2jZ4g7O+/s1YDj1x0amdbQwLFztdK0lXwfi/yh56GgVOMqMopfQEfoCsfo
6lVEn5lBmqgMD0dea6X5Yx+tferoiceRE8Nwu912cAunPy3C3ES5YLIEWi3poFtVOFsXPtqnbMzz
oFXicvSW+PCJM3cnNUhQeWpOf7lzimpHAxhBCbubm05/vKkVW66vQFT6PcHk6qRqOsYkh1bxSmZn
eWGNlkIMqP+xAAa53s2zy3RH+NQYbzfK6guAFytuiSzt7VxcChD01plGUZ63QqMsgc3UB8dNjHSM
KoCFryBwBNelH0hw5EhaHoEE65l9EixEMoB+rBRBGEPkctxcltqvzSGoCEBlcMtO8u3Mrnxq0jnu
/6l6qvQCBJieMbv2CCnKDWL4CA8CyxURg9DGbcFPxonz4/lU5X1+VMaD0iGYOylcKpCeeCD0KWsa
mPaL+z4rJg4CkTXbXGIGKcwyBULn54BH/nrmJ4fNFwoVbcODHJaCQJS2sJSnMaTTvSV5HSSZ95mH
YtMDHAyXDH7dVeLVR6cPZQmYKbsy5T43a5HqrMonZ1pBGUNbV1oGnvOkpUAnG5YyVsa1Sx/LEBFJ
9MUZglHSQkJjsU2tQO2IRI5irKY+BOdQZgkqRoi1C8zb3TQNNrtWAdmzgoFMK0+eILh/n7DEgVyQ
lqMMIwVzyGuC4GpM5rCrlaHknagxtCyWB/gxBhFpA2r8u5vTlmz+Aa7hBHXdlv8Unlb4/etMur9Q
dq8hj9vHZ6Zl3rL0E2wEMKGBQdf5Y5Cbz9lD5CmJSlqFSuHRS47n6yUeiu8GB0wdID0yRwughd/d
y5LomTtXREsp7Vdc2svuDx0qe9mF0zElRMmaKow/eAafzXLQ5moDtsirxjkB3LkRV87RudArarqL
Vay8zAn2TAAqeWXsqivqjExIZ+wZj+u85Cud/xrkgIGGpWUctpKR6wNIO28sgFR2Q6Myb9aAJBxH
NJapIIe2VmKtbWYHppuCWLg3EMPPwMJHHOMUIXuarwktc53Jsk2nAkiDKtagkV/JOefTw3dpc4d9
PEsLIjUP1gnsHDOfa/BNQ6khJRTjROqjxBUk2SsZe2pb13qDDXEwfx2bYkYDOQqURDx1VxB/zETy
3z/MQTfb95qV1Ll7tceUtJxHbF8aLsdYtn6LqIbb7rieu5hmye8YHv6/R+Zn2jG2hMLbURcNwowW
JdbTgAT/xfCFHE59pGCSEGlGBhqeoC8sG8DvjMPOLXNVpLIjOMscrL95v9l8Z5nY8p23p72Q9Xya
JLRCAnwd4XH5In224kA1nr6TiJaYxvHKC11gxVwRO1ELBZgrwNfY0xbruUAvcE32n/1MttSHRVtR
VeI0yLw0hZKOdKYQ/wEetWB3uNpZ32+jXt8Hg8R8a9pqcImaPa1Xt/ygxcBSLmW0boDoAutqC5zt
7m5QTWwAztAhac4tNLv0flIpRYBfI/kQBdpAYJM84M8TEf4r0/afWvBu0iq7i1Alb+RsuJkhJzWw
Kw5dOxlUB1ja9bZ893U7Njg2JVtotDJV+40a4aQoIgflbCBXAtAsd/RAkEpTI0xGteOKhdiUfOLe
qsOyMh3lVJl78UK4ZBHdIWsYw4U94kpO/N+o5XXG311iQr1asrK0KFczcVZKHFJ+NHxY8D9+wTFd
yt0dBW2A6rUU9HDZ9tMGIwnpT04o3fW9RgDdYZCO8inYue8upnmkIGAkScf0zMG3b2W9dQBx78LQ
iSD7r9QWLPD5/kNZO3rqdpzldKYErUkKyqTEKoy1olcJICLpcAvWsetZBeL9o9G5msN8eUTCrKM+
kCgBnuroIX+f6FPfs03qrOe8QVQwVZgiaIC/fq5XzsAH/2ppuQQykycFsp3BfZH2wb+NHY/Zse9r
fWO/nLb/6cmmYY+fVf9TkqkgzCi46aHBy4vvXLXnvZ2nTjXNiHZZqvgw28LprudE3ZrnfdvVGE2w
cysMZkc7rclVIGdXrQdl4TVpADGsadnZzCA4R4O95s9wMcl01MXBx2R5Ty1w5jSKfIYyVIDzf9D8
ik78BoyU/7E9BTDVg4ZLnG/vsb/z7QWl6CncuT6MFs+/RMOMD2Uen1vpZ9X7a1Kd9cES28TXEj6f
v/xwv2a3zQyN9CoiV7L79MF6FTXkF+gAL0ThmdPq8U3HKtSlUIntq6XhCIgylbcziQHIP09lXuWA
3XOUZ2YUhv6t76buVAM+kcYVP3Jna1JxpPWvLf3XC6s0Sao8lGg1YnrVRsOwim8iB/ja6IFhe1rS
cqSkMSo+p+iGHhVlAcGm4JlisfDSUuHDvLNltrBAuoi5ZAML1k/veSiOEYIUa/r+nRkwn0mKAS6v
eC4ITb7xWuvZKXq72+c1GBFLNTXJMF3+ZVgig+PB/fIWim7lXdD87N/+aR2gWliwmzqq27OYacKj
kvK0rqj/wl1Wc2HxNMLWZAtuL4Fc9MsQyTo9xda6Puu2UiguxSx1vhYmrfdfkVlQgyZkmUd7ySxL
/E7/qFp125bWblKZ/bEwV845kZ4EvFBvwlpa7GbYNhAqv7NRUdbY6462tDk/HOIga1nQgFNebViv
Tk8Pw/LZLqXk1h+5NueMpxN3POiaOrC9tELyCvVeqcfTGzN8+B1cVS4+/UR7Rc3ON5fpSZ2US+d5
12WG2CB+NsLm49ftUE8lLySUmqRGJBm1LyRjQhtdGRZvUman+QN5zSXAnxERR6Z7vEvQ0WrYnnZo
oZio5GsG/xoDZ69Iu/uDjiqSIwyD092kZ1mowlyWlblWuHT2CZ/imuIvBp8p0JZw/6npuanVXcK4
lSfDaIWCRMFiqCXf6d7YAIQ7pNf9KvniFMUmCnBVry8KnnSGVu76Pm+SxqciV1AQ48xVAArLPbkH
Q02phUhE8mpg9/g4Ecd7x+h6VrPc35mDGgNeHx8a3JG9JEofitX0k7WlFUPX7FHxhkaPzBpSlpw0
Eab4jNm8Wsgjpy1P0JP9RWt9UwVP1XGMkfIGUHzA9niREkh/zAJuo5D2E2dyKtl/iAhIi8k4yDhV
pwEis6ih3e6EHjrS0URPTXcirJmQbW4/Tg6S7Mo6Zdj5x6CETob5En9d084kFoTq0mZIjrjMPvzb
G1d8h9Y/2ePTB8kdb9I8np1Q3cY6988/HpGG0zcFl4+v/s5DeWusiXO3Eu+tRnSD7bsoHOqdu/wZ
PEpOpjBzXEl62m0K/2qrnNteeqNdjm8aLzBIy6/KdcByuLqZddl+VEX5Nyrx3VNc3kdS1Xo3TzQv
dkaZHhvKcDWJhY0P+l24xNhZHUlxZsCMvQXg5DUqRZSE4RA+Px10xWDjAggK00Ww+iZk1X7oDppV
j3OAelS7idYiQFRPLkTxxEScdDITVeVsRW+TveCusCVIiROBTmDOEC+40XwXgE1LnLUvDBMneW9g
urkPne6tGkr1yiRbRnQGx20xtrM9erNkdJMvyuiG7Mn27jtevPGQyHJuLR8ak+AMxnBOSenon9Jy
705oHwFIDV0KSHbir3UF+efh/+VAb/tBglVo91snrOSBo134eVMdaoqbJ/B4qln4BPRBOJhxTVsh
nt+eJsIwCJ6f6OSqitNZvAMc3/tdXzJ7EIhzek4qdYu57Rb9O63libJuN/eUSNTn0Pi5eLERDmA7
D9K8SdWB0UAbOPUqMEzCTePJjE0F3rfEH+x+Kjas+1IsMWmUCZuR2kSQgablP15jgdsvcBzp63tB
soCHR9CFz+7rLmgkpbRQKABCLSLx6W7FR7KsoE/UYPk7K7Eo1+aPCEcILIwNRqEK2VoR1rpVYNqf
ADCUJXs/Iduw4dfTNEZPqlFOL2aYtZKTHhJMgX/Nn6wTbgJiW7MeKMPnKsuZdwXxsVEwFsre7JY9
kNmqNmOjWukD6HOPzDMR3yo92pUdUWUzeuxi4BR5+eCpTzxyWnwlFaaGe5FhjZgEAxcDU19ATxMj
E6Sn+g6s/LGwCscQT37ZSniHccSUHyHRmtzW7GZDYiutJPtdWUR8e6wAI2RJtNLdak73GOC0iRr8
ZGMrBh6dBkirXV8h65pwCMUFo85Hqd7Z42843xHXYbs+vipN1rV3vnwyyK2NfCdgb306SbEp8VJy
r82XRZGx7vwFNTpOqdKKxBPVzoJ51vm0eHlR0UDXIQZuHUmGV/uzsfm8QBCmMuBIL03W3gQ72Rkl
EEPmjoLQKbZj9jBJaxCHRomrdjYvZbOLyDSE3wPKy0/ulfU+/KBTfYozAQ3h2c/rijfFg4FL488O
KOr2yyFTCoKsc/dZAri0TQ/L/PUp2oM3V8ZzCJexBEY9Py1X8x/mhZUi+6ZkMIOurKCujYAUvCCt
PjVDo6XU/fxL6fdzVs4Ra6Sh8z0xYXUuDHzFW0HemDbwYdNEqJ0rAaQBcMjPd4D/JZZkzcecmnwn
A5Rfy2vpx5W0n3R6JpFjyOSbDI8x6Cy0wZ8uheDNfzliVmaZHVmSeIpv3BRppVkZp8SrWEMW5ZMa
GGbGpgcVZT3jDdC+7TgFWHVPLjJlMVRzcSVMppNkga8mIHdA4nS3qbEbTG46WQKNcSUTmqocKYHG
FhYa3jNjNS2q5ZVC79eA5YJCj1uJwOjBKD8ii8zdkuZhHAsYrStoVHh8WvFNs+P//V6M0pENNKxY
aUCoGyLrMtNTMLWvteKGG4BYxoXbsp/IRHSaBrfsYKeXeavwGhhy/fes+4jSqBZ4NzgkG+sfEKmp
3IaMJYSm5lY+Fy38Sibs2XiyilCqY+e3YZdky6TuEo8rtUnL8/dOdmXEusM2zqK4otwnX+dyooRF
gXq8T7KDQSMt9vvRqSJiXQp2Q9ssqVegT8//wvQYKbPDyp5yC9FDlM7qoFSVC3LkDoZkcIOirFMx
86PmLrpvf0tjLV3Qq79tmGDQaSK1AY95jvJ7Yh81gSb3kkmIdU2V6GQui43fJnjRP1QE4cQvNr/P
bN2czuvf8lZJJFOnVCJpAA+9zyFFAE0nkHY8VQYf3SnY5kKIEKcOgY+sC77+vaFfYXXb5+BOjTTC
JhuQfzOd6uRCsyljugmFjZNOFrnJ+AJ+4YGoO8lrF2s2sOAecN4Byzg/VkoaJpNt2dcM6xpivHcF
QwxCxOfdC78TSQtbfEbKQ+syvES9psGnfc6NVKyXbpKYId40fNC7Q86SSj3nluLZpZpyAr1JK5VH
siGdJ1Uotwui21UofYmDHvzD3lxIsAOs2bmid6ux58rFlswpTWxtGE+fCnj3IxlDWzSzAVri021n
P5PTh/Sx1OoswUVxtS+NB40sXYbIhT/MWijjPmS1ZMtz1TmhhhkMrd5UPTjE9OAKqYSd44BC0N/H
dBjE+QliH+jKvPbqpaf4PpmbssPpyWUqzvap8Iod/4ZxWDAwbdIlbbmVbn9nQTbmB1PFVQ/QrIcx
GUYPDP34s+UnQ93dBTBvWYEGE+QATiI+E7NzDQ6kQPMxJ61vVi2Psuq76XqdRwfPYi67NQZu21uJ
98/jVDt69REFQPaleI+stK2dQRZLTCBHJziLdbRA0Z8pgY2gV0/qwBNWXn18mwY0XkHcGV0HkhTt
YWaajTYsr4UQslA5795UQWkhgulgXDOSThnpO4BNf+V8KYH1/QqCslR6hvPVAe97eXoGYv42Z3Sj
wFr92zQKdWYCLnFmzdtTgV/JF1nxSzK/FNAS4W+FFuKsFcoO3N/DsM7UZjmRnvKbVah0s5ki0usC
jO/Dd0vHFgMQFq6paCc0r9ErFcz1pAW63WHs4HU8iLbJZ350BfU7CMq1IrlGIeA+XIfboFtejwJ7
RoQGJltGlBqkNFnX5+u3Cx31yxYEgp2QWLRm7+totrN+/pL5oiEyGH0XPsymtpZ9TdjYmqzriM1U
G3LTsEv3ghQVA45FjlXMmcWE5uGQWVfVRiU+nMZmirjHp04T2jAaRmI/q+bBDZh8ou1gs040i8KG
0OBLHmXaFcWwdeXoBA+Ap9qfiP6Ig8e0u9aVwn0YQBCbJbP3BoZJp4Ayj5RGo4U2x8xMhSOe6ZP7
Rp3kDMNbG9pjfDyPnezHMgARXrRe/3U3R1YqRu0nbDBsZxDqtyB13TPdhFCv1umVIWvPuK/4Fobz
7b9lsxnLq5hiR5vp2Rk/QQaplt01be4GCSLRgPbRToEdlUBdKFVO4zSSqmoqN1TE3MPwqDJFvzg8
laKGRGemouj6u62RHftMiqBJbDJxwT8Ossusctg1xqNT/ckjlg3Imoao2x8jRykPAf3mfEPTvNgW
7wXrCYN/OWkpzpd+jgd4+lDZJTDW7TDQ7+gn5vJtfhQDQ9syTuNPl8fGPxXlOJSs9xBdPfU1hIYn
H6gOnfdRA5Rsgim8mcsUnWGSrKxbiSHLBsV0SQHj1mMq7cbJnm3YSiLLT/36dLjIoHOV+FjjKMhR
bbk8ZHbSFVcM7nPumTgDCl2saYN1YUbYC1LGZEHbNsTv40oP+WkGyPKxWSYtwj+FCZB1yvRHlCH7
bc/zWc88yl4E5vx2bpx+GsIs0yShE9Kpqwlh6Qe1P1OxGQ0cda7Vqlm7+szENU6BUYh9EF4KV8qJ
BANoZ/7OX21WLuCckM3pZg4XLhZDbWo0WjeuMvSLOZPzdvL/87Se5pR07fngc7gSzu475vvAaCb1
Hp4inWGghwEeQdKPhgjT4atAizCZO7F2HLoV5zszDruw9UkoJOAH3ijAC9p0CnPoQs+iFkfn0wH0
Dc+x0we9sKIwXdsSBKHDxERERAnPvwxiEbs01xEIhMWlasQAF9dFOeVq/Gaqe4FL0h9TSGZvV7zn
MkNWFjuHro+EAaClv1sviZkLrnuap3/GEkR4I/3O9ZyUSLhrb9snKjYkj3VOsTbkmHRV8q+sVGIF
1LfiKVPU5sBpsJLNPe7ZvikdmtHmP3ofhIMj5ImiPZWlaakPUT5FaptIAEAgSD0eczZxBOb3dSIU
i7P0L2meqZVNUI1Xc+RzhkAeHJpOR1sM4ETdnCxXWop/fa6i0k1LIeTkrSaHh0fueZiWEqDc0+Gd
/iW3Fq3Lq4d8KZWbWY1VHQ7+s6ZEjnkBVx/NSLJSwUFur4uVJRQY/5q0JPyr3CGuqOBShNq0SZnT
pu/NktxavlBA2Q0Cud16tYOunDV7LbD2Ne2nVPscbQS4kWwhoU3iIZ3os5PhmXi+dVeUp2KGhfZe
KdjlaxGiQbwVGKaO/inl/etzS25nDhBGfHiQtLaXLOCsVoZQaa3dE0pIP894kUh6rLoBo7U2VSy4
oBuZKrOHvlOIjUQlJN35LLVTLmh82ywgEVeE8+7yC7KcT4rtNDlbGn35F7IcqUiSGAyJ65bOXJGH
HB4eS0Jx9v2oP6Q/rYZcM0l0zws0djZkR2hhXubQqRs2Z0DGqvBXHCchaDfQernfA4MDxZacPjUn
rP+9umJFApI4ti2Ttl01toT50eA0KzTJqnI84rJZCvEinZxiiLY5F1ox1+gOf6KyYUXnLXo01yHx
hfeDCCaVXI9D5DMar+zRPjqftvYNr46L007fB1Zezw59ucQ06xHeYI9KG8+L8qVt3CmJ2NvNz+tm
pKxqVHnXTXvXkIMYZmrOij0aLQwdnyNqXA4GlqsGFvZPLEp87WNHv2XT8wXk7sO7k41wNDNpERY/
YT9giRzD5hrClDcRdePxkAlP9YAvbKLG5I3Kqg350EM2QHQjHNCGVDTJmNOBwC9Syq9LqYWvNwW6
9p0JfquSQBhkeTjE2qgj+/L0u53GBqhKoZ9BLvPgqm/K4WgQ1To7g4ntfmDY+qL9LL8jW6EiKl8T
PAdIYEP4q0mHEshltmBMnVsVYbCwuP4HqjrNfPZWNfquOx5GXA+iEbfhiZ41dPqlGWtJthxKlCwr
EBthasv2RHjR5hHWDvcVFsEEnwL7OcrIuhAPTFiiDOwf3Q0RXcGzR1AjDcs2+EnqN5aVzhTZ34Cy
h2r1RYnPjLq+HqRKQkhIAPGfVv2xzMxMhRA8MnTuYhsm58celF3Xwhc2t4BEEWlia5rgFUOHN6YU
pAocMkiDgwD4xPrBKdR9FVzqFX2F26yYqW1nW7TUIFQlpsuN0V4cW1UEtm97JKf8AdZWZC+caCoh
z9h+nLcQLVWItQo7cLjsGfScDBG25ygP9rpWCssLjPva+4E/nuHLWYYeki6b5VmCYPP7GeDk5lwq
dBS/WlmIYjk2Iui7j7JTnWxgrVA/z1C3m7MRh2YFvS+uHyKuT5lbVVbvgDMhOR8K9B3BWsRw60Td
5qyPgugLJzBBpLuWu/iKiD2CTqEcGjEVIeSs3N4f31n3+ON5o0lM9a17IWu1cY8rYdMHx/0Ujph6
bM0pSY8JCGFReEUMJEqZk5P1omGvazGwSL27EkhtJ0OPh8fGrQbginMYnSRBqvDRbtAW/ydREbSd
RomWgRbWZJ7Zesi18Th6aCVezabwZXp5N8a/Hv8f7MbSwQL67K4IBkMURLuEJDj8LkDU+uN+kjAY
WJHFc5Lkx9iVg00sFJDh+/GyXQGgRjt8M/uBxPS8UZxcMsFBnS2Dl0Cw2QKQQ8TdW5RsaFBqBmRh
f1Bo10JoURLkKOfn3WsR2Zo35HNiNOxkXxsnEGR9sv/ZZUkHdyhpBWyRWpzrHVNQNGG6mEq3PcCS
nZ605vRDEGmkxsQcemSV75Wg5dgodLBKfBg83mE1NGkWLqCZfjc0a2k76qLRDrkwkchiExMowJ75
AWDWsgBLLjn7n0HcqGmU8RMCDGqSJlaGF96NAhLK86Ku4Ti6M+GTVy5qQKkhnSIokEwAoQ0/GPGo
0qexDxLztCOSRqWf8WE37z7Pw+lu3nXCNmeCnqvlXpAL2zvuY8Ii8iFH6rDjaQEm7jl4EC7NsQnY
mJZTAKaXdzdWXgFn/W8QUbywHc2NxQWbIJCRz2uM9ch648Mb6M476O9eKocdkRvxFHy/N7wgoU37
BzFQ+CVH+IyfSaQrV22PmcSh50mvqgL8/R5oMLLVHWuOZqIHTsfpo/yoo5fcvPSGNc2lVh2qsuz2
n1q8a2HCYiTovTrI8y9gAJ2opTtAwtC2V67gUiJVrj995TuerXYtFN9UhCACS1Ftf3qz7kJ/+FPx
qotha6KQwtaZYphJCUVLgBGn/pinWjOAxT399DxRTgUFmRWEegFdhG0Kc3z3f21R7QQdO/EcstEI
WcpjbH1ktlNJZN3pNl8+9a8rKU1cZVfjiXvKycMvHqniy0TCHAzzvPIEtMEhxEQNZMAYlnGE0Xyo
2LFYbxOwi9xfngHJkIG3aWse7vc7cwJuyHQ3xIHl5Pc2z/lOVELSjQVCAV+Yzcyg6ayHLUdISahp
NM4b8GetvyHuzCgSBya4Yx+bNg0JhKPu+ID/mkFn1XV62xobth14HtHWjSe1vhzQ74wI+FDb3s6a
QcDHLLHTXVmyUx0e0+U4GkXwzUBl6NQjkTQ0HcM/wqMlcTDDX/2MCZlyhzyxbOxWoJlrGVCsqkPV
mmqE5Xa0k8Ma7n/znxFO6BKQQ9TeHma3lULYHSw7a3M6FRQDrRqnbl3X8RH9YTxJay8GeseOhiU/
ORKq/hY6I9j6vUByvESja7nZmjGJ6zOatELzQrijEeAcw+lapWuF9eoaq8Ld6q4Z9dxnbxDz7WpG
yp6dzUChYYFOcHP24/KG+jKNdokvkk1xJ/XOdycfELoRSGJm4zq4peyylgdW97pFXO1VM3TuGBUM
Ihr/5MLgwk1YNPOTm0xvi09i1U5QqPNSfZciugcsV4+Lgl1PAK58TB1A84BfEl8OATvdiupQ1uO2
Od5DHN6tUVj5yrlaAx52+UaY9UMpO60KJuB0S7EoYJyIVv6F2P5iRVzYq4TNcoHX9nDEgfOs2OmX
gKo1XqceXZ/O4Re+NT2CiV+lNOabtTzkaMdAKdjwsddue8Lm4d20l7jDRuAfde0p2wf3TTCJQ/h9
LQXV4FGFeqnXEBoizhiLNqb5nLlJGQrsgYy4Ox4IOFEX/D6T7Ayr/yDz00c3jPtv5N/QqIk/DaHH
4UT9LrpfTzlJkVqVj3MrABP9LQ3dLoPpCF8KqYCdULQIaA06maZcQQGT053gkJzJ0Uuc8nB6zlF9
nTgnRkmyOTFt5tSUcR85IDBZsTg9fQfdGjsIl3shibP3sdCRjh4Ji5Gf3M0otXBuTONjHIVNL3om
i1kIk4oBPd431HY+LVAcQw6KdpFWpoJtuCB4fzPSrSw4uRmf0H8U8PfQxyycyVZT8gScOANaacun
R1u9x86K1IdeB2dQ1p+GJJlLrKBQmkDA3GeH8yaLzM6nMw6xpDr2Zs0CU8TQPFBm+IOtHOQF6pcT
KC9+JltFyS0Dhz/lhFB95v/vgdDz4/dgFrSGAy5KXDnB/rCdhxF2inrJ8vCevEofghzK50SisBS5
LoOsPBweU9d8HT93jBdxKZFRlghJCrHYZRCJGq6RBE7zlL4ocBb28uNNWXM8eBb8wy/ZONVTuNfr
TqLH9DBhLIuLheZUPo+QwsL6IzipqbascryAC+0H0OlsO3d/9MpQRDiwIgdMpDFOViXXEBL/w+Z+
KRLcOwomOu6N7bdlwFhEJ6wAgJIXKoLtIn/VKON48eTSQblOsvCY3rjw7Yg0VUJ5YEuHgwpj9VAW
Apmf91BLB0cmFUcTQZY0TrOVg6p/DHYj0manglCYli2C+BA9jILNUg5TGo+A9onD2jysLGBe0kOl
fO0ArC1m1K2Eq9WeR6yhl2D9Eq6Rv2uIaLIl372B6TLWKGZH6HOvXkORyCkB6Jze8x8T9PtWzWF+
XtS4uLIFn0zJDrpQjbxOLhmQ83DWCwqsgeVg2mMyvSYNTw4oZkMjeawQgdCXOmce23v3BaNad0OL
6o4jUNa4dwlVEFnJawKuNtHNyOxb88sz6A4N3oJgsBYqhwYB0WSkHpPmI55IoEYtoLTE4LIQE2dg
vbUSlwWi5ydD4WlXaoEEEzj4OUtw6GFpLKoAZyLpQypKBHc1nVTKPpBMssi0OBdP+HEsc3ixwDN1
8/PJ5Lt2+cnw/GQqgGp2JQ+/09muIWGCFS36rq666azughToIXo+EMz5eq7AUOmK+u9xs+mCs84C
6G0ueMJhd4DdyD59StD0558pA0FwPE9H+0qE20edGaqzPsZhtluJ4SA4eDDJFLxfRPMKA2j2GvrR
OdvWn0acYnQtTrK5nprge2zMTGCC+DOL4V/9EUGcJqHFueH4VZJUjEsg4f7Mw+PDIl7CbjEUCzdR
wL3H7wLLvNj8dnpJ0udQBQAKlRxFQADm7lKcpV1+40brWyGuTQwzxdklO9viY9j8umaAAWvn+k6r
XyWy6s3y2TEQW2Pjub4cJ1L7KOaTLyaPMq78p502QeyQlTPdSjQm7CrfZOhW2vKfprIXDLmIU6Q+
yFciZPBPs9AWY2upj/+tERwghZg39f4ZjHlL/QEnmnhISmS1ukPFlekTsdZZH6LEIit9lxnCcHcv
OwR0bORyLS9+gN/3N6Z+m28fFoh5E56/wMhqpoj39gqjA/+sNBd2kEV19cbXT/dCAM/KDZCFvvWP
wgLXd5DwE/8lJqjeV0UvGDYhRTGNmWd87oZ6cU9FQPSZ8vBs/gvK/hVGJhKVzuP6+WpIEnRMinYl
lGz5LoSxFS3C+JQbOVO5WwBznL7COlfFYEKy9u0jnjcPfQCo3L9X8+F6u/PiMaeaN69FJbulJcQx
ao1x10HLpp/ul2lWzCL7OL/NQW8AJqcNykiWxnBM1Pl5ssUdLfJfU2VQZyRWVdUUehMyHV1m7jDp
y2Q5dtN+yG5CkGNUxtHNliBy+BGRlR10xC8RyNw7zIXiS/gB5y6k0l2vWtrq2SL2rdj202uVsgZJ
TS5UbxyMrqq0yq/FL6xjHVKJscBC9AXxPiME1E3nAyC1KoXoyNtNN0dz4hFU4wjMozfwbsoe90nc
cnuAQx9Ps5+hbiLT6aJwn/OvRFjpliaM/ICPb/iOAzhm36RDgSkxDijbOFaGBcbMk9vpkt5MYb6Y
3BfBUbTUr9YvM2LWvU8yqCScPV7iXxOg4etuOJLBNcXEYPq/0xhbEe58cqi3ZmSSpAytWvl5d4D3
zhgl0geQOpo8XUOkkiW2ms3AGvEn+zI1Hu09cR92HVS8rlkyzwxRfGFCihYMou1LozoRmljKNoc4
iPaNk2a/dRvcSnyak7gBBJXIBztlAg/GMZGgcQBXDmhFdjpvNJBMoz+aGSa+rwroYEtvVDXlgc74
3ioSU2Pf4MaX0Mbw0JtNHtKIQgyrS+ptbmMfajeCOCcpuLYwISYYBC7zkntZCpGvAVaISZrWFbN8
NmjkJWR5LlYJiBR5BGbPJyI72u/R0LPCMjuvfV0vZy5DmdqlDBHGJ424TMCTS4RTupg6VVNJfntF
awdxRprHvqYE/200BEQJNhOiUzt34ztkdREp4gZaooHunGPLlmYjHEn0IUSyP7rX4zZVnMK475TO
VVBcQ0Wf/LAZxemjoHfKDMcVhyzr7XfaBxghUL1VGyDhGzvfDMxk3lxz+JzDY6BjJCKtcdGF/Elk
INj/jrP1UqR76DYxsyRjwjnLYjUvsLjM+G1b9dKCpApk1nkT3H8m9vl40GFoHrvn/9qjV3e4+2yJ
qtqpeskZHK813jwJSR6pTTDzOJxJMZ4aBD3ttpNt+RKDX3FBvAmYsXb1BntgEJh5WVcLzIJLLJWf
2lS38g9Yp5HPEBFqplr55/t/XPQjxl804OBhzsxgqP17RidUiNEN195E1cshjfqoLLcM2hzGCDCw
NbfqRHX8RHTlN1ajjCi7V3xn4u7JftAO4v8kH6rPOQY0dEYzDGJXcbAVbvNKDBy0OCGEc3IvZtL0
IhfpV6ZvVrXiwJmtoEwkk0hcqZD13pmsE9aEOnZa52iUvVIiLeZ1239Xx2KLR9ylIbE37Wku3oC+
rx8KfBWgFFaOWExeArHySvdXL/wtEaYtuTT29XM1jngvbww6jdWYtHxDSMZaSaBdk4S/3P7AintP
NkFaIAfSOuVyBDcL50sm+zNMdCms3QIXHM/O6xoqadIZUEjJBZ12G4f4NrF4Bccjsyw8BbHzd9CI
y73ofJoQLwcj3+WGFeJjgIRYbCif1kvVjcmmKPCJUkMV+6FdaaYJEStNtDw309NNmQMid6Fpj7Ms
acEagn8aF7006GKC60htlizkiOv58uXJh3AIKr2jvqlCONRPZR3A3J9mie43ZzUsNSa6TDNGZqRd
+dVbPSGSfcd47yHxMUFthEP8J8MMVCGNwYi/Eust9dE1eV878IgVAPhymDSvDK8Kh7G9PmyLQ8E6
yDK/IeWdCx9s/fBIbFMfhJ1Rp8mWJEx0zwFGDCpj7bKNyHgZ+5QDxJDztiWj51JgOt6TJrwJ57ap
MZIeNeD8UYU13ALHum1jpHzlhxinfF4j3FDcvBklBo2zzIa/kh95lEfP0tRNWMLPM4AXYqDSNTp6
JrqgRZs0sOLLcN1QO6PtrfN/mrPvKjFsuxK/MM8xJdXUDnR5JhU74JB999651GYRicHD24G0aI4F
4X8fLazwmpzrHdRpK8Xah94ApfUvMEVWA257e0ARhBbilMzgA1b8do8N5X+PtT8SvY8ePxGxuqW/
ovGXfP5VCAqPXoJrypcXKub0kjtH7Rn2IIETkle4kno60CoOYEaKAYZvTi6BxrhI66LcsKSjfHlW
yBOhzmkQVJBlVhA2DQ4E5E1V5Pwc+r8zVahS7XwHBpK9eSbAzkKJ+hJz0S3MHOJ6LxkWInxXN0vZ
jlJNN6xf60HR90PY3hBFZJ3lUVGLllaapaIPq2JNX99jNk4Ndpq5zg9rcKK1RFPikekAt0i0kw3W
+KeNIRFR477qlPihgrCbBXy9t861Y7zmwPVN1/J8iy/5WCII6nPoI4MhmHtzwXVB0vScsR31l8xd
f+JetOyyqvrGxFp4sWQBK6x/b1K5sSaDvp4Qa/vQSSWI3fJ1pQ5/H+fM4W4Fjlz1sxwvbtV8KOw9
gDKxvrCSROazVCdshLTbeWAD6cYIjU2sj84r82CbZ9cWGoF7G01Q2tUdI6HsxKR7q7s312pzINO9
BSR7Pz72eP3CCC/zKUYuvWSx6FBAGt/upDq9K5LKILQ18NC8jrXOD2ck0F3yWXr5TP5/HMzudtnh
JsMjd/ImtyfxN4xH6bsFXdankEi5JfB3Ug3mKwLvwo1+UfHqRyy2ce8Cpbrwl3oxTxXg80ntJ+pp
ort/LqMNqhOAgSc+MQJfpJkON9NjVzie/k4UFdUWAADJBvt1RRdGkY1MnsxlpKEHOH1UAzKvJ67s
kYS5w4hsN5TBwteODZE2s7kXxUeClBzoTK3GC/QPjbTKadH0z1O7Dr/KtcBdp/q+XWToGWPvvhmi
3KIgtX/0KrtUOsvfnHfyFz5Z9wApjYged4PXjaKzUvT2tqiFEM7aWfHOi3VgYA31Nrjc+n+PI/IV
oGVOGIlhFxNsAXb4R0QKynZ8I2ohi3XLdT6rqIsPpdmpCmdPYEio1Px0FhL/lN+KX1QRBQXZZFCv
wpG37Z4szEupVuNGJyheZ1wV4QCD2PCagFGL9LgTX0RkdQdYJbRa3D1Qcfp/7V9uaMCm9GnhMOnP
6naoglm7E1D2vXbBICnaWviHgA+4xTrIQ4rseeh4DksHg3U6O5iu5tgB4pIGRNcx7Gw+KIOJP34S
ve7hEiiX8cRUxDicvt/OzOBRz/2j+TOvrLtr8+ElaUI9aj6HCIvVQlXIPR1SgjIA0Mjr22STpy8Y
2I6RJJvxa2w/fkiZPlStMu2wdATxW8XFtGWjT0QT4Yef1HtS8wZs6PgUU/hjGmhR42xezeqqwnJm
LIqFKzdNNRBCNdlPgBqkwmBoIICQJ8qNOJ40rgUnmbaDPIUPnlfH0ZsIgFvWMW+F+Q4cYXByE3Xx
OIfKSsRKWVRfDWpZDUGcM3gr16jH9gYLnuxIad5imberZXDwngHPDplxaHSBUh1g0ahX7gYuvWJ3
tRwrSf2QRfX5XyZItXdC/f1PNjBGQLo1BNQXIdZpvcXJa8f4y+fx+YhxUrvpahxsFS9D9SmYSztu
fHA/HzqxEjdJaX+jsJ71ylqnHKREsXPdw4vQOeerPvPFgEP8DggIWHeq8bkt+9GZs/UsvA5PJ6Uh
WyV/fxGZvKbp+VnTqXHidFiBd4vbOXSXUCDg2WxstCyNTsKXYmB1C233fT72VovlgzHzQwquov6c
9b4skKsMzHPdtPZlaloqgOuQfyf/CJPFrcYPw+1aF/Kzis4WrKXUGdaxIoL+XOgYWcqPFFDcs4pt
s4hjWWi2B3/5q71cNetnj/47MvG8s9gY4uul95irs85htTK/80tIDi7iUnl/N56mDGhgmU9MszT7
5xKrouWolV9OV9pc2Y4cbytHMuE6QARYzwgx4NIKKSUHCXwnvd5Yy/Gn7ihAd3RKnh7QJJasFl87
90cj2GgU1j5qAWoajgcHcsVLtHChbC9eIu9fEMSD8T9eQwubrPiBusiqAKEA1HGyAno2B6SsxLAZ
mczm0NOi/w1f5HM1kMSYiaialjpFZmwJxE7H7TrR5lOdOQHRzO35XY5mgRfBMuJbS1zbFtJlFtYV
1iwmu4D7QKDYbpehiu1LaulN/5++VcXH+bDZDAs580yBoYbiEx9hQ43cOEjcb827SnUXF4ODRUwu
SbcC8AaChmroZV2Ofq+iMnOoVsytGEYtl7m4HBdgVU7TI+f06K/jCzhS5Qu6PphL83EGJZKMZVyt
qcQVqhksEOukinaD+hqli4JxBk7WbVuXIXq4+tOHhJEAFwIdch7T1rS2eFYvEdWlT948SgC0FFjb
bCT7sZiIGitRjuScfExL6UIKUGvDR2Sj1sPPdy5bbC/IqnHNfrWZU1OlyerqVXPTZF0eDJFlY7NS
1uw9coazVijOQ9Br9KCpDGrppbbKUBbBswQ+T6/vpYMpsJbj6mQZKW6L2ifczaNkX3CELUq3OSVv
th7fFUqAByc8bTn7VEPJXN9mDpO1EoqHriSz6Ce9ttadWjUetG5QDMF0Sdfd7mUwOraDeUjdzZ8D
ajWWOskavpAgK48GZpgnWtccHqfOfsOKq1GVLY5cAmRIJef62ZaeigohLvCZe6Ru3glpQZjOCqcZ
kdaepYMsVitHrEWBgT3sp8EFyBZzhb2OuVEwx0NLJK4K2i2IeM45TB+TQVqnhtyqsXFnAQsluLl0
JZelc4KkTjz047qODEyJMVgNbH56G5Fy5QtBHH57GabQehxIbN6wIXJTQ1v4brWobpHD00c68gL+
rIlu2QkrufImpj8tiLYIEtLX2XJ/RuU9dCvex8mfyKsNOoS+jn2FRqpXu3vQ4E9DcqkI5xm/n0PM
nrasUi5Py+wKPoPpe0sakdiJF3yRf1/C7UQJ8pmvCtpl/8MBdq56bfYKCDPuBX31IJQ1Tlpp8Eyy
fDJcBMQBYP8azti61h+lTO1Pzf6HlebeEAdnKgPNoDLXnDWFuwbfmhQ2BM+dg153f2PuqL7lxoSS
1ZKiD3FDRRBUz5YqQS3vLtnsjHqlI6IHP8qCfCSH8qRWOL9PASsLE5MV6+qaGesCCu8FsuwxU5Pd
VtvwEohJU9be1h4fJBV7l002iMjNEGA4ECOSqv43E5u9dBX4tBELFWRFu55/DwvVVPTDNrsZ6RhB
5eutMlLxdvpCOp+btOFtlPkgLYhAnRMp1yoiNpO+mVMLo5sk4x8DC3oD/qBhfzb041SBhip1soeu
WneEdja0HuccW045zgpzBPal6e9ToMXNSN+OrQmbSmBoNMFlevHqfZkvTQMREHoDMD+QS0xy+WMe
To6tVnf5LFyzCwLtLmpH0hpl2IBG0GqjCzsIer5Aj1MPaZ+tVJsJ04ArXUsgu2928gSwhR7Bwcvo
ZrhM0pjm9FyUSngkH5oOfkTpJS2ujBEz3l4aGpdcNJh7HeGHouYZ1nUMGj1iCT786EL4MmLpVPK8
1MNG7RJvj/9DVNaKeHUFP4a/qR6ZR6XJLwqSkZWFl2V3e1AAbo2VrcA+YidpHhaq/i7D3dr8daQ3
LewmtaYlitJkuucl4+jKhTC5eYmEZmJIGqm6oHSIhyqan0MJx1S09N1eSKLSdiPYB9gX0ZpBckDx
T3viQQNmFRmP07JGo7UOSji/RasJwCIPMwUNoyJAHYl5Epoj7d9jfh3Cs1rEAwRQHMyTyol4V3pW
97fTIvbBejYztMMhSMrYK4D7ikp6NrqxoItYjQC0n0hM/V//eXKVdP/vgYJQ9hA48gJSMBiT1lNJ
D2WDo53gHPeES6Es/LbsloyBqTL4A0YfatFqHWeKl3U0av0U8w2MBetSn7BB0JejIZLzu6p1YOvz
aUZaNKdC1h272+nHhFrXSNF4q+MPxdeLbJeCfc2UJlf+WG5o9eQNe5ApelkcVVf28YvXAv7fT16P
YmmnOFaB1MyAjhrbD3mLeTtw6GloJF64WTVmtz+UgzJ1bBMOP9MA7nEXdN8CZdO1aisoQYuKKZk/
/oj/L1vbAjlmPSWT5zsFeomkk0537aJK8WiuM8/NpJNGbbz1YC7f5O5iDS51qp8gf2JUfaAIwmrb
5n8j6IdBklfbxTbKH5WUpBUU+sNypKM+gUJvrdq1k9S++HO1OSDy2sbWuwxlvOCK8OPEdNF3Txwb
23STgRtcU2Ek5BPfU8QUdtCRzQhYBk53beqMWFiOU63AmgUu7MRzMwrZTOhPFOZtG3yCA03ZeUqq
U+gi0i+5yXGQZBKTSet1zb/ARkmWehKwCakf4yFDlFo1SGNnmtr7LIoYtZHUl1vAXoe77TWtCj5d
UAq3LGDCiN3dvyDPmX6r2mPJ/priRpANQGEMw0tXdIXu2DFLGWEe1skS4z4evqQqKxzwg5Iq/+Zw
ZDpnoX4v2j3tczFreVEeADmOLsQRATKHCpiWa5PDHhM1WKKryaf5GWHmzxoRMp3qReht4VeaU4hr
LuUOFEu0NQgfeRENRt6t6tJDQVIQPER+qf/rv2uhptgSQ2IRrbLeLnf998SaRJmTux82OObxJHT4
ZS4uIj1BbaNw79vtsf5nnJmXyX/OUDU9w0iRfR6RMZ8/5oWaL5LfEnMbouL96CVcqJhWkRcvfAi/
3Bq3w8euJzIzsm8oNd4YTDVNRelZ4NpGtGfUOPLeP9i5Kx07qDNLPDI/N0EQl1hd4GvCfFn9rR8C
heIqLMAohIkuZpoYJ3wNwMZ2bioY+T/KEjgV8VVTgLmUO3MgC7KEFVoazYOZ2TRLLqtLlcZGr5Yb
cxUsOHVcKTIWzRpZf0HibOXoi6AyulY/C9JUGAfc0vwBDz6cWVqUIkrKLGZAWguQhqfRT3Uwmevw
lKXUh4iyMvHqtURkBcISSLPYpmycLUgVOX4rKFr/ss6CFsfOQRXWfeiawvH+ZCs1WZkiKc/GHeyx
Ck4/6AsJU7nZEpsYSxW0gk1/UE6LAZ8R619r7KLlSIf+0m35PknpUANsq0/6BaaJnt2owZlg7JlS
W9zPvLPWjWsUki643DJQu5EyQx0OwCqfJoh+gsufUm04mrV0i0wU3e/H5NWHOTlXDTSBzR5es6Rz
GDplRXPeETOK3NYuko+loB4MpyHXn9taN8E72HEZXyztkKnzDnVGHJ5ObhaidG+8m835/AMXlGr+
3InDJ4bBGSKc1PsmgRoi4+W0sxW9UgGXO6uogzvLFBV1Ifmwo6KDCS4RtthgQSq4roNo5+Q5UMH2
NzBsmPjKYTmaQoinmAc99Xa8dBoFcHeVaZNUMkABS9bONVvhac2Pj7qfMuNcpUYizztqRYNnrBoP
dVjKGMKBuHlj9orr4BxyiQFJzuEpUBTVwFuvjjC+/hIzSfc8RDmIQaUzKaviBvzVqn6ZxiCQpPru
1DS59Hm5me9Vo/0oIiJhATcUa8SkB+LRl7rmIB8vkldKQ6w62Syg2XkGeg7+3YA6jdU6jnDkrIAG
irzhhwyCbcJqqcQ5j5Bh4PFQCzRMEHNlwpmAuxAEjCgBAw+00qn7eLs8Qyjlds+6IRuPOGXiy1Jl
xh8QtsXc2FfzX3a5RdAiAgWkKJPxwHCv6w7vWiXj20yNW9mqoHjOe9tZRtEa9jqWyrkFNOeo7VEK
3m6g/Sw6xin9PSzkEU5RVxGrqLMghSGeY0gg3FdwNhoAMHKOwI7ZD8UdeQ2ItJF50pHFa8kXILz3
NdrS09TOsR5D09VsYFmrAX2XINwKPxPH5cccCg7PX/TZoQzTrpXOPEMDK/rYobP2hXaZdUKNstf/
DHXEPLucXdlJyB4z2VeTVr5zbzV7TTfwYfdp6s+prjHrvwG+RVw0wGnZq+Kl0sDomfMywGo0kzQJ
wXWHLpFWu1w8Dq+dImnTDfiTQNXYF47mNPmyOx1oPw7reej5gZsr7xOvjqf4PL40geQJht7e//zX
c4tgtu1KCKHZBMDFYfYZXyfsOZ3NggneifdZNVzu/D3GY+5KQQA3tkQ3GF5vQfKB8O355FVH8uRK
UzLhtpp83PnP4MprK2arT7TQq71fIQakJ6BatM7Z4TS3QIBcjblXfj/qKXDQ9fBq8biqTNFjtcCy
IzuM0ipFjgLwaKZFtYWzkrgWr4c7U8R1mDgvLOprTwltHr2C83f4w6NZaAFAp6FPbdQJXCRh66lp
sZEpn22KNraWIVCWK46DpO4Y/fvBGp/Tfxap3ECSdfxe4z5dTrdzHtJQsSrUDuQGA19wtTWn2tOl
RE+GmuhRybudOLlHU+tcnF2vtpzApFtKEOwSxR/SgfqMkjpirjfYZbbRzIPZ/afHFkQhs3Z/Kt0Z
LnLXkEte0HuHNW3rveGnFQOM7PNGa72zjRPymnsqCRdnAtyjx41nF37eFyccmn8yujVAkOygth3S
wC994jNfXpvtCgCez9CfEdGRFF0OaraZtYov5g2t4FgTBYb6C4JpEcPvUKaLhE7FrJQbC4uxdSfl
kPsY0u/TpPVMwMxnw46Czpsx+xXJeUxrer7D5Goy8NUACZE4euXBTfFyJlcPg4xjvh3kg7R9s6yI
uwYAHdrrZzhsd+vY5NPkukIXMEKGLVOmxBG/f2QltJ052eYcCtRJtxvMiRaoUh52xWqZIg53CBlA
7esL1uwPBqmP0vxif2IWN43x9qf8nWCCEja1CXDIWY6kLt9c61vL//RvKU+OBxdR8y8MsCswPrLF
MClGHPOr3FANkWsw/GkcmyKKoZgvpo6fTUGjR1BZstUCK/sFI9EwicVq4685z87nq63joWTs9btx
hrq2WOlNT/B6pWXaBumaOMzqKAsRVGnoTCiKtTVWrhG8V9qGvvYqtkg2EpMwz5M5FxpOctTuwafz
JITH8k82HhylnB6Kjpwm0WsALqkSXl3VuissThv0QdlRLly84KkOtvFP0tp8B2DjicLkyf/9IHW7
u+IceSKi5Jg7c1/oTfJhNPHoHH3LmAUAjwWRLdZlv0AfV0JasZ5A3+2lhF4yvMWPJ5kcBDW3/xJn
xktfdkyz1CSxO5w4C15TqFTqBfQSb2azB0aFuF8nsNuW+xgfhntzLzjY3sco1zHCuplg0EJg6h46
PfSeCVD/y5SpOpM+pnmJO3BOXAOulKN9NY/RldCJHZwRprNIsUaXQRZ7BxGjtcePVyOIqV4Hhv5X
BLoc4qreYJEejWrmjgTC/mLFR/GVncVqMyZBoQooL5Ixkm5i3sY15wJtCzEJh6B6ijePc1XGnNN1
+r2nHBCkcLu6MJazsq9/q0mg4TAgq4Fjdy4Na6zciVPxapsGCynULXS04aQ46jNYWT0YkdL1KHNy
VpWLv5fK05Z9cJUpLGOawMU2XZU/Ww7lYmhjqoK3fiUbVh2a41eyHBVFTPGNzx8Jn3xeEfKjvkS1
o7Ea87Yu2Zs3xSYcmQj8cMTB3ctdIgpqUXtylXNNRk6Yyksc/ErHLpuEHyKAO0CHh58Yi4IXIKFW
twSM4fsPM+ifBSzAjmwSarucYK5/l91V8LiMoz7ZQ8xPBstvJ/ZIvEizPEi4qQE7rSzMA4+etAiQ
7zxqPyJk70T2dWK5WGy/q6GHEbJxCymX+7Y31QiI79G/PrC8dRL6UHvpdbLIgW0m7te2o8BZvuiJ
jkVt6QMGZRUZhcgPSWlrhR/U7To4vOo6zVP2E0Ag27u/IiDMfMdi432kkvMMKM+GJTWG7MMzZF0E
ip6duE6RYEuIM9ikVpB33Qn1KE8b7dGeXbPHdHzUJrPGnfMkn2ukjUOxi2okeiQJ0HRbC8mBx59t
qVL+njtsdICCp3Rp34ke40aolIiDBVBsKTYl65nwhCvvVYkTwKEmtYAWi8GQ8h4PUJ7P8QIWak4C
FszsQKGK5qcY5Aw2plFpiAl6t04FeNWb3fqCc83uIFMWWiaFrhF7O8J/zuKzeGViHHhlNalnGS5p
S80FFzrAeHEYbrjBT1jjPNaC87t8KvXze/MF+WY5cOaiAk63fvxGZjtlg1KgVLk9fZz08tsTbwRY
Cf4AJFzmWnxBY9tCrud65HbCEJ74nke5BLri2e5A3j6evtyjfaKXKZyeSOWN/RI7IFEHpK7//uBS
VS0DDa8IYjafFSz+Mvgd1+pby7/lBewH8wFeARMGOvu1QP5EVrWj4yFzE54d0P1r9ROCIRIk8vsa
dfxW63L1hpdvxBoMK2JADDQdte3gmSepfyMNEKrlbjPRntGLNpZX+HsAMOcDJymXm33fBO3AFmws
Y6zgX0mSQN5gvG54Wt1gBIdRRvut0McdzWehjEyfEXYUFxK8o45tlD8xB7tAB6CZL/0EHcIF5f12
bpIKSzUW+j0kNTYXqhHLKc3spADefI3HMJIYJ+Na/suA567W6oHTquB5Q0jkAvLnJBhlgSH5yDYV
m/YG9z1RveUtsYn7auxHRlvVP0U453v38M44T27hXbhOnbYjb9EtRlnw78v52GaBoGpKJ5yA8DHM
l+XKLwvglrwFAewhs1GBRIHiJq31OfeZQoAnAfQn6ZyUHFnYURA13foo0TXpeq5xEDWYXNrgIy9a
H2Fv4jZ4l9AIEBzF/0eM1RZHDPg3HN94bXTUzLTBy59JjpP/RHETYboubW9PaDtyinWHHIYWURjj
bcRDQzNmRbn1CASnYGpJO/4kbBgKJNuP85zfA5smk//DiiIF74QqiAZU3G+qaPQavCzU685ZUBq1
pt61bs8EE4yi1e1X6VawatyMGKcYgip1z/0ss0aaiWN28dKzDsEtKkd6lKkt6nxGC0s9YevtwSUB
Tg7DIqUZ2ZIk/Fxnoos+3/OiSVD4Pzph5K2vFr4rhhx2lX8DlWMJMYpzM8N9F4Kheq6bTi3dOCY+
um8yCY5T4S1RXQ1aYyPCGNLMHs5rHmyBJw02doDpIMIpnLkurbs/PHPyLEn8vIfcSslzxSH8XlI7
4FcQKIrZ280Q6H6/zQcINOaFprS8z9f9l0RRmc0vZbhSHkBMaWqNSX1Qh25Z1+ri304PvKnY/tNC
+mGtFN1IIxUmuWIu0LOnJZrxjmuwovI/G5Gm9ofSlBWWauqOmBidr5uWTKNHtrL7Y/IxCDdVP+/c
QDpqQbqlBcZeD6MTgUawx9uqnAptpNB8Yb2iHUeSN/UL1+O7/5fRB/UoHbF0oaKxKM8t+kyqDBl4
zP9KoVwf9nOk9XnLYQ7VPAsFfZ0jQoz6Y9qS2JDV2V40uaTiNZyC9CrERPwT8GZj7xqgBNrqsV/O
Fe7El8nng0GK1KAOmHOdj4Pif4DnI5oOaSd2o4QICoajV4oUbjUHzRmoz/pzHvdmCjsrMJXqluiG
unSiqs8BCH7r9Fp9VbG3Q/qJpN0MS4O3g+G4+MBCRzleFQKMR0b3jGR3eENP+e8tuz5yQs23x9zK
028emRofTUw3C17mTwW8ACc6VvVM/cztYY+CBGTimuEK/Qb9qoMA7pdCU6+IUAHNFa4HWarNRjY4
48KhGDc2XiOvquEA13EmqU6tX7CAIq5lDjP7F1ygT7k33hTy7BZGBMewVk/nCYbqA9iCmYIS21gc
qqW8xGne91Kv7Rfu6BlwVa3fzj1vuaVnLcCp5dOy8xs56ZU4Tlo/Cad1jUjK5UKrBw/Y5X9XA7Hx
Yc4gMTSvtdUNcj0m46qCNzVcSAhDBlB2M7Rwy3yfXDqRLJIg7DQgl8Z9RQyXWZjzWUf3kAcx5Qys
ePegkcH5ayJBp0b/j5NG9jkwc1Js4+mTe+i/XaybkJIuF26j8+sIT1IkJQfH1hW7o4op0VzAFRZG
8vIsbkmITvnvnMEHhp53xEhPZVduuVIAtDq6jSi+NaHy+1R6QmTsqcO3i1KS5ZWaLRkS9saTlMsx
+p6JhP+y6JEQ81QGfUw2T9aCAmzjQEXi7my5KqgN7ON58P9UOAooNF7ChYAFHgpz/iu8RawFoUty
yQnmzPk2KgvBqnP1zeooe/jDVnLd7KMDv+DtWkh/QqsRZygmnPc0r5JqewCpxcYeBEBPOckcUcY6
+xrrv65/x7pEuziz4QmRgiPdbKsPsZbJEzxijUrxBCUkxRPd3HlPQqkHk4zAcg8yK7/Epbrgkz+v
4V0paEM/eDdOHRxaRev46cLf8dbAtHizaL4GHDlsMDodSpTRYkdvQprgZGi2AE5i+KdeEyAX8ko8
WxHpBzHyUEG4CXsj/zbAIAsEacc7c7s42u6rkSwMKNJHI935NcIh5ulhwsOGS5YUCz/v+0kc4WV6
8TZo7k6Z/dDhOo2ZJC0k9O+C2xYUxnQkwpTglURk+YkmN1hyyunW+I1+dRMSXhwgkXKylZdyyvdc
C/xX21lZwi1v0zLHN36bOreSp6QkuuYuNcV4MEoHgWuB/XRDFhNJikEQgJTvJoNT67bhUEuqIZCT
qP1vs86TpNkst3W7X3k4V0nL+nAAh3p2X82D86M9DnGGHwKmoOwIDC5ztdSyUMnvHEXOOFGjdEzP
zEA4fhso37N/HavcEe6Ha1q5/KA5hrFsfLlPKjMvYB6ZU3ZrYjAm21eoKsv8kl7YZEmAYErBv5ou
cP9ynYqTtrFVWc99q/ltGGLs3G9anZrxMvnQKvTeDTSYE49iJD+shnX33Yvd8/r/yCZAuKg+GLC1
47uZvyzyVJM8NvPnSRRidqk1d5TjthcY88KABWbJvn3MFuTMt74MZhjWHUpm76dbWkMKR65gA3et
qVJxNMdvDjra1LrkJuDWtzRM51+Ns02jUnhUHIlgsqzwBSELk16rt2farvLQcrWsTFvggbakxwu2
gYt0LDHmSGwLN3IsrsvHngAXV+VLYDXkpXwY/a9eFv4AzwSVZGhpuXXb+CswPfCn+325dXyn/har
ik7yT3gvqcUQAZ0faJG5GgV7agH4mNrx2xBRL/AaEY+W7CG+zb4kRG40Ek0Z2dIsTYjijADGpw+b
uREgS69fs2mxGghg3cmca3qtV6BouufaRCphQjRjUFvnZXboRQiUPjYCDMCxm4o8mSKhV6zHC+6z
/icrz3OAQGZngnrfFf4cW8r16Cd4M47+34g7bQwvaSw3b55co3oZvKMI1oWtR9F2kYD7Y6Kf9PLB
cMeHpi5ILoAvoVYeLe5QaAkr43+PZRplAhhcCFGhsqBXlv7Gq9+agXNVzfopGF/CNMGE6NZq7Tpz
an42BbTX7TYFgfrhdKulSfccumnekYGBNMO9iRcqjtkoz5lLDiRyhkZuwLRFJ8HNvoPIMNbSoGg9
+mO+Y8xTwEs8iU5plxPK+JcGHAELm12NEe/SYNSjSnB0Wp2eZuexLmIaeW40uAtB00azaVITKvHY
86wRmsH5n/IU4M6eI1JRQhaHdMM+AB/CH9PaLZSx3dive9KOYLeK+83M6xdDw8BXIeR8xQVN7BMf
Vx3GzOA9aSIpBR/D8kDD40T1skHx4HzY/n103wLmD4GGyLtWpZ+xk22/gmHqdLgBE6cpkobUz2bI
hHmtUNvZvpLkhjYB/oHHM+p4WIxk/wikOlMlUIcZiEejo89uNaTcaFAucF/deE4WGcEV1ERJIVYS
lVrY3hxvo7SMl5/yV7Ibr3Ory3KgIh6hClt1/xZDlr20u2sDwe7+K4h+IJS+Kl4OEnTP98lwMJ1z
L2hcHbSybYR2gKy8SgylDXLxXKg4iSl9aF9mIlflEUGkWAgZRulRtp+KoDXYcZxkwqXJ8GfohbGw
zXFqrx+an4zBNIy37BuvzIly4ftJouTGQCOtRbDucE9KwCl9/JCN33ZR5hkF9geX70vVqX0n8KS/
z8nrxE0080zFQdU0wbIIF7RSl+hl0FhWCOybkMgHxIczK1/cjKeQI6I2mFysAYrPIRWQFMabD8bn
fYKzz58s0YrUbzGkHEliatFuRSBqcF+QdjIy13TDmI+8N/TeyiJnfuWvzocg6L0GQpEfFr3oPZ4D
pyC7pCWtVT7DcaCPA+4Wjx3YuPFSyFBr2pSsBR4/1NbVrYcuL4QCFejYV7MLtMGQO5DbP+J13PE5
B1kGCGimWUh4WEEJGFaamxHIhChaamU1TV6cZ7440UugyzM52g7Xq1VSEmvxOb5CzpWatni8E0us
kUMbqdWpQo9/DcRBTXOtsKzMmwjmLP2xmrbr41PyOJcPlgBSey+AgLLqyll4QMpAUpDIGqxd7laZ
XgX9yuBz3lfFH/qDmIvoyWeOSctzOjz27IH9YRDNYwjLnr+g4s4zuaIBUwUutlO5kN9aqrlo97YY
XR06XevQW9Y72MEuQrPvcaDizpkJlttHLJmlrZjM4YomNXgGdr81f0OGDz+h9WXJGtxDu0eFQxLY
femeV6do1kAdWgRlwWHu+VoITuJAiXmBFjov0l7lpkz0t9JEEXh5fXgq3vLEa8A2MYKSnza5Por9
yVHVitZKDInYV0/QSvgZ1Cu0DVq/glI22qikKTK0Mz7KsG9DR5uSiu8BVn+dPVaP5VnsYe5q66ID
2G2y2cL7dB8yc8yz60p1IsjXw5s2UvYyfPJw58XO9Dd52mY/6fy3XA3UMg+1CYhZSHnaIp/288ak
KSviWG8Ba8cNN/rMone+Z7FZmXkW/nPQ7nZU91a+orhegwVsquh0x6VyPCvM7NJ9nv/8QyAMircj
cREReASuYIJ4bkCO5Qhs/bKbimHrxYOcJ3e9vFH15ZvK8d7OYLyQFXVDg2MNE0lLjVeY+vMnyj6M
fracba4QnxlXf6uBqS2SnalHHss7AknNPbA41HTno97CKG1pssAPORZWAeHttWS+rUpMHXeeEAXl
SiMvPdfxc8G0T9uOvllnVGZJ+bzU/9tsCV3C4jLyZQy290PO+905CuYphfCLD256ng7v+l/RRSDV
mtkPIAxdfcwhvQAPaJJrPq/cuYhYJjGxlngzUAygLQOWbencCUgWeNGnavMk8/JKWvbC4UovIDgs
79pm7xCm0Unf/ORjvYFV8k0fEijMBAlxSsfZhYEWhhc5Pns5WkKD+r9si8yTeNo9Q4LIF+0Kfu4i
NlpryoGbJE5OpZerQ0nZfrmIOEOrhTEqWudbhT7xLVk/6WB2GqoOPBSETbVeFmTFz/A+J4BQtAyA
+2XvPjg6+8dM/S4mVfaijbSk8pc0cXZosNf/i41lLhy+L/ECr/ZMECKuPO/HSDhxwW4IKry0tZJQ
assRyugxHBsZ2v8E8AyRmlpbYdfLioOTrRi+P96E6xx/UbEethi8n00WrKaWwQrWW6jgG+adjuOk
8xVVuTFHWvZ8+PdWYRt1Cyl0+XxL3MUuvlTQNqw0itSf7xvfZSs6XDwdsHMGaqPXaFqVVkKHWggY
aokGQ59xBZSaH3Mg14TujabwqavziMToylvSW2kQyx3FKtL2HzxRrxCnD7tD5KxLakQgeDMv4CnS
Vbr/6bW88NVtrQ7a1gIqzhmVuGBabzqH06LMYHoGKjtMXRtSwYzzDg/wVVA56MZtnlpFl+P26UcI
UMrXPl1Ici6g4YwNb0BfdNiCOUNA0DQLCkdEg1Zojml35qBeyaorKG2a10X9ZfHUT+waftd+gpvR
43DVeX+CoKlx0Yt6LWVswPLbUB9Qw0R6Ylpb+eD7z2feWSIvaeEMkfoXI6OVXN46dzPMdMfY/GgH
UkvImNtcAmHwVpFFho6ZeEIDdg0FYSTmZ28nJtyl5lJKkW6LKdbP8e4R+vPBZsAkwYYuR4HCt1s4
7CFcajTGNZRuZvs6dO5nTGlybCW0ij0sgH8UfrBVZHfEc9ofpnAyw3v6kIwtsc/GVlbDt3S/qlD4
T+YV4A4bk2cE1BAUSECU7GNoaUcM9upzSWEzBMqYITwhlKkxtfZ2IZfTKLI9P7PhuzRf8K/uBGyr
jooFv2KJP99pInNoLPqc3fK7bypt+UdGOV5R+1GdT5ZJXoeA9SzJKnj3odq1jeXO//cQFL/FvLuW
lnANT7A+2zDGJKVdEAUKD3VAJ4L4wqPONu3ojArRLOB0yAJZpSlIKFtC8bibIAO50i+7wczc6FCL
qvpqNQopI8f3vQGYGZEyZdw3i/eHkxV7L2JVjnmJo8YqA9W/eU/TlxbwXO38p3Y3Oic3Z1G1K1+G
d7fcjSVOObZOFo7BQTlLmSFlD5pRotV0dI5H90Q6xLPtyLKKsJMFBvo8VOTnWv//4+JOhMfjZhBu
FqaM5zdWwfGc0fuFOdDOZrA+2IveYX1odK025hrEHsWGfI0yZzAIfsckMoygaU7aPAE6eVDVEXTJ
alFPuMzXqAdiYc7TZFxrm8WxaK0+8Z+MrX98i+bGb8QZpbwdeCo/DNv1NOff8+b4bhCYXOPmMVJw
4HQbPRUCy5ymYX0ecZAOHyatFzrCQQ4A/iXcOV9pF/vqkg9W3mOxNdS7FtcJ8+1C4jBqc91d3N0C
8Z+iaUJcINFjVxBKXdoT/SfGeUQV8vAl+3miP9K0T+NEtsf/JIKiHrnVihvKwaJX10z+wTYxT48K
crjd4hPx1PgRCvyGFpwFRpuQoTH5SjUeHGZdPiPTEPDlRSDls7wUc/tSyuvpIC9wr6xCG5mLiT2T
UtfoRfKo6ACt3xFEQGF45VPqtR9hbR7kNftdqrSePIUt2iO36v6tioaz9naqeRPMopaqabERXRO2
/9dX3u8Eyq3HujGeuzZOt0werSNrZzwE1mLfehOSrGiWgPTFFGxsdIoi/iV2/zo6whdPuvnDzahD
m+13SWUG0EeSoU89C9chYHlrHKlGw55mipBHxKYRz+hVGIGEmTum6s/ocI9CCVPvfJUoVea8BPoH
84DX238rfdejSlKQutVjic59A5UUq6tClVahMId7Rn3WLsx/HjnsZ989VNGu79L8I9UkWjpuPgjt
EJBfIEwGkIsqkuyGGvRrAZb4ljWBzXEfaVtplEPDO0GB86y2TZ5EeeKb63qgEIcQtVL4tDA1w6V/
IaHKaPeyxrXMwtq1rh8aLRnDPrtc9QHGgJkerTu5KdudGXZSZS2MOuMiKOIEknqml/B13THHNnCl
9JEQK/hLXUdxuxkzZDUVSd4QwoOzsP4VgKKVWxiNMCTqpuDdmlVU0V/1ij+hoSErXjjTEq+L3y8n
BoSlWla/+4nWrm8VpdtzO6uIp/oiXglHrZAP+j5+GrngY7i2qIafRGAM5+DfNsd5z8KJ6Y9I9ACZ
bDtHxagrF7a6sZL4zVOtzkdBMzSDCNsAQ5cPSkHADliP/GKRQa+pTQtpkqlp0FT+p6tjJj+mL2yy
aRDKIkFEty4b7fS/QS0mkTPB+eiXkulPlohmfbnoCHJ+IFMJCNeKg57kPINidMZ1joDYfvk8b41c
YAW8AV6LjAp88faWrfzyeQLMeOxA1og2618bDOdkL7IZNCj4xV7nCGPzIPCEO2NPB5Cdfvbspnh7
5uh/mBCDBzWdYirkvf9vj4kJlr3hdV63dAdIJ1femJ4j6EG1ZEQs9/8/mbYe/5S0JbXkCzAwl8C8
Y3UzJS/sQStBpSPlVyhhCx5BZjLAZTeD2T7ek1J9uvZ4q78y2Yhun3NHo0OXile76b95Qb3yx+vL
+gZCqwnQsC7NA1l8JOvfdHGZEwgS0B8TLogusnLMYPL3GQFt2CHsI1mY3R7DG/1Rp4xhpDcLPdiD
zJC9Hmdt/23qpMYawjvZ3T/A9kFvKuS5T/DPUqNuIXZ5I7uuh09eMQ1mrShzKRuJTpVRhHVaAIba
l+UFiIQ/pkVXYe+1qevW1Z0TU774JPzN/eVnBZcHxnhs3aXoZdXkALn86lqH+s9n+uvCTZxE60v8
K17a6rVHeGpLGvU8PL94vvP0fSRbuHh5qMTaHQWOkCmum6RwWDkul4wXP91UQsSHpcucANlNG4Tc
BGdkhhMxQ3dnrV7XCgJCW0EoWB0TFxMaoAGYrzQ3eVaA9Izd0HpL7ETLuhTfWp+yJWGa2OKJ5XJk
ZUmePeoeJxKMXNqV2AUHapofRtVRRC5BTcYDDvdUfqnmU2HM4C8YuZXGeO/S/OGGYlRxUTo63lK/
bidMG83tWyltur7D4HGerBur6A6Wrjtq722a00GvoU/dFiHfvn8MUucZ2/Ssx359hzuY+BRt7Rnl
7GGxP9altZVZzKtzyGnFBUq2hm9oIFmozLZwjrIvtPqO+9y0n/UM1WOudHgRAfYlihU3UX48CR+l
8X07HiM951j82TAAWvvd3eN0289wbZYUo0DjCopBMIqgJJBxypvh1TD2Q+5RWpgPtAYiyOklJQig
tLJlB5uupY1hRMDP2rQHUH9ElKJg4OLyg7RyQDW5NjsaHgvj9uhiBL0EMzQNEqKsfK3MCyu8wZwA
5c8s+AHewnATz7c0cmVL8hXjvQlSfbXnQk669/I1MlfHj9A3Bt04plTEDj+uvrPsjueNlWDhEE6c
JR1XqtKpMcxSjDy4IfYRIpVwkWJoPfo72I/9utnD2OEDVqVI5P3Yo/rJRHwHpyK5eEWfd/ocuj9w
oWQvd2B0PXAWfGUbOmx7ybHSPAcSv3Cc8oKoDph8jMGTFyqagy5PNPEqxj3gRAnndAwIDHaAsy2u
LwWwuQd6Dhtmfmi92uXvS0IHjt6lBIOayDvZjkLpTlGQiXLQ6rLxU5tStBMNYPzNcN+BeY6Aillt
YilBPWWQNOoeAvUM6GTMe3Aui60kqE0codGcZQa4v06NCQJrZFydj1koMvWNx06YFoM1RpeC6JPc
AVvPe8+mlUXtUi3RdQf8SObHqvnhCJscxSlz6IQiFh78lnEiDFC6cj70sX52atemlb0EfKU1mYLk
EThr48lIFG4tqoj0Nzj8idH6pdYMhUV3qZ+1C4vsifmWyj5K1yItiW/iLrjK9UKdMOQN/kXfT1I5
lRSuSErIXVXl+eao1UsaXBiPK1qFQKX8pcminCghDhpDwuGKCbz0I5YW/J8teH/6V9rADaACZbHm
YFxE7pC3Lqzq2MNLdSfmlT74UKVTdNjs1XjvA/Z5ky4plW/DT7cGMs3WNiUGMfk1Pon+sHEquOrF
VRq4up66DwXlTY0t6xu6r1xh5HMzZ7SoWsv8GRZ1xABGkrSXrMkp31IzDkMFRForDed7jJrGAaMW
2wPpQjepWw63dQCj8VwkFvCUk4Ix24lC2Muk7kLRd5zJKb60HUgy4Fk49jApvXhSGuOGY601pvvB
b9MDNBE7OE/WyZZk7Ses1tonSdi+javIxu1o/JFjdohJ+V2iJTc9aVKNT6j9JQGrMRmx9FVMaraH
3iXwzgiPcg9LIhOQ2fT/tq1Rm8HPkYvRh2+cR20iFE381gtST9F5X8XTY/kPjcNo8cI5xu35V7hb
+fIkuLHXF1JKO1ESeSFTIipCJ4LJgcwhlJ5zi/QraXrv4NyKRotvjWdJM4PdCBEOH8oiuuOQ8+SO
V1c8/uLO8SFqRltOV07iT9I5phyeC6h3TvYaiDKPQBJn4ag+zvo14BBdVaMUXNG7W4glCDniuAyy
KBSvDfXh8Vodh7qW+16KOcmUTI3Ty+PJmPbzo1lAT0VM/MydJs8yD8OW5EN6LZfvIHamK2rWDLhH
tHw4M5UNKx9LdkwvGq8DcXDaFWrArcFznyufXE1p8ulpKoUwXlvDvSlejzaqTLRViQtF9yrKmdo7
XgLQ7bC+kH9MQ70LgGFMFvVMOQCM6OE2u1k4VeLQAEppdxt3QB8P61cArYEpCa7CUDalY5mdubQo
yuPHVKSjoNQAsRFlnCIvCIVGKugzyEth23q+JYwCSwRMdVGPyAas8eO44yJEvSmGZcy5aJJhnyQG
Dj4zoFHJhzZebLJBygSBtEWJN84StfaVYz9h6i3+6cL9eCOgL3dGXa90pBWJnku+UOQuUnUA0Q8k
8SK+RQxIGzPX3iDFR8p9maeNlxxoOlAgMLjUz1Znf4fSKPfNSLS2XA60PYgw2acZjnsezVDtXW3j
obwYZw/iKx96fpHzBe4AGcWvnNWvaF/b7RjbIkMWSniii+9sp078fti90DlE4GjSBN/UEqdufRgN
u4u8H2X7dFdW6gylN0lgKCozcsxeh1Cs4zxocxSgEZex7ai1DLbA29yTDTrTUsJatrTh0K5D6qyC
/orKoV3N6R8AbIkAexlvsuv5qAhNdM14PGXNaBzmAjTS8S6w/tV4OrzrJPdA+onGJiigo3kJrjzO
WON03B20ElI2kzioUbiv9iiVSUp+v6kv65b6g7Fz7k0u6MX9SHPucQp0zGwY+FOKGUXNl2YVYJrT
htqisPkKsSaseEexELIndAkiFjCJl5nJNVNjz4JaAfqv568a58D/oGC9XQOTsMzzcAR25k8sDkTZ
VaBP54hFwd/up0XEWqMnEyM6kG2gd6n8nbjFBeQEEzDSf8fIm/wCiw9STRAgQemN20FRv3I6SQxb
i6x6zQh7783WwAsFjaaIc+ESNQnCsgloNdAjhPJWkc/qi5dNGp4bgq02XaiwuQhUHRQtFgy3VhQn
TZBdv4HFeR9iC7ZAnAysOhVZgnBjKvJjzfXb+onNhVGEo0bUhYLcMdw6ZOsx6z6AckrtcYdneG8k
imp6Of9EzuNZZCtsFJtArmh6QVbmwJWKshCmwLXlKV05pPb+0tMQWC5xSW0C7SpMp4RnLzCuQijb
QJkMikCuIIOTCd4cmmJ4qUrbbOfOH0Bdz3Gzd+LO6+cGFRkcuykFAo4W5KeiEdOhzbt6m0pcSAk1
UY1oXRsN/Yf/3Cxz4ZpbECOTmmCYb4B4eb1yRGAq7yhtpZTqcx3xE/74TOhnrh/igQDf8ZcSrvrT
LItYZkwXeTzTej8YKhkJ4tXRQEM91XPOBEcw0Ogj6PbQjX7L1CUFefCwnPBqOrxALVK7D8MIPTV3
7S2kZgSKi317OyLvuAbQpugyUkbw+82cNo0AYxJoBseP356K4YIvTl7Xf9uoKM0fP1Xxknd3nGXW
ZgMyNvIxVU8ExHNL3wj5BOZ7+/0xeOBYqNKWFETusbXpCWTHbmv4nVY0lFNpIbeaZiIIr2FDAkWb
xHE7W4KyDiwd676YQ2HJp5bCQH0obuhT+wlGbKyiBnTHkjUTwk/24x2GodZ65L4qSF4v8yIs+lWB
zW3L/CC+KJnMr+aJ0wA6bQFi6O7mrgMerYhMbTOP3DHSX7j7Wna09Gt9xpZBUxO9fRoS0P+tgdcM
mMjLl+6OYvQXRwTf8yrV0kmJSwJS10+M60N48+RIqK6basg2TEPyMYZKoQMZFdgx+S+xmf0gUFjp
VCDiosoxEKmHrDC0VoOIgC59MKyF+/hE0vo0Cux7kAdu7wh///v9KerJ2Hc2rYRtUiR5QDhM+BwR
zCK0vQhW2bE6I4B8DoFyLEfVQzRiuzMNZeAzYpHqXR31mf9AJr+Yro/oixTbShiIw0ts2BNkRbYS
fEWlayBcVPYdApZbype92XigcCGAOPlNuXFX816jj/6gWdbQdSgl/l+pSiTold5S/D3E+iZddI4v
iVrOcl7y8va39QWwTnzc11/IaPPOuquLHoB6eOf9hV4N/OSLHUmgMBKZahmekorrlNfDn4kkeEGC
rlu3QPvNMZAS/yJS0j3K5pu10XExO+gVH0AwczSJxCUdlDgQnDn8UCkRq63uQNO9UlL89hhVaNYF
nPNbF3zu3GrdSfJGWQX0qZYI/R3dap6obWlpUN5QaK9Ow1wPXiXgL124u/4krTIPOna8FSnU6/P/
RWMFBObzsfdXxuxarmHVztgVr86mVsAcUyIZ/I/2yUyTVtFUQ9dn5+DJYQWCJVyIvKjPfydAJF8m
/pRUfBxxvZ25YYhEIUdOIVLmAQLD5IVmw+Cn1NrHbe6NO1Jopbgjt04rcEpsRuqT3+c8YRlByCOL
2+O3BRy0ZRB6/HuopvK/5TwP3ROu+YcUHIi4RzgqscrsBfjBt+CCo3ZQaOlkDzCAjOsaXU6DhgGt
NLWc2NYTNhOiVzDOB6ts+wsfHmbmWTI9ENJsVy3uohL1L9TLabLwULp9+U7WlNzrq2KnJx6DXscw
uiPOcbmMbya2XyJ4BlIYuUY/8y5No1f2pOsNsNODQjBEXVnj+HmXjUQMXxF9XFxry2tDj3lrzOKU
VLQpJ/b7+fWIpfl6lSq6XnIfB/PA5ChudNNSeqsJfzOT3uNkXSwcUa/mVHUY5jVONA5dk1rYeBTj
ZRD6s2rLvuSlTngCFheibw9TzT7/hO8WJbCVNFZXGWA6n75McOWjs8DQDHOjalaeKnp3zKSX+DoJ
odSSGZDE3FOyKltjAjQg1djfB/bdvupOfugkqZ3QsCcW5esvkoLsqyt3EIX5Ny79CTpl18rjwmZE
DQ4fvkWRfIeiuCc0cig/0SH24bpuJhween2Q/yk4oGr4h/JtGbu2z0qAm60s7zu8p3QGcm+ktFI4
mt1NDCqeLnHklXCUgQzlWVqHpB/NWwlpvh9bsCLkezAS30sOEb60xvu1paqGE7ZPCNhTp2iBdnoP
eFbWoQvXKaAmA/ZG9+BlIudRdxcI+mUOsWplZCfgt/Tp129KUkNqbuWCTCp3e/Q31npbqJppgSOn
Tf3CCiu99HHAuZDQt14TrEDCPowTo4ATrVtQ7dSAilYACJIVO3Rbnq4q52NFDCdD0BL0eRHh207W
jMzwEll46hoSt0dJP7kvyEguJyqvxdfdnAwBIb0THmUnvPey6Smr/RYAVz1yvBgGjeKiDBcubxux
TmWhUk29R+ypmFA8DXJH4ThFX9TgipReZe6C19Doxj325al6vQpKpWgyc1LcsriQ1SrzTUvfgwPD
aH5/3I/W5+Q4tKC/q3RvN/CLqNaetZ/UHl0IkZeSN1CtMKbEMhIs5tY+Vcj/hTAFIiF1Th2PbBYQ
imCrlkbMIrM7pbpEW+m0R/te4s2iZg4B0vcOxKxFDq6wzLjULz+ScRCUVnRV85rJiK9t8wQOnBD9
12KTWhdvL+yaW48Y+6mif0dBhmtOPNbAzMpZanXQOloDwOU8qhurHRIr+3leBYaxBhR5zwCn2oyB
93vm1vO7KnlxR821N1NueQx/DLq6kRIq1JzMmeQN1W4WG6w0hdjyS71MvaLQO8Fmb0wRz5qfNZs6
jsFkp3tcsjH5mQ9GcDDwGAVNylSt8jKJGan4JBeQNZWWP63ur+M4+M9G4TlMUoVRAH0IbWi/iRy+
ZffhmTTBnfDJ4VQ1ejZaJzHzEBcU/H6dyGSOs2P48hnSUw8+OkPtu11CqjnMUiCzOJK0JrU+GiB7
0cZQ8NTgbDCcJ5QBPVy+kh66PURnewxraWMxX0oaphkN1MXC6um5P+opSbE7pGmlkMUFdu2rTQUp
Q4yZ+qWNtIY3B/mgx0ZrcwvuTH1UyvJe292TMRVzjFM6WXEbvsU0jmF8CrH9PRaHNgzmzvVvmE2E
Qeb3sLzkW2M4hNzy6hAGZXlIGZAlww/9lQG5VCdN9EPjE0+atwfFGd/evHlg+wsUQcP0LM3EUQOW
79b5q7e0NXbd5HEgrAFTKKvZt1wHmKHsVc20JnCYtJaukf+BofOAyJWdPGk6/QIDMFyrohdwHDrn
agbfzX8K+zkbHU1+2jFDUDtZTuQf7Jrvbtqoe4K/vafz976LtJ1+1CNEmIfti3ki+2y0q7FRsQFq
PbiH+0V7h8M11Ni+phXLZzM/uYDkdR2ZiIhSetRHzkKwD2fbdpYc4zEJ4ZSCAcnynK1Z1qBTcnFV
Fy3vYe+LIxhYLlwZthKiq9zPOPTJFmnDFEJEgecG+Bbii0fF7NNs/m4WmFXoXah/EC6f1IvQCd9W
mGLBYKLruoTWquB8ERca3RLZGiDuMFP90llAw/t++i/XVkrLY3hHDX/cYnIXTcbwXSo2wjb11U3E
n5eJGSFuW2/BynZoDOKR0Z+dbcuB2hpc7QlFEIkooNj922iJI+rBjx1ui0Yf/5dHTZDzQcfQLFRh
IitndbGBfYgJFWmB8LCRve0hnuYeYAaoGETkYIHNNaZLizAG+7cXYNoyZ5VRjz/rueC4VHzVh1Vo
Ec398FTf+VzAROhptPuOC22QXl6YonG94o113hiJuAixPpB+t3GY6pwESacKl3idnsSDJQIpo0ZV
tBS9UPBw7qIaAwXl3QdH4bU5791oh5rOBRj3sw86ojqlPF4UAievmpZLKBb5qiMv9Njil9ZdAoO9
HnXNea4gdJB1TEEsG+ixJqF0C9Egxk2b0eDEsZXdRvOYW3no+vNwhGUYkRuHNkZ/viex8twQU9bm
7Oj9aCUASzIfhxB0yH15CKFXFEyuu/f34fNPgq1QYpW5Rv47/G6zNEWe8V4chobVnK7na9D9X0s2
y2NwF0h7b0Q0Sd2FgtVZGz6KdmhcOkWFrUxRYhDq2NiufM/fa4iB2RBst9rUMT/Gyd+eUSC34YwR
bmuXP/47peQhRk+oF8RjsnbiB14EBbZRoV/7MZtZ9uBsv9Dh+66JhxLkPAoxF8/5IFMmjKsgo8nR
sSNTUpxjdYIgQh/PK+72Z+b8MK4vfz4MYWwy5J7n5SBhtd2OUNao92+EqU8AobaS3oHB1ZuhvJB7
4WknyyeiG4paqNThyAqo6EZsXDlH7dgH/6c8z0F8YtkQchH1Ui3Rq6fcUmuRH7SBxd4uueO9oqJy
U5DMAxYjR8OyUfj+JJzXSvA4PXtmmsVpldo6Yit/t2ugLHFAqRKEEO6Xm4p+/WaXASOR0jW5JbX2
Q5xwg23Q89LPG1J8R6QjrBGcnR15DBmI5wwqcwyRltUfrBsyNssrIdQuBINSFbWu4Wy6AQlxx4Z0
w3U39+CJkJvASGuptAZDc+cMEFqfQpmnZGY9zsi12cyTuJm3Qf8+buK/u9rMW3eF1IyZIoZkRDu0
tGaxkcEVzT74Kzf8QOzScEBqBCSGQayZyzaXiH1RLmIdPy9j43Ksx+mABs2Q2k0WHeS8Jp/Z5wF7
INmCOwkbiKnpXf57yZ/494X40F1tDPDGElPjWlJ9H1tx+JNNOuApCai358quH+uE88AdtNvvmY/Y
YyrYGasQD8/eYAVWjbTXpKriYkilEhHpRCErrLGxvKmDYVVp5zWjCRFqtQiICcFqmL5CVsjtiOa6
T14IdJuQ/AKCr7WEoi+pcnuaRcOn4eOnCzPxpvIMcpNxJ98Yt76Zv0A/ZeGlaZG49AX4LgadJP+T
dM0QjDKAyMVGlCQsLGXm4gQnlvXGOoODO/R0lXBzZytDO97OQSI5InkKDL0DUZsPDy265TxM788B
d9wOkEpS5lAjTT1L4eaLzKz4wqoRzAWLMknUCT/DJO6RoZTxox71jJsxZkctpA5Gbu2HyzcQougq
jKHfqCFgchcA9q8uGQTCci71ahsju/rMsgbLXhPDe4hCeAHZ4wm88iYN1Vs+jMT+c4GidLYgaiE6
9cbykA1Q1KkqrHSivsxaLQFWk3hhKCXVc1mYaAH2D8ZhmFjsr+FvEk+3YbLGPYEczXZCw/mK0zeh
prlO2nRCxw2mfK+bEo1t32DGAp15n0J87FKOCYqdEVUfHepETo923zzmoRIcnHPINXWCJ7HKpGEl
/tn3gmCZIBd7SNdjWu672SFDfo1Nv2GB0BXzqhUXc+Ayaf0JOkbQHWusfHNq+n3nVFY/rU2THNc/
rXRhQRxTVKrTsKIhegfGZuchFL6qdJSgycZ+xaAvWcTWXpGnJygpiqO0q70htaeJgOxB06zmNvwn
ZIy/u/tIL/BllGCfv2z+cL7eBnEaczGY3kE/8QzaianHfbe8wa97SufDq6M4wZchmebiQpN5WpKA
/4akwl7RFcWF9rEgdL40XF5/kRfshiYHUBM4RphcirYiTbp5/u71LtaAP5T5NKB7JI0vQMjOUpBE
8MmqPjaiDGm6eGd7+fgZhWhyISjQnGH8v5jPbEdb1k9uQs+pcNgwqmXUCsWGzkKamWGHwl2DrKxb
2aF+kSrK0hVr7KTaPW1ESX6DDDF9RNvKz84GfATgUkPcPoQrOlEoAWjFMjtlJkVSWRgxkn0st7V9
tyH9AJBVuoyf1bZYQ6/yD0NJzOkEzsnsHSex2Vzo/8xB/OmEXT0vAlzDuZhcpRQP6Ieb59VKY5Ro
OiN0RVjd8E8f/qblexQo6LERu5G6eNFea8dStU7EUcG+ZkBc4vuqSGLpUX4LhssVKfd0sj1azlNJ
ON2R14JTxFhBHC+zmCTNYXn78+j1/NbSMC7Mb0SjGLb8mZpJuFXBxkIcp1QWFwjTdr8rpyH+Kol8
iPWrUXWIex8m13XvNdgq1blLxOjLhUa9BqQh/JKG8cZa8XL7JeQpACBeNelSyoR0jcfov/wMLMBu
5Ft+D1WotcHkSM+uZ/1AkmyLsTBIW3zs8C7359EnNH0PINHtGI8mBQHJbdOuz7l3d/C0RqiFuO8K
6F73sU2u+9wizBD2NI2TjxSCUbvd/cZ6V0Xvjluei8wYM/b1FM8HZ++Db0iDAkwhgwc7IJP8/PJF
WX1cYDVXhbnd1219dqyuAB4cWdVbp/x2yHk9x0HwdEyDKOzeuHn5MPkA3Hohs4nis9c8ajM8fTSc
7C7lHYjPA+KZKL+2mMooyAIyUtkguW6yvrv+kxUdwu3e2v/0junba7WE1s74HVm4gs2y6rY1Oel3
Rac5hYJI5A8Us5vIqbiI0pnQZ4Btrk0DMraPsCavTkVsU5knaWG0hii3HM9OpC3x62pyvjChofKj
5zZ8hvtce7kNqNJuak1MlgLBF3XZB/0TPJKipfyEEvnSXRX2W6Qv8Z+fa1o71lzoWzNJBBgQo1Z8
jG+kalPtj/ZEXpXqk5+uoYEOPUev75KKFRYlZzyNtWAKSY6Yz6veN5NSkGrnC3DwMFDhzTkZAV3o
i6U37719duHGEzSRoczeEH7qXDmqUiVbfvRmeuOClqK6RUOlRY6G3MyiEnZpg7qkokty56VONDTk
aNUymaGfjdc6JrF0u8XMTQncgGIJ+TjX3E/8RoQdxCk8q7voSLFkIE1O7pp1BHDaBOkK91ZuCubW
6Yi/kKp5Qtcitq9CDKQu4efaw+LeHVJXAAikt4YmrG/fvjvBE9HpaxN/5saKwhrvf61YEeQHgAh1
SaLkobdjRSHeOyPm8kSmrRXJcYuHV0i3BC2OTM7onia3wiRpj59UzjVOPkYXDQOE+nWbOENfacm1
2jG0Ab+6W27RxH7+oajP5BSJZ9tEyMZo0e68Z79KEHY5uQkdQYV/M9hvLAIunPh7mQEsNEhXE6U/
g1kGZ3r2uqBKirBVnRhbnGKjsmwX3PdBJ15/muqEkmSuOqs5+vlaHvbtaOuA36di8veyKMXETDZ3
qvjv86YhJlPmss+1OWOiVecUto4Dp4BOZi94k3m9CVU4NCRnccvfQz2Kr4MAwaLeScfp++6f/Fbj
Y+QXQ0PGgjqL7lh4ib5w59AtflMmPUCxtcAn7UB0XKl7XS3BCtg1tAdtPiJ2cCgVbul6Bi6+YltT
fLF3/NXmeUkPO96EHg4TP7iebkt3fr/ghWrITjL68e0uPyQyO642T/ahOiysrAgh5xjEWU4yhNqL
+TXpmkqRwsqqb5uhBinO7HhmEiTNUs0fDaXXluCbhaJmjOGs3PiKxchakqbyc8jK+wr4DCHzyi+E
U2/uzI0D2WZAvb1Csnwsug6/gBLtjNM/5yPmLcLJOykN7o3oOU5Q/kIgHfgdkaq6rzNOweZSrV6c
1wvM/WX0Fbx1JJR18dM4AsdJy8bsSbudCmhZkiUbgyVc1MUGDvkISbfaET+IrxS94Qq2x9I+bEqZ
ncI/rPzC5Swc/Jq3uGk0HpUyRMJ6/d+yHOT7M5j1sWTag69NtfWmXb/TweX171g6tnmEIXbwVAnE
P9Efu1Gry7Uqs4xaNsP4WU0fy8xEbsM8VX2GT6wBuzS5S29PTHxl+Xy9K0+0tRoQVb0U0+fZeIm6
Tdore4E12xIlht9X0BOkQEXJNC4ZOISCj0I7Yg/Fd09lGlwWsBjCg1VZQ6zkFQCW7Wxyz60e1OZe
x8OwfbFrH24k4oZk2UjO4/Vcpw03SHqgC/AduVOrXwx3yOwEHTx3F6yfEsosvk1n/PXOHfvbWfWk
A5wz3ZoV89SfoHqTjI63lTvoFTUOpLYCRPM7VXwiqElN5rJRaYvDkfCREzm67pdXuaD1eJEyvJEJ
PKYPBzAwKEZaBSl1pchmfhSMZ4mya8HtJ0E3bonUhtdsZ3vxwM4b6U8OWiow0LIb7DLB5n/Ki/u8
UBXcRZgRV6CwZ7csPdUnc+mRJaTLvGwjKdOWbtpJv+7dnvJRdVnWJEQU7ZRoaRP428C2r30dPTGT
aOLkGzBVRsklBsmmqMmTbMXD8+5cfC8uwntoBoBiZpgCpyPFAiWRSd4F/euqavLw4Bx/jDG9NBbx
UZye0F5/ZgNNF7uP8mCsQJ/jYqoSq3sHswXNDeBoJgTv4DgONYUCqdhxmnxfj6ybq6jsXg7b9dIT
XhIHTTyp2j1UgCH/np+K4wqTWsLXL47/FB3tPdLBlK5IVTrFB1qPCnL9o5iROHZMDvaTWRARZiuB
Hv9hiZNcxNcTltx7aEcE1itmH7sWG2DK1lmc9oCXp25Z2Jdc2ckW0Znz9tQO0Z7aaKmdDCxJAaER
126v/IjDHHmYcHKPTYZ79OdRUJmQmfJ77Qxz8t6mCFnnQnoY8D4M319K4SY+jOhMdcDXdMufytSe
LQV1PloogOKjAdDFzdtdVDok1y09C92oPXHt8SkX/14t8fZbnIhoaYkKT46LudRX0NFG2x2YdR9S
oQI/brF20iIXUgXb7untOjQV37kngcajgiGsviZxEVZ3jcb4e8igM1TfS22G3sRQAox6leJgJjct
/pzoOlNIH1YyqFEOjiAczUz1bBFoGSYY0o3HcE7l/upn3tc+tumykFLpEfNdcKS9c9jb21lEyC1e
TlyqofMly8rvHFdfwIYaYxYD4Ai01u/u8AP7tmlfE04WtLx9Lycom5toPjg73rboQL0L0jrpdDCs
CU1rFx/xUZzh2ZHDpVUoUjr3ikoXqiQ7itu8o1midvroR0iT7yeAQ+ywpzhFUKQU2kBlCXjAw3eQ
+C7Bazr719C1oxSumfnzgnBAoxKgMNooILeKovu8aznQGxABmfW6q+obwu6Fu+S4A+B6FyPBp/Va
T1/4TiP4m5jSUvn08w9y0ehDbcrfSBBvYUpSzc0ftvupT0w5sQFVdH1YlmTHpaEdN6z2HsxHP3AH
sUVCJQaclszvKSjB6dXVoCJfCVRXsgkGfAAod3q3Zfqq1UabkOd5+ohmLy3ISjdKpax6HSfLXJ+D
YulyJD9SWCLOvzHGhm7s0Pk4HBDv2x3bwGujkbDVfJbn55coYYp7UdAQHZfYRuZAAUK14Kq/Xo38
B1tYu94rR1CzpxaCKMWzZPf7xsu7cm6FPjbZQefwDZtv9URj0lZCchLCsD3AxAiGz/Ck8I8c3ksm
JAfbbyqOgDI9c0VQ2F3CF7aWotikLk0J7JKpkgvBSVuEsEHjEgh4f1O4qlCl3Fk1q6z8CNTjpDLZ
JoIo2Ax/iXo/U2pATDrjDSMvqIZXpna20vXw7EqfQsFRFl8t0cDUhnmQBJmq4nLMdr13G0f12AX0
NOgaf/zSjaTxP1o1AR+TjKp2ah+hcz4ZTc1/X8DQbDz4lqQ+poX802ubqqEMHfmndBjYr7WT+SJ7
qDVSi1NUPSff77MZCHzCQmU30m7YHjpCr60H6+mSlwYwUZkWcYKIoD5i1SiPeXn3rEzsl93v+pWE
Z3DDJ5PnMtUwputKEMz35hh21wxvA2viL69i4oKGZiMqQCYeyopdL2xGTRvFeXxUGB+Cj3i7o29h
z8kE71XeVpM811kDXBconGh7IaN+2eAgkPdwOx9c2mX/eK4YM2B7zCMZjGxoC97mMk+tLe7em53Y
Dd54SvIBqGIkBAPzx4RE03k2Zh1mh7/yINoampOzXFSF/EAUVp1djhffAq/bANyMjUuxn4xH/2/P
3gu4Rf+RtlZiWVOXMgnRHsFQow8oG3oEtJzkK1vwibzup2/M9NaiBHZ2KXls2BlYv+Emp0kFeDKO
pw8POBtagTZoWwRfPagi5xO5/TtdNWzgYmvH0Zleuo+hcjTuj2voJ7SfhvXxkVPo4uch9GtHK2/g
NZjzJeDIpg2n4C7Oejll3UxJfqw4iui6OqdwjsmBDlyAr+lwitxEAVQkKgvaWYxFd6H+PGkdfTLc
veC6X1d11FTnAvJOnKKG4yZVYzRR9zxImRB4RcuJMc5gF0JsunaOLzSwNGkdkE+8jcrEWIRucXBz
pvnmQXOycyHWRdBxfIs6W47epS066T1I+Xy/FZBYc632QaFlTkPxdJG+gh73KCb0gLCKkneJjSnA
9WELIdTyMDNWQ6uP9zrVowddgtjcKc2zu1ubXl3tpbi6HTgFsvR33TNWN3ibY7wRFJa1psW0nWTC
IR8DQvUylMJUpO2rmwwAAlHf1kLr7O+B0tbiXXKtEP1ZQFn+Ts1JMNXCCTJU5UZJ06eYkjpzPOTk
SsHlt2OnF5VbgGgQnmHjczFSzynfnqR+7VUOYrUTUIU/k+ySE98NSnIOtaim1sLehNsGz9GMefUU
WsPaHVVnVBaUYuRPLxqM0ELf7DIWONlJICtIPJlBQZ+YZg9DTHc1k2wXAFltQEd65Hph7cPE4Ani
Ton+SCN32QE7mJeqPVTgiwCCwnmBcSNdeGhAHronEb0RARUJ10wYhyjgbUnVG/YV8wLYzwoFD/16
sc/0pz1KSp0EMk3hft6hoLMajwRYW22Lkk7CGDY7witYI8Tx7e5673TAkbDCtOf/sR3PwQFPWncl
S3pL+TnYXSJykPKsdcf6Gu8CfMPnm7MTL+PgLd8usqfWFvwbLdUnCI+Ryt+D4fM7uAWSkRTQx/yV
SN34gAu7yGrUg9SKr2QTYhgwgoKKLFLKkj1AW1kdQ8+rBcR8v8CntbO7VMUnNdYOxTvLW3KjjB6O
FW6cf51PSZlwY9R81wIalcPS2+BnXCvnZ4aqyeO7eVJ+ymyc46WGDRC6cbkukiry9Mv1yp50Skxd
8WTD5bISRhK5dEuGdncM1HB2YQVGOOBVQAuGwzIAHxk/RViYYgVcElmQPQmxrgE3ysJvIRRm7Leg
SXczXZtIB/7P8XntEa7T+Z+q7L+0ahW7siZC7VtcDF8Ki4Lp4HTTkUnVLSAkCkMJ7mBRZyEmg+4/
lPUpEi7+NwuRasYGH8toNDCuUMON769s4Yd/ebm3jYccPY1sul9yJxzz6Rjrec/OjDBQLzjSL2xQ
Wm6eZN8mzV1bcYS+Q+MJvJ09a/yAclWVnbc2DzLhyOK+/j97jMdnPgoTI7SMeEDRJAM9bbq9neZ6
4PbYUcVqncbL5rRf6tKXMkgPuVwZyuLHGDXFEiYhh1TfaKbMgtDuQNgW4hKIyGwSdO18UPWMNYGb
apJEZQxPgxI/n1Lw+uWKM13JrNDnQROyX0KR2LcU8oGThCgqde5/qquMMtjHBDgdK7SD7mW6PV3j
3ZUPxq2KmpHXaSW8S4MtUWG28ZYzLrNXNGJ6lI3gkE87jpkRjVMbJ/OomORNMfiphOdoYpNDq84O
OAfC7NJTF1ubob6vaF3FClvWB2DWqQndaQxvsjO8iCbeW7cFZ6wLw7N1QMnRQ/YJly9HDjCa+5/d
TvPdxlunxFEirRIB0exXiXEkhwk8EUFc6E3HGag7nJ/+DpTrOwQ81ZNdT+WAcM8HeapxtpQERiYs
ywP/WmK5JSu60P6Zba5PEeqclWuHw/KYW9pl2ruo6dBI2yBf31Gi1YsYYd/LThLZ4VwBuCe62oZy
xqb4sYk4g7HJg02bXPAzglydcc0fsyyJ1fpo6UX1/U9EKBAuNuhu64Un0UWwaARJuO+yBoLkmA9s
JZa5BMFKldR0oA9QVFwZ56xSKaNLgPF2eDlTOClmeyyzXD9kCWI+8M8OHkWlz9Z4gwz6kp/Z0vvl
17VPFdoMTNUoyubXkOinsdSCGic8AoU3xoyBzsoBLBXp5TbFA1yVI9Bba37Q2zcm6fP4Q3g2PKY6
CcH7ahXSEsqPhjbzc0kXvz67C+TVX+ACvR9Pt/fqwiFmlcJ40EtfD3QiHLA4srqMyxUNc4/USMcr
V7VAOkangJLrhzQvGjjfYTYTGuonmVjLp5YeVL5Vvv8Jf/bX1Ux235ukpKolAOg1p+wGOWaLW4MQ
xknd9Uru8Ctf4vMiKBXDg03eYVynupYUCcme7pKmpEqQYQAiAZaQkLJWQr6E/oo+BZGb6iAuHwGN
qKltr52jIcVjErNHs5ucBLVrAj7srYLliLz9Q01n7pkdY956ufQlv3M/SBFmnYqgWwmSQZo1kV57
bl7mUkIHWcKl5YycLylD4eXsjXQbJdkQPJC2wCZdrcu++F7dVL4yWPQCBHv/JjGKVD4Ef33W/wZl
70ZNsOcTqLKnLTd+VScG5mp9p0cg0oSqDvo88BjS1T7TvQYWJWaw7MkS72pxGZSbHIpeKfKm0dxH
D+ylxWEME0NsQ/b9IPR3QbLyxxZ3B9JnjEwNyNEwS1qFKurBJF6o+fzu+wjhAV3mAQ2jXpwgVlOk
sW9yaxyK2xYiA/TEVoL1+p3hbf6Dd+SZXsKwWEgV5/jD2p/fdE6dtJ7ofW9IuN3bA6jDSSaxiGJG
roJ63tdakwvUgvBycci6Lotsi3mP6J/+ByJ9U6/ahqNG6vT/r740D3vAywcSn147PbOxMl6wXN8M
cEkoxWxX9/BSiLeOfVKvCpoiQ9+63fJy87KkYVDDUagsl7zugltChkQbWMB7dDR46bo+/tprFuRc
KHy+c6PqghDMAgnOK/jG08uCzGzsgR8KYYaNv3r1AtA5YVFvvFP0orHQ3YxLuEPUwhnNOIr9XOm8
p1mi8tsDg41PXfB1rtJFcjQ2TotIdNFSwtpQ6QXTezcZtPXTu6w5UJlbdvoW9CfQw5SbyQm84eGE
RPyKl0N7HAk7GXWisBRJendZB3+3vJxqXJbPex+T8eo8WXnE66WjH3R7YX3vsZfwRi96EfnujO12
stophZTFecRuHccDTEAn53Z8k9Cy4dspELz8CKO4NATpGK8pVN40JRO9QG9IIVgmKE3xXruJovPO
UG0IhNyELeW+TzLAXDUe/uLqa+Bo69AefO7XyGtoplPfGE5GYqljXJNKeSq4oIU7TrG5gW+Bb3+X
nZWaXOE8buCc5eJSLJCSQUJn809oL57XHN5kPEauy78TKf/TxcVHHXmW40RsOTVGdBg/Jfm07yAG
GPImZoIk1oEK5FDTM+RYScJQmz9gsVf6Kkz0r13BCB0hJQX4sfZuxtdR+5QDRBJbAuSMKxt1+GhH
O0Z7obMIwC5Sp5cQeuqWOZ0+Cy9KdDEbhtZBTWVDw5FGI218r+PjnUP5mAx3j6/12mdIxcJ4XnAk
zWQ+acgTnhNvxWzeHykgT2hdTpDIoRwb58K0qvbkKIhfhFByENs7K4aVBY4C/cO/5fJ6gb2A5l0H
SRrurS4KXjM8cUX10dCBncaXFWzvoQS6kxPlDfocTj5OAmgEKMkc627r+REQjAzZkHabjt4oQhYM
EALm0iPbgISr5jU+9/ePXeW6R9vanKMFu1clR+Y0nb365lLBHz9QRDCcNaBqidY0e053IRiHnAe0
lba7osey4L3QrShIOnFrcd3d1UtwkFRWYQfhwJ01L5Kc4G8rWUN3OdPzkKqdvcE87dZ2KkoF0GEh
gVwnsXsYL258XMV7SovLkB7jftEyV04B3qKHDRODVXwL9sdUFYP4b0fI1eUuDgdEF1TFUmGTQlbj
x3ZtKr1VDhK4vtULEamOb/B4rDWsOLkhtWkkYvylfltTGHAbfFQxNCcr/UD0JFhESrN9jcvrOdxK
zgK+ghd13FgJpRk8OH1+1Gtt+U11dyO6t1ONOJqIzBaPZ8jmJNZ2ZOqtygUFwg1lgIEXsojDkQox
YTMHGIPiDIz/M7mut6E7Y+0ltv4+4+mN+ctUMRxQCxnDwsy74ENRaXEErRowmtwb4ZkPBSyOfciu
jJT14elPAk19exg9YRVs19G6TZN9yx7weXbfJl0uiEQAtA+oiuCdAx1z5rDuZ9/oLZScNdmkRn2J
5wCFczFJCMhhmv8qugwohuDqg1UzqtWOC/hvJap6aj522x2s1A4HVeLHgmHUm1nfHdJW06s2b+2Z
U5czYC0yRcWbr7ywqsWFpMj2B3ii5TJjP6yxqtaHdcAYADuWYZUpI3G5+k3Xq26e7kCbSQOETptR
s+jIRZYkLdB0nkCJGWXigukUj0MfqaNU/nhSof/7mQMDdft0wAIsyki6sJb6jpQsiNAV0QYtDOrl
UXf/yRaLWX7w8GUp57BMckNg8Ti5jtdLG5HDnurMompwEXn0F3GGDznTpW81EVx7OquR/m+fY7/+
T+IZEnWQQ+bvzhxwRSYN8Qub8/vkwmhZxYulOEFJPAsUEbjiLohwXzV/V9ZgEKEej+20I0+tBBq2
BuzOg/LRzhSZpiM+b3CjJM+/WSBD7EqX+EYInZJTP/BtVBKAqeoO/QC/UcuSwKryLAs10Jhu3LW+
VgD9vDf9HJTOnu4jIm//a5zfpKdOAJhzoXGqTKQx2qv9Gvir3l4Cpxl/IaFItcZmwsk1BvMj9QD1
qIrzokV75nhW0+E/jCvtAziv90AgySTdrv+XxTXkEor96Nxwwe4biTmGnr4xewTHre8cyf9uqK52
wrbqVIoi3PuBOxi9uglqBDIZB2Tot6GD31lX3nyHZYvBPlwXqECaS8YkTMZSxYx8BvMk32Mfxv1S
kDOHgo18a0VQIWThN1iHcB3ZKC1oly3fmPz1ODz2qKX3r+hT0310s6Hq2okkFc6F+jPTi1LB5EC0
WCQnAnLt+9EESO+qOdmXuCeBw+6NXhOnzFIYbCxdwvqcUHgtih9nMJSpRdFQMxSV3IV+nr3e6Di5
36ENUalJGj3DkXrHLfPQOeWUcllxzRwcNxh2MmBiyyVt+XyO4EzCINILQ5voogxfd9Ftg8rH1OhX
Yk5bBMb3C3aHsrE+22iYAY7KfvC8n4ytAlhzMFIBk8AOOO2+y80lIYIDxWSk6HmXMLhY8tXvYj/8
OUYGUNqDUiCrrgPUtjS4LkxzddyjQXmjOa4Wy67KwyV2F0gauuKICWAGy8/VXnpUtHJr1tzM9jUV
mwKBa0aIKLhLUHkuWFBWkF70Uy1Vddv2yJq3IL4pDKCzmljyoL82GsnYcVD56XP4XldJjgLU9u0F
HDZttUU4jnS8ZzB5jspjMTXQy8d29a2XblBQT0kZRLepqhZK4s/aZK5gg/sNyUaRgMVHK+xVL4nQ
K9FCnQTO6eaA8Y3W2NwKHG7y+bS0dKvV4ZIGotuuhkAqLlFDxh1K+IGgwlK+Awsc9U4voufPFcHE
GKkZ0fPn7owCXTUSMHiy2osNVp18Dhfvj0trFH98k3qKHJkZN7/g0i7ytyM20igmHNp4oLyaeJyC
Aa5HOSRNXWtrZMh1igFd/CKytLdc4BlQQ9ot2Ih637RZjGJzYRU00WlMBo9Pa46HEwOSsQ/R89+x
toijfU9/KXqQUqBD2n/GGqu1yITPh9HtXlQo6r9M0IUxftHO0ZGJdgiXNHpXYkLF8VcDjFCRRdoK
yx+Lzv2Leezaw79yDZr6rQT/vBd+sxyftgzhttcbuAFjo1K/AqNMfyZrvB1l3gCkSmGPjQ2vhsDK
xe2G1/RoLoWK5aVhpPRGqleB4s18bnfXjQ2tGZ9aveBAT11Jon0xNz8dus6Oz51WMbmr90wCmDZA
9z7IaQSpUXHYxjSS1JX/PsxUU+mvePnB9jYKFGOy7n2+SQXGVtmCKhbAzS7QwrnMresSBq+uA0LA
hAxJ5scHI3O3ffnezZT266JixywD/WJu8l9FSLuXtTeTqjsJU1b8SBlKdaobNbzZsyTAhSNifIKc
2miAgLq04bhM5/jfGK6ysnA2sYSmcsdub2AIizUdxFPoI58cUEiIHhyU8eTE9R/WUVqh2b5qmByp
o7uKCz7kDRJOkCDhik7qjAM+nsVQJ+sTWXPIHMLu+InGlbtGfVKMZtICBuC/Qe2ML5Sz+MZkcMKP
JK/jPSjGjgX4fSKbsC+pOkukX9Unx9dNwgxcVlUn1OpdGLhFicQ4y1qGmI3FeYdHiZfZysBVzm66
fZqGxMc17Q3dbYTNR4b6hx9xTAPRMmDt4iDbE0VXbitS8lJWWKgALvmsC6tQJX6ReGrAqERt/GKY
29qNh2dDxF9JL1qfu5BskNaJqdvx+eqOa6wUmk3kIEKQE8snyiEQUJeKo0rlcvTeC0xB+6FIadn1
a59ZtSLWIzroBOf15wsTwAmPM3xRocOPa9Wm9GCC/k40j/ASBr5UTuOGQv4ufcWFotIAtykvlPcs
zBcO98tCHobGGB7BSAxYW/HNocdprlqho12kHgIDj2O47K/betrZHHg8R2ZtdrQdyND6orNz5VYP
DnfY1Kk7uHYmCLq1AoerQFdH1YQFP+hd7kj2gqS1mIxKRnZvtkSHImbkh7U5Ehsrr7L3ncCkGUOv
vwwrr/QY/374dTFJN0X/s8I7C4WzWlMjZGVTwzMRvypaNsYIQfmwSUL5eksapivHI+dP44QTfASq
hX20Q/8XashnONoL1veIg3ZonYudrF3bGR6dlJqMzVTUeKR6mpb34TOIBWUtI32+ro14YJR2MUdI
RseDb8hkiBEvSk5yL08MkCApDFNbglybkRrYpzjhz97galXCpYIAmNofzpe76YQTl2bUv2wZcWq8
pZNkUaMxOaZxqdILNHopn8VS2qp0dsaJp54LWjd8rM9twWTwipfN/FbU0i2UgbyQRU2QDzfRx7eJ
J60blbq6p5JySpO+MUky+miHTNCnY3qGK4m/lgZ6YbtloRSvewDrLgdZZoylMTnDDCl/2oVTOIzl
mSvL1SN0z4ReMxQAVj5nbfUSV2K9rR4SStGpeQ7RQf+cPOuX0kwQgrGqRWiWwp+gi3Sl5O8ivqAU
gUazTzdn/+1f2F1FaveVz/pyie/xmO45AWMxobX6gdJ96+0MNy/P2jze7z8Eu6o/qcJa0uUEROqs
9gs0dgiqJ35klFblKwSWCQSOTTRJQ1gErjcqeO+x+hguHizfikSv3R1YeQAjBzrIFFLCQls3PlrD
U7F3e4a6LcmhGovfPRvXwsLm7UaNM7VPh16WPAQRj787v4EwVYDWwy/rwGr2mzPjGAm4Pm6KJbes
iE+NJ6pEU6mQfYnf1UanR7aEDDcC3RUM0RTlDkPZby4Y8MaPr9dF7ar3Dx8B738pp4MbNnQr6B/i
1vhVXirgl8PDTRAALcL/6rhulsPcfGrEL49fh64716YyJiKVMIYjgYD/R4zgGJFYaRF4kWDdg6tl
3CTQVeKNam0pIy17Ue8WJegXiUUxGc3laVzDxWsafwcdvreD+sDHMCJ4XFjAp+NvQUJ8de16Ywrs
pw6Blh8vuJoru/TuN8Ptxbj6UiAF1edWHBQ/qTOtH/jKnMbtnoFfBUz9dJNg99hsMHEvArPjJJ7U
T4II2wrPf5LNwH9gZxJTpobqF6l0SAeD3GlpUWLDA3Hg/+7eCI/QWqp0zKaOWr69KHgafac4+cZj
EnygU9VLiPe6LfCHEKumiTkbFF+jXeyu8R2+3AkslpxJPwqntTU1nrdSC7DbsF/VXI00gvtsV6E2
iETbDzvospUnQgarwws+qvoFlUqyuBJ+xzQoWD3JL6jYQyQ/rzet+zApOZGDJ6yKE7xu/ClRmasq
G+2mS2zClTqDFDuARCRLun4b8PlFj4+mwAqOQYIZgfVwQf2NMu6PAuhdpBZxlrUpbm2rPJrUJh6e
LYZStrjeSFwyWYtTtRdEoi/wSUBzYlIQq0MsqWyQHUuWYvXE9WqW/+MwUL3GbiWzmw0Y+aIrssUf
4dlCRqLR7skv5TItj9CPtxDdzmIs1/sn+LJUhB1OpzknKPKlSDI0K4NjUkm2ZnLdTuburHqO4rVK
5+htgZIaxkp5nv3bbzznozIgRHAG+EKAHe9nsr+9ikVC77WijAXkxYHNCLyv08Br6LNMgU0MaJCW
dqkGEWqKKhH9IswJwV6SUlL/tHTEcmIOcqbYao8RsHcxGxTjLpc70hRrJFOr1qJ3D6V7jgkZNpKh
JfmN3rK30zU1xJPueLxPRn8IqgnBIpojY367gm9od7s63qjiae2lIPPJXwDW4+F0E11d/5wTvwQ8
+R5JoC60vsJ0YqmW19Vm8MJOJ2TAAJsSZHauYVjcsx5dPyMo3d9IsUACjJMrRlBrb8V1JgCpG+5P
JmMUVzJycP3dEskRyyJKVCQqZFiptyFtbeW/9bkGCEpjMnBhVw63OZI6trKf1Hpuf055mHrIAR5r
RmMaW4dHTbOxgxqgHfXUq4E3N3eoGgXdmBf3VekYpmtc/I3vMt6/s97R0fTYVzOn15p2Vqhp1nLC
mPttXWD6FL+oeGJO95SyjT15S5E5uLex2wOyNrdAjVQBNIZVi5x2541wfiFqFJr7g8SX7l8gnLR3
y0lA+XBgJOwiiiKmFp9COGHh+mPNPs/umAr2FF/d9inQzoBiJ4hIsPiljVXD7hB5cogeh7r60zHy
mJMEvfWnbyPKkY1X3IXggCHLtwie1bW5Xhv4U+cb6Vcy+FuyTFU4JPc5iOK+YylAzG4pa7Nh3HLx
yYWZaZrfbwnSWTN9BUnntyNfaKjn0bCNc9JR7AcSwO+UQIpZgKHow8v6x1Z10IySi7aS+nkRoM2x
jurBsjMmS4InEqt6EBvCUV8LR8BUW1e3nW3YTgctYJT/nYGpEpGi2Xr1Cdcc/e5aGly73ivKnZV5
Ik/pZzwJqNltTHPgmixzgJo8jJBFC3qnqxxdY5l8j0yutUriU04gfnjltacRpgg6UnXeQ3CU6CKI
6eQdBNVLveW4i3C4bKocvCynWqYf/oyaGli45u5+ZnXOdk8t+sECxn27L4KTHsz0HELY9gEoEbzN
NaWFAVsoBfd5c/akNmkteUoZGQdIkIWOq1KKr5YxZWve9J77OclDyoSYuRZeV+gHub33fXbEnx6J
d8ceUgoPLEmWANV8KborqDjikj2fdFIZ9WH5UcTGuEnI5Dh6bQqvwt/1HQOWsFO9yLWl2CjhgZMH
VzFj4BKUXv/P1TIn5GnUTzBvvkb1rnfiXtN0TLM7hapSb6NCoHdOX4j0Ix3j+5dsQ3slD8RGhuxx
sIeEBe0zokNSuIHm/DVgFUfbvQKcQi+rtpQGIYbb9Z42MjR8jpiFXbsNyCamUsjQkBoWiib0+z6f
PXbesepau5DV5xizwKhwmoflQboQM9Slr+PtLnTbzFk7oelooQt1xJrto9c8RftUuqI8G297S6ph
GzMREq9wnZEhyAQAfGrJhV6tsk+bV9smpb+6WkWXTBon5dyGsH1QhFP6m88tTxTJK7eMbB8HxLmI
sv56jG4sp3kWmv3/Bc5TaCEER1sVJg95H4GSx6kiD6XOONQ2IgwyHJOD5JwGRzOOMJ+FyzT2z456
UHAdP/IdyTRiJ0niBxwCBUET8lDlEwdhNCil8tFD37Ghbaqixf9X6KJhPqxHLyud9NNx+XF1+EOK
aq13MThPu3BThJYw6dwwKKtVy78I8tBtHlIdZqGG5ujO0YqbIZNUSDweUHeqAg25SjQAmMsnxHbC
uvNN4jJaU0nASH0Jit4GM2n2eAdd1sKJHLnKpHdH2PRI4/KvG/cearaE4XEk8LlAuyPkIlkws863
JTToDPnF5nYaUJRWFBFCYQbjMJspw6xB7yrhcL7pifXeuDHIPCEASZqP62jVQNAU5ssVHxygygjE
gMDt1lLoO4sZpon3Qk2GXe3eSGA6Qx2ysDN0fM8KLZqJBd08olyBu+qh69s4zIEwweGgr0X9HgdX
d6sB5vywvGJlbDJe9PYL8bwg3HXnH/Nt1Hk6G7KGv5kIdKIdbjFQrBkkul9NfhMDdAI+38TqjCTM
FfuaJU68zoXoALRVdyz6Y+uH7LcAQGj9q0H8YY3vhu9qxYyvcnmL0Nvqfu198oySrwBdP2chcaGT
/k7bC0nivBj9crZQz81oSScRuMOBYJ5ACbGHCxDckzpVrLzI4+Iqi0KHWYwIjLJW7mOmC77yT6S7
kdwidS6bLVe8LtFZMM3kI4kQ7nZu3+Tn2xHdYdAAl5KSsDPyYshveDBpPWD6mWtWV6TR6osqI+JS
IP4esym37T6N7I2qX4BaC5kIu8sE/QPzPnFmS37e2E1L/YCZp++mfxYJlhGzN1naO6cVMygf8fDr
dnql367RLJKVFsXDRgaBFr6IQQvaYZPrnl9UaZPnH1ldqKXM0amkjeXRYcK5uxJ/AvCX5wwAXbu7
DeQHCGoHqsty1zGEFiEpiIPgM5Uib9uQyXuoCFIeDA6IyMhKgtReZWVoNrjOcbL5X7kO4GqWDBJo
EgNqhRqW1DQ1I+pgWxfvGl3Pig98PH0o/e4EDOmGAykDan35M19L60hUnhuU+fq9v5Nol1+B0slk
gw0fFleUBYg1sfiTBun8uQ49W5G+mPHn+qi3BMridV7KHms2DURmY5FMRz8aVDa178tl3waHr7LQ
3lPuliLIEkv8a3xGGlr5oBYMedxDKWI/unjJB8yb6eoPFajfu8m9a2iZwuPDKRmz2heNdc93IGt5
Ml+zGq9bBgoxm6UK1sUB15AZBLsh5pGG5IQOnm9M8HLt/wwDlMgazL3XHtIRWuyFEqWQ3cVga40l
K6gmV6zkBm1uRmfBR8KDyq8MPkKB1d4xi9ATj76xEC7uYDV7hvjOSL5DiMCHmBL5mEih6QbZgdcu
zjgkTMIILXNKne2BaAuptZlbiP1P+c9KJfuVaj5HA0wuZjyvDn6vULrPbS6Ln0VIJY2vn7NCGQQb
rdTiGEnxojVGOgx+a83dWYRFv8zE9OAI7jmaaeYLdiOOxfuaMRwkbyJK/7rt4CWR96olHjOf4fIo
458mNu3GnTCq7WJ+7eQJSO848S/9SeocKdSLY8RrmZFIRcGO0APR59v0jHz6XyeU1ozVLcpJmfZY
79MQ3H6QtkW2iCp/DC5qcyYIDwSdtsGAaXacxFHbLULolypfO2X3ue/TZr1yzvnrTzmjwfJqOQ+K
rotp7L67W+jDTjqKmNXgh0Q63Xy2Bct1GwnbwJZTcMcEjiesWuDeGourn91capoB/gRbFi/jDHWe
a9NgJRhOCf7hEqQchLUfF71coaLbHSRqaS2LtALc8pHBdnJNJFENBIXfxdNTp4TuyCFYYOF+lOte
3D6m1Z0WDBmUPh/MPdStovunQ1q3KXbRf7RsbUPslxX4yZY+RhaotzwcGgEEP50xqo1jjQAGckg8
Fa2Xa74qPPIaU1q0Izkkm3KUGmXI+FDF9lqK7PYLndMSSBriopSy9MA+ICd/w6Zv4cm5sDBFgvsE
67PX+eL3pjZ2PsSppt79Qtty1nCCiyDj4qaDnTuaDXSJvPX+neC27wHn7skMnwEfkDivk/DY/iMY
GpQF5hizFxzTejzKNPTZGcfRFkvbdCTHtwGkKuQvzj4xnDIC7yj8klhqqmO0K/VYc7TQwQLhcBbK
x1H63QlfEfPdruon7CUkCWGrCg1NtA5ipO9bQ2axD8/YlAssls+H9E6i8M5eqwcSpbnWW4Uw06AP
9CoZav6+ujcCDK0GDXnx9B0rcRgkCp9KWROj4t8eSjWPAoWzFvHPn64sez1rmn73RMExhlRmDb8K
HZQ3Vto8oPJkTd6sod83daA0oERdRB4tRmSFV5oQIYu9AlUI2BFET0w103uCV7Ivv0zXhLSGA2oa
2K8ladsRTyZp0q1jFXdSSkIp9BYg8D+gYxTi0VDsA9bnDJ1denLnbVVolWMb6VromLjmuuLJod8a
wT8hDSOYyanEI81SOmEY9ZOXEbW5DJc+6NxoRaUT8SgkfvwudPQWybWnQC4rkjpmcSEoxkUXBu6S
q4q8/iEz1aJBW6DMKw0rsf/jAd29edrayJDVhhTuVzv29d+Wj1LqhfrrUQVGssrd004a2W8pHn1S
iz3fVwZ3/hzjCFtO4li9y35HCu2EhONhQndXcJeJYrJNQdQHRRIWanFxuFhrPqVlT+O026H1ZZds
iLvcSVVDzf4SeGTbuL/hi7FmeH/aSgSV5evxcnw2CrYLM9RDujbXnJ1vYyA+BwAYOAiwAIQHxULp
kuEE/X+3ikMRoYycL0LnE+sI1EOCjA4RbBYI4R3ShG2OAXF9w0PyNV411Ploglv1x5AsV12y9pqr
9QJslY2zw0IYQluAtx1bxZFnw3f37wWN63ThEPG7rJQiNqmQ2XBduD3+tkCF+vyn3DK5/lbDHG9k
CvMowT4sh9skT7C8E8VBj0Dt4mV79cK/7Eh3rLwFx3WmGuJUP1c+5wylPgsojVgKnTfFKGLmSFyb
18hJftMzsy158m9pS2v+6+zArALPR9fuXA8zW6s6QhX35QHE84tqX0JunIHlm+cLv4tuWI061bjc
D5w8xOFh6yM0opXgIoXkt9+XX6TUS1Fc9F3Msc17TfF0rRhZxT9HYllweylFiHj29rV/Z0gDC/I1
oEWXXu+GKsg9EcvqRzUdlsQBMLUSUHyRdaliPlHa4qHt5AX8dazwEkWzsgLhaNn9wMVG7QcGqaZ9
Y3xUHp6tkO+6LBWeU4jwBgkxfIAprt5RcTPiAIXZD49dxNtqcZ0fRMeSgHh8o1IgM81fcNhZsnrQ
vL3hBMANwMDWJFhSR5QGtepDNAJdoj7iEOqPdMEMofmgQklVjdRMNk9DljzzzTXE3KdQyuI+9QSO
yHD/ub1Z33+w9SIQRQj45kG+MiRmATu6R9RlSe21F0qQpkqmbWkkkPk7v96F2rY84SaxJRErEs78
Nm7o9V+3mkUtRXNJqkukAoJhGkB84QA/X0fw5m3HsT7R+a50RZD3FHcvsTXFKP1TI+kMYPx9xPfl
pHOEA9WHkhGaPuIs+cu8AdjkJhj6FSFExCisGfgoHluSqfYxv3b8g7Dy392vIpawe1oHta9ohVIM
797OwwSzEpDjHKWU2U4Zww1UtJ5AwYrmGLbj6x1H14ukkrLWSm3NjSKeo1btegzez/X2u4O7WTRd
VJDmIpdznCECXLTV1bp2KBivDbdDzZIlzA0qCP6MIG7YJmZSUpdeCqLzVqbDsCXyn7RaVm1WLYhK
dcBf5y1cRDbvzieuchWgr0f6Q6/rHRYTKSVy2Vm0j2dwcpre+KG17aDVpCioG+ot7T02OiaWb2XG
FR7V9/lP/hzeTQGx++zUQeyubYgbxzn3V0WTq+7sW0p9vhHuHTvQZlLk0zO8Feyneq6r1BkBK4+w
1UO421EDEGTVHbXtG3N6tlDNQi+WSoxEUSvzs33593bpr/in7v8OBPn5cCUyAS0Se/apq3YuBipb
x9xmfHiGBxfP0zUdW9d/iNz1GhQRzD9KGCgBagSKdoXstLgRu8crzVCpmyU2zVtzQzf9DFuWve28
3T6lBQjgTXQzRh/2euMBxEuE5qGLq+nkpcdRgfykC4eZQrTJR+DAogccsH8M4bKz1QK7j5yxmK3P
C2Heg7gIRRJhlo+kEhrHyYbrpzWJzN0v1IxZZ9ZwlavVHoJ+CiOfDyDlpi0I/fwsFQz+vHK6XqgY
syeucPJxHE4OeTE4HRA0OdN5cW60CZ9riJaNfnrQ9MOe8AXye7XQOEnrL3NQT19urJ9lMpjbgcNI
3Y8k5Fy342MnyojXO02P9Btg0ISLiFD7Vj+jpQrGg+LNWnefqNYX6mmrS1JoWqVPnaUu3KKtB/I5
WRkY5/f8SxRy+5zVS5X1cELAtoT5b+YDJpoZftUpD9XqEgU7vG+Eo7ySaGNkknFwhGAV1hKzj/+l
RtoGulCxUlVVoXGLBvA8tueNST8pq/NA/JiC/MrGQ4LlV1tz9MvD7PhKS7e1aLGxHFvFitlOGWiy
Ai2ik2N/PViy+E68X8E10/pWIedsHFC4H883vkwU+dKFoWybM9rYhGAKLvltTUH4qLwb32bBBQm6
jvxC/IYikt7xWAmFkM+E9BbH76yElUenVzCTKTm+xg/tWxfH3b/R9+iZp2X6qWUui5usW4Hlgi7r
3NUkW4R0qDxZMAuXlZzQogznOyCqYQW7IeD2xw4s247K2iDOZ0dU+aPlAQ32d1tTPOIjhTYQY0Mq
SdPDL9u04SfHwjkC6PPqD3iNiWR9mNhnAxW4h+Tn1y56ThzwwVdGfbTyuzyGRLGO0JgL5UVGZIe+
TlHmP545vQJxOKzcqQ4yxp9jMU0ZLmUTF9Vbw0pHnge0oxn6c+clGIah0iuVRxkcNbykhnlPM2VV
HNWbZXd8UMTjXc+Rk8su575IelYAkgp1UHSN2DxAkqLbf9DoMfwpkT7AXXDqEHYwvWEyH74k3JL1
eGLDUOvwxgG8xECzox9sk45BlN/S9oPf8Rkh733ArshqbmP67ou8NessTJCY2ptm2m3F6iWSoqfM
8w4EA62RZkd9FtabL6dbTuve1aQKh9z1QhjwfBpIk77lAyUA9IgMzUC1ajltCybPFG6KrVIaE4Fl
d6NQeLSK4HFzsQFGOPM6FFFhGCylRpebUoqwbVWQX0wT8QlGztEc9fHy0K1q+RzdJaStqj+Y1uYa
FBNz29rLhCD7psg87bKytEf26KWAzTpkRiyLyqqrEn+xz4zy1ou1SbJxBDXrG+T+iInsqHvWlTaB
B9PmpKrtskrquCh6PnyU7WOZad85nNvwLPLZKXmHHw9jQLhYZOzoNUfWXrns8/dmqp1PfbI7ZCjf
g9SRSMXz/SyYAlGn1lfim7Oaq3MeKVvsx9cMvmeLfCjqMWp1OI7AwB3qaoSUnTmtzsdcH3JeTm9I
eciNXYoXZCrPpE/Ijd5Jm0061rF9pm9UfTW8yMusgsj3rk4PcOpbuay0G0CRbUQa7sPdy1zWOBb2
zNHKqvUMmbXGt2dEiOGGqK5rmWKABOFBXqhF+CdhsBZJD63N2lnOqWVIh4M03pq4BjjZwxz0r77p
uIuBgHhiWX31bohZv+v9U8Sa0tz/q4oh+QPbzJjVXKaS3NbjtQO2cg+a2ADVb60677cN53jfyOvx
YAYlAUqbi5HJeW0Rigtn1Aqa34Mc0S+uRXCk6pZDJQNS9LN0z9i4QltYuqclG45TKGX9Thky1uBO
VwUlkWTmP2t4G3QSndHN/c6u00ocLML06XXnccfp+n9pck+6NKVJI1454OK9L8aYoF/AdVRbhp6K
GYPYvVFNUA8Ir6dZkE6ESAC6Eh5vyVo8wrd/2fZxO90zligv3RQmEnfh06Z3bkQGzSeNa/7o/M2/
vnh5o/5nlbPRdCb+j7ZdxbihJzLgYplKYVkILrA/xD7NnKsibWBZ613GLRQoJaNWSrGLjiT0of6O
kpaJUhYWIfOu4J7kxCDc4saW/FftZBpqMZb0QGyJtg+STP+nlLazxdzDoNpHeNUlHy0qaEXkeROA
s7IhMk84Fcai231TXdIY78ePaN50B0a06alciLfxWKS/EhqdwNGT3S2oSzIMmQMDI8pzY+/k6kiy
E9J5w4i1yRdrWqzTxungio4apDpUWYDxUvpXUevN1vmtF/P6GSJpUISS8srxLfRnNfLNBCeyHBR5
lXzJRGU0uraAHuXAcDATv3G3qJUq64pFaA6Dyo0Zne39/MUofa08iK90NcA4h2NrNggZjlZVpsts
QVCBAr1aDCcxNKHfveV3RenAVSbIJzmga5p0GQqE5oILx35OGE2YlCBKCPme+JCRpx3omCS5FM1T
g/+BKYBwzrnyXywyas5HkpQlin9LLZgTASISTvA7JMY9hMsymubJN1W/6SNM8YkuxdRWZqR3pc1P
i3SIDp5FpRrK2jpiEunxQ57V9m78B3m+GsECwDupokMGk/p9jKOWEF9ZOTIjwqcsfZIcqmhbyNIR
ndy1XeBsuS6gNxxOMKjelpk7oWJfx+L37dicJbXgXSuh+MYmjZsCjcgUQw6rrvkJTRU2T4JCwDO8
cZzUFdlAg0LBUrVBkvaEIthwpSKMKPfvneIWQdXln5oWIinnW/WUU4mrwBkxjNgXz1Qd6LRsuaL5
/yMJYNlm/+rhjtNvwFv5RZzZHW/mTReshGlRPGnVlcFLtnWJ8Hi3NSPoM3mHACM863RcPGr5XBu2
Tkp8AM5SgZHijC1QstWdbfFo+X8jE1jTbu/lLyrfEJZ58mSYGj5zwZDXVF9eWZ9BgV3RQhrqS9Z9
fsdS1GT3FXh/tYHGryr3rOqX2SYl49OhIIig0kxxggh6+H0TwXZ/4MK3NS0vabe9n0ETjpkX0j3j
/R/Xij+BYgck+7TyI9CmWCq0dQaz9CumRkwyUfaGoEf4OcekYGp22XuuE5DYO/NX9TaMIZal6GGF
2ujJV11f7QvaX2cNmUq8wPDOwd1G31T3NWns1FsB1bEU+Ckkfa1MaVd4zPzLP2ekyh553lUO1f0N
CN2bsY/eqcEYwsEpRXBWHde1IIMPBVLcy1eW5CqlPaeeYnYYnajiABsAuRPaedxevlXV9myV7j0i
aSzn468WFzaJk1RniEUQGWoWcfFUTAlmizZZID6SqqCqfF3dt0pb7tW9eapzRhyduDXUeTeYYq1q
yTSwK98S3blYISPJjlnl4R7asFW8Qp4KvxupTW8Un2RcC3ux5M1dMkxZBf6DTX2kvweJwtCySmYk
n0NYWvnzZz1XScA6iblNccJAU+Rby2GDB7wRQAOmKiZ3Sib1pOCZyxXz1ZXc+H+DiCQmExg7aXjO
tBBNokJZlo0ELwcxX+2Abr3N8AMyl1QRYweLKiW0v2+LGGY6wHB94HfHYNFZYdF42fsx+nazmT4e
L5W36A3IjUulSiA2KzRn0hgJdovNyrG9nCrnAuzQPlOfCBF9kyf3Xuzu9qDa8IRVRCjvNTp8rn8m
nodLIwb6KWk3tWd8fLIbUnFQulK2eWKAZGWCIAWskqlIPXw0anT/KEffeWfgtFzDQvtfou4+qGA7
Zad6HH8ubekRHgu8VrNqII0w7K2/YutBADtTtCfK3VLoK1jl/wbxQJ/cb0F4fxNEhm/cr5HONbCC
xBDP9ocsB7OlpfVOiAn6pE+o1TqW0lwEn3FRh5qfzIujc+MgtQJJZYPlzpe7wCGuuvm0GCiwjwZs
cRsIlJ5hqoJhhjN8GN6e1pFWBXoOA5JmgteJjHwLooj8Y4Om+THW3UX0GWJSeApul4qwVxM6vkE3
1j73oHy3B2HaxelU+eBkra/UtV6O5TVQUlFjJ+ntfFObzI4QK3FI3NHMnl5p6qlR6yjpyBzFEb+6
oYdqlWFv+gYIUlmRbEHqcEJvbKwPT7lpjtyynA3hTsxSNPbehTBn9t+xDhG6jmbszHeoFrCjw9S8
CMG061PtB6Bn/qyx7z2V+VbcKE50g5LhiMUD4oiltZDQ89gVw112g8bMZDiGomtyuirlyUj5NQLW
+gZiFaPuCTJCV8bdUszvwWuz07VzHFmvL0XTbMZsD71F0XWhKHjY8ijOpzvJdTKrrlKb8LFWhkAK
GEnWA7pIDs8h+EFM+taLA/FVuXjH7fyyRIMgtH62w6wWJKT8jLj0HsSsoCUSpLAbXIAMPR/M9vW4
nsl96zW90DVl+il7sZjmovDHc23Ne5nt9jgJRePFVZSh3CzORMp8N2De7KJjUv9+xm4sri8WDGh0
6kONViTlM8IsvLsv8ghYkIXT3+qkKwVqNyX2UUrOTZJkeRsDGYngqSsUbd1UQOcydFRBNTi4Q9kj
FRFsUj0pZICsxDc3h9PxZW4onmYp2gg/eCZRKqY+6ZW5r1bPa//K0AordKxI85MHYEfr4O1BZkI4
fea1PP+L/Afd4YqVxWNXeqcdeWnC1Epq+S7k5fVTcqqJqfESgFRGqMbnhqYuOJAqHZYUH5HADgKk
1yd0BhFrXi/kOxZ9Q3vZX5ZEwtiklrFqZ/QCmbm8eVtrGKcjgeo4IfPg0owZgu9giuVWurUmR4kO
8OwdNNsaSpr9Be6+NY0sxr+MZBnfVEEyYEmigg2/lRSQedJnEBaND9kvArobFSavjZMyz23xlZfb
ErzOf37IlIyRigtEwZh31zM1RbLrKjYcesMT+aFDT5xLVIyhkIiaYe8tqg+O7RbM7INjgBjKsVSQ
zaRrrAKt5HcWr5eLEuthmBVEOGJ6TiFVa1J+TC3dSWRR8bhn6eiUeTunP45MvX0LGI7Flr9hNfW9
Y8fzhqo/2U6bECQkgmx5kdDHR689b76GDMJZFlgZZFv6lueV+tGufMAEJyMWChDD1j/BBHySxNgE
Px2YSsOI+2D3rx5DIM/QrG9BVRDBPYzoR7vBRqnOuAh9NTXHJ6JfSxc+ePjwQzyF0Ldyei5wZqwS
Lug9LEh3fRD0Yql9noL8ZYgvg5NUMit0G9s+pMDeYanzUfXSHpqVtJwdMam046tAb0fNH2PwEPK9
wKOsvOdC7y92neAal9O6iJoX6mWpwraKnRy/FiCFecSypSUF5Iu4QlmB41NKgNi7DdeztvEKV4mW
MPzTMBHaJPlJhUaBD3wmfER37OcYcSBF9lcC+1UxFTIvqXNtjSHMS7qBxKHPDvFHzh/t+wqcyERK
/Uu9l7XrDVSGMY83QZsCChC+QRwxTzSV4c6pkcPTKwq/CsTE2R7j0aCShWGLMevQjw94Lob1ZFiH
/Z0rzkomNa+JB+elX+zmBZDx1X+jLLFPePq83eqdVbiN57ygWXdLEbNoIxxQosyriSN2+k8XK5Jj
v3ybh5BTrk9uYi9IseB6cJkSLuIZAXA5wAtHMywfvQsI+6KkSKjjvxqsqjy88FQ7Ytz7TOSHT/XK
j8rN/WWf+++wyvbaYqS1GeK1aVayrElxcebVpxuwfnb+rAooi3ZNXoa9QnrOW/IxN1OnG3Joa8ya
ZoqXHHLznO9SqA069Q725OCeuct0hy8SKjYFFkX0WV0dHbWp0cBpS2MS3Tela/B8IRANk8piqUeZ
P+1TCi1W8fqGNw90nuSkp5IwGpfAYwXybkK4ZLWda7iJY47eZDxqIIkq0wR/5S5CRHNISV1syzEu
PDPYEeSW62zk7Nwhyt0RDG+hXY+bgZrbJcKEJ9c/6+J3jNPz/7wAEd4veuG11xWaKcqYik+pHeZJ
zGyKBKzxHvQYDNBb5a7GNejnpBAnBDWb7dqpuCl20xBmPLWmmZ7L8nNgB4Ski1iy2jVMXE1HN8iA
JX6XiekN9dxZi//TRdmFyOJsZupDTDDvx/0B+08c0pQ634D6zEBBesQlzITtEgnYvgohm2QXi2iq
rtHYNmzj5SXLf5bP4DGJuELqH41rH0i+ZI6CrOiI6JkPjz5DE/y5BBAlVNJYiwz9dQO+bWVrOHU/
7MO1VZJNDb+EpNvqDH2tE9+zgI0BhNo1gWNW0+CRIJo3mpdwASvbfxGo0NdMzF4uLwvfX/l1SRaB
5rkRvxWyvMpzQusRVq1QBNduAHWlKWKrKhRSDYEfHko6cKLqF4YEcgNd0BqFR621tBZ9WbKOCb4x
LXEL+HnC9Kzo9G8h7ERg+OuF3w+plIk3Y0hqJy/c/YpzlsYdddWig3Dtb0G9JMjmw4eZfAYiO53t
L8K8mkZU2rfkbDDrgtgrTxaQ14/taKPnUdkKKNWDS6R3n3UZN9FGDYuAvT80R2JL/RATsJAiNdVs
99SlA6a+AC5nwaKB1UHAJR8niwe3Qx5r4mdBgwrTMQsAyeeRGIu2t36/w76rKCnL9zb3xxkWbAUA
ttpApB1KDN2dn5rtMliyt++qdhQb5ArHqNsDdNFTaQvHkmaG1GxtPZoL+30nO/8AnVk9pEAzSNZh
5560JBbvNzvQuXX0W7Z/OchCgZGe/Et1EG2iNuAra3iSP5yPmwlJGmT0xgiFkXHfxDogfuP8p8/z
eoICwS566jGEd58DpRiV+Jvx7iomIGpjaXzfoXe6sFZafRVLbA5Bm1SwAyN52ZH9VLZrANK96bGr
G4+RQup2DDFeOXO5dJftugpOESVO+q5t64qJlbNx1j8Uz62VoOxy/WGHYH5VcpIcABZjuBA4EsZu
ZL/F0mDledwMRwYsReKkTeLTSMgBczsI9Asw8p72qVDIOBrW2FwAd2zomYmWb3jIaM5Yy1nLA0h+
0JnwbtVum8lrk4XUm9e24pTw9uoWIx6IlTpHfigxNNyEppYzzusebP6caH9K7d+pAigz/qVD+E/6
3A+gJjFhZ1Zaf0Vzl9SkiEfzgqGUte+t0jtaRcyt8im40s2mbqCl6/a8v5KuELipQw0OgzR1p5Ue
kXPPNCcmOOfTLRVE4Z6w37CPtvI/vL3pbACHvWnpBJRiHjnIaaQU0CPAx838uD9RaA8xBRPk7PJA
XdL1smmtTQda5TGroSRK25kAGU1hOrrmDOL858pFmPQHvaW/iZYaUCFMGaCO+iQfkaKv6Rgt636H
L3irQsUI861i8dO/htYoTX2lmUgc5QDRH05y5fUqb5LgAjaoanbQblean5UJXkEQDTyOMJfwWojU
jH9xZ8iKax0/j5NfVNlH2cuxQBKq21feHIcu2kC5tmzxVSqyQCYzkW0PrOVRc3rQCAXtfUfEx8uy
oGmm5vCXHMOyGnVQvUbdalCjWiL//8XnU/1Hz1nYozpZcsHDbXdBhUQp4Y77wjhZr5rHR3we+jvr
YdxFAr0zIj3KuolbFFm+IrOzUGlynAjIu032hPB2Hy8ZHDxF7AE0LqcT1iF2g7dTIRwyf9BUA1Cs
ewllyozs77bctIk/FaXkYZZfUC6Lsk0ul0iN/P9OBriY1Hbdc7IsnvbTmwuBmpOu8MxcLKKw137i
JwVf9lNPn4agyaZP6qHNsVNhhUXqrPWlbmz7QInhizCOOqx9xtHVQ4P+LoqSd6IUvRJKAEL3xcGk
N66TVp7xk2gxJ+xgR29uBGHWYex/bj8bXAUGec2eQnKALbRib8NwwBdhdBPjp45YXY3OJ9aqqEtb
RIHyepcoBu/9Lq3VhF0wduUsghbtUQceWqj+ldFEgs8p/T8PD1p1DFjOE1SoQbwqLRMpl8lpp7KU
LsAdIzsc4++E0axBQVoLJ7Q8Krc/mVDxPeFuy2MWvR9XJ0PFKeAIguN0T9ZhYFBAjhC5/RswLej5
o56A1dQMdRIQe0vX1fGYJUU+BaYJrQ/xbIJc2gLO8pWN9tVAD1MafyFFIFT5coxhDNBjaxfDhvGg
XDghEvIX+t89YQClI9zLLClNf5kOqFwCmCQ/vXmj/sXvZSyOVbCBjivaCkWSkH6Q2PYtckHCT6zx
eAyAXXMxoDlh6Trs5UJJjoA0ruOK3KK6ZVQhYornfMP/CpTLRAbwBywAkqNESR27HoWx0rrcRuBR
ZY12u4Ed5rG9QDMcDmuqCDR1k+niLFku1rv+6g9mzfAXKrUUf8KdJ0W1z+IKsxYQKece5Q4D5SM3
HSI9GGGj90TOdGkb2KWJNy90EOonTyG7A6ADsrTDPaxhOrVtoKhwY+hpLlzy8o1SzWbUEbhrrv15
Hn0JzTZ10xZ+73G547Ddy8T7qYyBfxd3VZ7obRIuhxI4+aHPtB4TkVxThY7HsC91pTkTc9HBg2yG
pRlDC5IlE4BzkR8DOAQDXzvIjMrTBa3wjbIGso1djsJzd1tDgW79QZ8hQ10mw9DhR3xqUiIPavzj
mxbaicOYwh28BYdq7TZtfkpFwVNspdy9Zma6XtL709gafHdfKbCYfQETlnDabtpyuHYHno1qVSIg
nE7CP+CcSRaK+RmvKTNd+ZQVWi6OpTRO0xWkUgq2VBDRSF9vS+feuplik3AYaTcsFzMH1ZaYgZOR
lwAKvBubvpNIACpQJcfTCL7QE7zxUCfa6M+c7Xy6g1h1YVDXB5c2Sh2c+lBIWNI8KKGURxJKdDCL
fhew8GWGaaEL6OD8Dlqm1euhtjooPE6lKi7//dKFpEISS/TeYFkVto5P9ev0JPSEOirIx4xBlegf
/55J4ZY7SYRTuF4lr+kyKHkMnzR2mlS+hmDPPogMW9VJoMJ01YwnckyVE61bXnfUcaHvdVgyA01n
JpVhNiNeDnLF5jX6P1A7qmL7cvOdiOpJjjr3l0TsK564kP4VNz7xFog4PB13rDKH/U5bQ/HJOxbO
VQQjLoLoQ3lgNcTcj88d31OxeMprQ9jCBKriUh9q+qEDO9e+FAOdoOc6cSbdXFPyep1C6Aun5TSG
JKRv5TtW+eWFqNhy2WUFtGNASBbR9Wa0zrktv9HajWXNqlxl2AhLGgdhgOEPw9X7Nl+3wTRW9cLl
TBtlyxalUSWJ//i5bhQAKCbYCVQ9MMOztqQd9LcGXcwtfAbqYbgP9/VE/z2S4xYHpPARhsjdp0W3
MDDi1D7KKdEU8Yy28w6TTSQyEJeBIIaJXyTNqi1H2o+pLR+9/COQZ/o80oYo4eZp0GXhCvluheza
sNorAH39TPRNck3/uMq1QuvUV2g+77Ej6OvMi/Ky4VRm+fuAB6m83ZfTUkyAuVKjZY17MqFYf/Um
QMPQht+VdBlFNbN5pCJnqxFZSOfw+KrY1ZPNhSxE0gXwrAVRBJHEh3qDYfiVHyNbMSd9m91AL5tQ
y1keDB4LgFLPPgrckqabYlierzxq+ph1IoAbqymgWo75kxD32ZBXr4qayzqDZROaJJ3gyVzCoqE+
zpg3P+rDZzn7I8Q6jI941fGQoURNZcmis8b6WDT3MQFEhC4Z4cUFwP6mR1fEeMbzAx8unOjn5XfW
A6kgK6iX1ZXQWZ8ByzA2qUss/ag1n1reWskPvC3vkruw9nOPx/4NUygIEMZbQVsjuWnzVD9hJKDn
zbVQC1eI8bH7q9bdaUc722v8D3jdFy+RkP6eebIKPssZw/YTUMt+gQq9c1CJ4vaWGvrG84rTlFfc
1vM0LoXzwyZbl/Vx+GrLGmKLbThNijFst9bogADgkySxRekpbffi4SR1WLPUf+Odrx8Y8LDq7o7d
DaQKBoHYmM6EeS9xlhv10F8XS3xSQUPHLU9i9TEfoZzoFzwHfICsJ/84kfb2FlTkTi2oNZfrR1wh
te1bdbwAmIsrlYA4qh3jL9SOMtKou1+EkXaPLe3I7YdAyv+JQq/zQlKvClcTjKVviixuF11/kaTF
0CkJVGrYSEeSqH8DkXSUavxnP6quwrSWJKDUzB2wWUURTsMR1Hb9TT1VcPD1CRoXTmg7HIJOk6cE
uuxsfGdtOKFOQHsOCy5ZSDtwqjxRJiEKMD0qz5PITUacLV9epZYQJHgLKwhoQ9n5cqiz/JPSfdYj
hTVg53gGiIciZ0JBnfNJCT1ectppxB0Gqe4YDyH4UzDNaynGfQw2cnbowu+KhwjO52vhF2L/4LPK
muJItXl9BvGnZKKXCOwCMWSgBMWMPAdWUNvJYYqQUTKdfjxa4/sZMD5nktRXXR9NDt3zO08qIkv2
7jodAinca9syNGsj4IDDLFA518X8ofaFt9JpMQOGO7rks1RTmaPbWS6gTtzZp8auIaUVkXAh3ZG3
cGn1xgy7Q2rC8FVc9l5uvvCywxeYAM3uQvwDBVZVaToejVpVAJDwYRJIi98ypKx9LCWS3pmlYinf
czffZ95CEC5w/zWKJOWjd8ZS0FnBUc1Wm5uo8OvU65ZpRQVPeV8b268F1GzBWiuMG0GIe1pzins5
kLZAwQYTsgkgN9e6v5A+09a4Vx6fQxr0o9Cz3Z8wWu65d0RmvXTQ07CwIBaN2y39Ns1eEnCjRKgd
3hjI3iyvGVKbMwizyC7jJPy5unGZ1fUQzROYQMJe+B+QwK2DRP5pZTND7rWpVef3oYt1AA0m93Uc
rbdFCX8duClClc8aL475YKRhXEJ7q9F77qQSMiGhNZi8xxDGCYwP5etqgIZMIcgF1MXg9U0k7JTx
n4yys+cYaAnBSrpQW5PYDHI2Yq54PV66eNCJuu+CiHw3xoMZyJTfg0HQHhdpE9IP3ULYtQVpbRMz
oZxcpP6nqcKAGeh4msuVfTqifAOsT5jhqyjQW4B9sFGe4ZGPiL6SPnV0SWwkAOloMLmhdLNgTFbw
ooX6M4Z+L+NBeFBdWKMWDcIrVdeojhDBZzZDcxfBl2IJDL7iW0JPVAPdAslyKkQ1eKzWSFAJdMxp
vpqF6detVUBFBbg8vuFWSA7A85jWqbU/t+X3ML9IeI0vBiH+GNSlpLsBtOQujpT3rOMQ6MHyj6jr
XX3Dm6HPfbdSBStsKBb80z+iAYiFYjeGgepRznXv1dajVtcka0UEOnlk4PmcVoeQiVBjEiLUwR/c
pu60oebBUG8wdYqadRSTseCfrkAevTZv29fVNP9E0qOl1jHQcTyo9gpvGGyqtIGgz/praP1au7Hv
vclPPDxCGiVVuIqP3WvIqCMAQRpEYZJYjIC0KfxwAoQSWDf/M6r7IzM40FP4iWB9L8fbb+c4X0gM
XjHCzGdfdotedFhtmYQElFClXAoyb1LDWEUUr80oQ53kxqYggQguLG4JU+v7voxD6jZK2wfi6c/2
9jOhBLWfMpZwVoFxmRwHjXmLjLEBtBY3QV0nfCJztzd8qcqMSjuMGh+nK5ktRhUtUM5n4MBb7PTw
heQCuCrTy081RILYwNphuwY9sugn2+9R7mhF44qvU7P0hldJybptHgY2VUqyGQWlECrOzmiLfOCx
62S298/LWdDut78ulhXkm7gXuw/fpHHXDFgUZeRQlEEROL2v/ZFfCbXNZPTDLPDvwhi9HrgU1cQ7
LdBFRJz6zwF08j/jeIPUfbyfGDUgaAGwMnFE82yM1ROaxlmbKB/S1uQdenhQwxHWL1LOePaghyqW
NmB8iAjeb+alJ9ZgDOW7Bgs7KJ1MvOGb5PbjW8eP76rkiXmjP07evSfOYqYrbAVgmvfAA8DgWKKZ
zL6hgCOJu41nQ9XZjAd5XTGbd5hf5PhppmF8MUZNHqbuMp7y9gK4t4KNK4NOj/ZixI49iB6GTr1T
5pDY/gVs/cpt2CUdnMGm3vhOdodYb5SPnO23As02fk8/io+d3CRUW1KEttCcbhcx578rXwpY0Hdf
y+r+NmqYk9MFmOmQKWpNCTh9YTQbPvA/rLlP1nbMlbrr7tgivq/wAl/8q4tr/cLVNdHSTHlUgiXv
QgWO5q4GyllJaeIRj9QS/ARv/Wq0cK9rYXW+xnI5OvdIqfUOA31e2k5sCbohblLsbOicfvrtr7kD
lhIiy7tgwIxcN7qmToG1nYAtHqxoO15c6F8HRW4aDGFKv3MAIFPjrafAfyO82fUa0Y5aWJn+QXhW
uEtTdz9ryHJp0WulDGr25mWoNrRLrxTPtDJTybxNEo4oPM8mi1c7jXL+Xe0a2FCLioxJXC60jLFO
ocVFMjxULwtQQU1gZWks7PhygchwWUcXSMNufJ3ocbcLvpKjYG1DAtppZEDqa8OKgBTJ0rMGYHUY
U6zA97UiJbTvGUjEe/EZDaLcSdfxm3wcHH1Soz9u2EW1kgyxx6vJKKjGZiiSZpZSlXgSK4nBF8jw
hZ5nEmpMKucOdx9aiwuGWlRJOsJb5Fnw4yXjdZ/JSyLIMFMS3nH3M7G0lvxQg7ywUXvdPN8BzK/t
cgLXCjxXB+RUkc0BITvlORMzsxbFUy5Fax70Jh9nqGEWCcXkSXy/PPVNTWDvjKe3gwD2ZWbUUqVF
vKeK1I2K/5K3IWL4ubvOqYwT7S1r0mQKFzq+MLHCii/9f/ZzMeRohEuEUCehi8r8EueCw0t5KfqM
VZkyiSnV35J5gwZRNsGbq08cnTEmJ4yEu/LQhkB9m6qjAfB17dbhtXco8jI54zqTZrHTrubdRb2w
N1+BLSdHygPnPaNY61AGhR8wAo/3t65201/EweYV4Tzm6E2J14q2sJJkrQ0X6sQ6IuWf+1lJKhuQ
EsSlCoza/jwqxuARlumwuMHJWfiFUvtwz5lvkF/WRa5YkaZLMS+lGFm2/u7YAu7OCn40sRQMS7mX
aTZu2dQnTBIB0mi0y7rHwlQ5uH/vBbihdQOaUwelHZgPoSrAM3X6zkgNp4uDG6I8l76LPwnRDOx2
7fm8hR0EtXxaTD9RaLU+QI1l3D2I/ZMuYzHrW+e91sODBVpV7yERiHImU2h+YRCrwnj6+wSMcM+3
DX6ilL9L37zSwHQ8pmxsCDjKV7BNMzHoHL9EcndBf6+vj9Ovape9Za8/dP2KgsGPNjlyZ7TvNpdD
XU0Bj9L+kUSNm/TPPhjnqXnxxlLBn+vpVh2G0bvguhy7aebMHj1Klmz9JeKXxQN9QNp3mobFeJ9a
Tw+Gt9rSmRI8iMm48y0cEEsSHdoNxpGq6gXKLXWXANCZ8CDSQ46oxL3Tcg4olmiOA1QCoUlkkEo7
0a61octMrzD3VKgZKjGZxC8+ZLBqg8hwjRhKfXQPuIHJj9fHEKiV7FxoFPOxvRxvlutVxUfO7Mlc
Dm5+ZieksJ4P4gS0Y+24xyBgyQbD4PMkoo/yTEYs84Vq91Bl6yFBnKrguaUWu2XoEs5n4gG/bBLv
udY91u1Sz9RNuWTKBMkvChZQlv064l5RPnMDc4NyXuEWHnWZqFpsj0j2U+46NoV7yCBoC27fSe7F
YpAsqIu6awUbx14TYXJfPRdyK5sTGgmf33GEpUu4PPifCBvXvaVblPu5ryUbeXLnrirJK5v7rLrs
2IwHcfzckrYcYiDoyJs6uPOl0A5c+I3iVbbreXkUGRyN1SNNkiQhWqCyDUskXMMIx/FM2tvyhupn
TYmBb5f/n4r4uK8Jk4+XYNNIXK13tbXvzeIICwiOLlH1sxsSrL+p1qLYOY/RVgOrp+O/PlTDhjFe
cOoUFKZ7V5C/2e3YUcKRFRpwtw+X1m4UbOFPvA0p9OzO+vB+9fHJ5vJDnZCOib3XbZVWSpCFah7S
weSlJHz9ucxDBLSbQe0s0rJ5a2qHxnPAKHDRpBE42UbzqF1w37GDBv/2Tv6qHiQGSCSHsp3dB+zb
wEDbap0kfY1oYRYiLmHpWp3PsnEGAMEkKGXidfghyazFJQQ3t/Gs/Lq1VLK2f500iH99fCH1QQAs
+fsxAS4iP4ABHqxYAPBTx8scbE1TGJ4sYOtX/TPhItr9K/66QTqKF0lwbV1C3zlJeDzpIN/7NK3G
+N4prf6OZL6WKiiZPZX5EGq+LKI0eZWZQkOITl8vHDI5/CrTSc3QxB3ngxQQceRQtoxeluyLjKxX
OWuLCiG3o/+LrHnctOLt6ldjE52V3O9EGYmEhc2IXEmK7z49neB9h19nar7eNoi8oPRsMfJZIWzR
tRuCMOhIuurrdY5oRgKhbT+VwjnomHR+dyWYgohxvcyFwynKqDs+NGUTkz8FDJ9Jsbf34gwwYr54
CbTtq5HEbVfWpZH7BVmG+pMVJGu8JN+B8dJH7ERFNCHmgu73HEgTlAq7djK1LDmvWy0AwPgjh6ei
/I03CwFxwbJvD3iBs1NZ0ecLTt8UIA8A0c/pR584lcqUWT9+UbUfazV5XkEdAxYksYvsGYhfl4+q
71/wujVtUot0FMnWwo2lnu2FeOkfv+GheJEGMafvGy8noIB3zGMq/+AXQkX7q9iq0JZTkiE+/Ceq
tQtSKYrznnODzAFFih5HjPjkLz+U3aoKaqgERqePdL509aLWprgbnTtpS3l79jrFYqXTi+Au3t+J
Z45/f6RCLfMRQ7O7vQM1ulgUWzE40m0c09rIsR3+HgA8IIzxGGYkraULV3l5ezxdAjYPlg2cvVP+
qk3O45sM7yGOBFcpjVu9MNmrwp3wb+HWypJ35sgzTj9eczNnOrk+kjrQuk9c2L9sxpRlbve9LTdy
GhehiXSuvDk+7fh2zq7IaKDJ5k5TYZfUFQKaNSRbi/ErRwPcPWxF9qd/P2TgrbTLcF0Z5jzpzgnR
VgK8CBjBGZZFYBhcrT3+Vn9L3Tja/yZdD5CnGH6WN1+emq8l+DVwqYOEtspqIFztbXXTECGPlzMH
g/5xRT1+NrR99xt5VHNjeKufw4fgRmGpJ0nAxPhOHZtOvArPkIDzT0dI4W7zP/ht3KJUr3ST920R
cDwTGoxDh9vnlGIMKt4qeiquN4HanpLEO+pGKD8ifvU+cjH7ga2PEG8223apSqqQYCA79oF60X+r
aPrDvOWlV9yEN/ybfHA/wPJ0g9IYybHmGOMiOZTQRSY/5F1sITrWVxCir+KRKcKLxxGPAzfbOmzm
dofmEmksLn4wHia4eRjaXdF3Ob9IgYGo2aXEdpBRGy1RgEUHaZVZ0QkRuLAfqLs60sk7Q8W5Kqvy
I31KaPTKdu7IcBne8LaEJQ4vaT8fL7o6g9QoQSKxg4DvNDvDSOCk2POAMr/EKzoPk0+kZ8nZ3Wje
P5jJcTXTOzSD1mrBxSsYqvyFLXgHu0h3xnABlDCfXEwui5VJRWaMxyvYkZaJLkG2v7uYcXc0FGcR
CYkS44D13YAkaGaFqv2R6GF66LylDvG4olpOuQ6YS04zk19KtG91qyBLnA6KmSnyGOHo1IGyCCQY
Y29VctslB7AjVFfAM52JlALvxyBHNeLgJdzOkPBYn4TRvZaclMfzE/wfkaZ1Cm9dzvE4PZHtA5sI
0lD/9F6OCderZC7+2EMO5Ks/nk15ckHild/XTEIjsLRZ7M13JY9UI6Z2aOA5q+zgdmgPvyCJrjnD
2mnzaFTMCsNB8z0o48T1jtfEopBpEvEJi0u0GIWf4aPaHm/1ViXmELlRLN+zCOXEaB8BBl4o3rvD
y0IswRwiitny8JBpqAmmGDj4B6YZV2oqyrVK2FbHt8sVfqzf5zCkN5oIdyDTOtjO3gGF7ZCDgg7S
G7paWUKZ01rB7CDJksu92r4fpp10owXfAtPh3dJdYT3gbRdrH6bOvQ5IedD6tXKPMtrONBcJzuuU
Y8/HObTXumFtz7nPZ++glsZh9N6fipdY+MX41fv0eRA0B/vATKfZ8p1QNqrpjC9WF9lbJ4QR1L6i
4jxEMa3fsijTovXaD4OFqWq4uLZpVaVAqMd884zfvg5/t2pKyB2zOjak+bZLkANBd/fqKy2wAPVB
beRnMTgZq/UjdKCJmyRIhdfnvajMPaL81wYgOBfexE85WI50aDCN461NLb1Yf/oh/66C1laY64lf
sDs0vA2tc+Bjxr8cwdM0uSoS4NdkxNvI4BrIWZ1Fl/GWsPWN7BSRUkdLDXDEAu12jAw08KiJrpMY
2AEjlIQ1GX3I6yKjuM6uexOr4VdoJBkbyd1uILnoh6GeDfF2Q3uWDLx6X3fxUw3jFlKXjA4zji02
naj3O7tcitCgX3a68Rw/Lt7uTfjMmHXz+OnXmqJbbGn0YFopj40nd3bcn/BU1Cx9o7wYuHb0s4xb
r+hRVxL0ywola90RgMyACBXd/feCmfK2O4G10iTvvIP9R7bEL0bY/wsjnXGoBgCDNUE8hXfRrgs3
Wl+gC2Yh3WFJUTPW3DQYRq1B19YZAEoGsVjJXACt5fru4gv49RS4SQvUygEl1HgxUQTpF7x16j9J
g4z7A8g6IX4A0Cp3zrQgcLzHa6J3ZOnNJ83KTjY+QXh+keIrNQd/tJvCt06qoFV1hAnUl/E/n3Kx
0ohGiN+DilJ/K/CQjBJcpF7QO9sQauN1dQQ3wtBm5jrlpGAq2nBSS6vGlY1m0/iSdT2PyEpykVkg
sY4XQW9RQmkPSINydQHYT8/pq4pQprebyzHKn7vveMXpkwSCJ7cQepJUjneeIb2I+fKihBAGVAZC
3BqcK7ISq+iZbqxo1/ph7eKexsygmsBbLCPt+bIaFGjerwMH/yF49n+p4kgMQEzsELGmio2kGRiR
1xDGBrNN/V44EdSGG8iuVE9SgfGFiYFquNKxoW7YCPlsiFJT1d3AsMnhG5utvS7KIHkL4RlkiULp
HqmgSatJB0bwBoA2HZZIGMuYSIJTeKnScfw9LCDgP0VnbGIh1Z5AZfUkGAbGwJo5RJHDWaQl2eal
qOdpSJfjy60hJK/08k3pc1sOOwp40v4oPG4sgzvgHzz65sRE6FVPRN5yDrJ9dL2mnpzQnsGccFra
GDPgLVLRyIMbLaTfE0qB66jOkm3HZ9whnOgjIcwfjdXQ/PFgybsSu9QgG7hQA6y07HwkP03iCz4W
FCze6X5JhLybRk606XN9vX/6Hxx4rqDuep6XPFEY+drNO6tDnLzD2JYwN32U6zF4qYUnN4XzReo6
M0jnWE30DSfNUwuZP/RNyVkvihHfYg08Zrvue4OK+zupa5IMzkz3g76EhSfk0idbWy31Pq+LEaXE
WBc6YeqiwEZWQjWgJoRoQs+S8wjs4RvJ2fswRUPQBWabc0dBjiHpJPkmebVD7V7dx+I1ht3A10zJ
1uN8ihNmho35LMpyIGmo/SRQz8lI1g0lYUUoTDTd2OZOjkgE6vXDSRUNEGlzrja4LQihObcEk4d0
GMFXr8BKxu9EV6+yOWAMENj903WMTczR5An7PnPE3zQMNhlS03+jxNraNWbwhh0PNXdp0aMvvxdx
u7tIFJxescdCaXCMraJ5syNvICIzdVT9VLBabh2inDo60o4RX2hhImc5kka4aSNEAKz6P6u8ARf5
pXPTrBcS0oWEhfVyZkDgR6cIxJaxI10lZxrijgw3+oM+b/oZkJCKiq761QQqqyEIaBI0gKmiVv2b
vaoH3dJ+9NO38REtL3TvO/w/922MzUMcbq3oXh0CLuGKutKEEzMeHWs6RO2kCaCykNNXgCp4bU3s
WU0FYABL+W22/KgAtoP+LJ/4DN5GObb8uCx+4qIqfQjvuoUGQdOLsUOFTseb2LS46fNrSBJmlO2y
Tsr2qY4ItzqizUmMzhSb+oW8QeG+xN3/uMeW+MjFCWzXrvJ1FPSiST2n/Blcnhk69+zKJDZ8xtJ4
N+BrBS1Zjj/tWMaib/WdhlzS/hjVmT+V2LdH4XxmvstAt5jTOrBPza4QCQWqq5eUmyfYnrkITumo
dGDW1M+XzTyH2HyGV/jxzniWjXnBHIxwcO7BHpaCwoDyC0TgeTfNgbrPz3/crw/T1EwGndjgUNjS
vQLh6j0AvsX8ZxA7SVPyh9Tf3F299fuszjtXMOxFOiDGpDR/37dzEWC8/W62O4CKMRQ+jOa4PXs6
e/RY1/dYBarcJ6JKL0jZyP1DSc1s1/65AjD7RqbRhmTSX/IRUdVC+w7qhJkXR26kc+4ySb3oVdvk
b6FISTa1/di+H+McyEzoJERtqRmw8Ib+5FMyTKH0Ld/mTdINgR61jQJLiDOGZmtrbJFBNqE5+g2T
kRbTfpa7btvVkeSma1rsIqJ3zLWwrLLOcxexdkiFPtJSRbk8BrVTs+454C2ilWBy0RWj9uxC5kjN
X+Wk5iH49nfBxwBGG2VmDv8i7dswxEnrs8Tyq9WpfnoPwU8QayOBQFUz8h5gk/hMntyo+RGn61b2
ywC1Im46Lu54gpyyB/kk/qu2UJG/nxU5n9Jj6z+NDLE0t93mzkAnHd+0v9sX4zDfn9DxJnhhbcPJ
44lvC1FBreI41N106i55mwX8lMpw6GkMmiKaLCBm5nDZ5Av+3GWDnZv7zQ93OMqrXt7HcUmE4zKY
CCd17DXz4TjTvgBzb69O9llaXKtijnTeZ2etgr+QKLVbBO8KDjiQlfEwji3S98ehhxhHOwIoTXq1
MPEGL85Q3SxkVHt0iHQ8QhUBJo38RDYQ/uQNMxBS9wX8taMtyfeHT8NuTGZFCzhzMdcog6UkQaFp
69tPiG+Z030FQ+omtFOfH5J1tenxl8ELBz8LrzKIqO9j3hnY9OKt8QE9HvXj3+BnXOa1NanSAf06
6xkqDyLu5NX1dsqGcS/YqFHPmAgyBw44IwGIBlpINuFGN8ceFS+LfCIAjbXzIT4hGTVuU18J9hfH
ZsH0GCmWE+MnlkX6cV3SAZM5xPfNQ5mtV3dnevJcVWCrLWEi1+LsKRLwDJy8czPCqeU938dhMW8Q
4UZXvX3ym7CATtcsrbahcW1Ti7WSnGo6r8BdNMqwEfubyXfdftav2uuTyLgjpeDwCTTVZrP9KFsh
W6lD6Mjce1fhgbGjLBya4yMYq41A7G2f4OVPui9pAcCy3rEwekJQcPw0whRuI7OGkLH87kTqnzht
SvNtWFZKq6rng81d+MGRSulNphtvjfBxdwojHLw26sxzvUV74mEsZPvDY6IA+eSsdP5pHf5rpuEw
KVvDM1pF8dJ1HaJS2vcRtdzJ5+7noz0HQythg1ha34iwd4jKn7Xc0JNt4mBupdZOP0GKVHbAhtAs
sXjqtmYEEHmVheR//K5y0NkIspnPSDPE+jc2hQHOoc0ZnNMN1ip4v6f6MqUGmM7HXNBK4cJjNvZB
f7Vj8G11nx17wCu5f0aFE08nz7B8UaTuzJRP9egZt/PoJwERJM16aLrXY0wb5ggOFW7ZuUv7boJL
2Sp6efY2XVuxYp/go2DQ/RT5gvIAmieF0BfGxiHASN0rS+FVyVlSf9aSJZ4Ob2Qz4hvE8Udhpd1C
z4HPvUu0MHvJ/5EkPxvV69oGukdVtvdVbGhCxFbSMovZLcg27AYuzDmUMe3LB/qZyABloy1ygjXY
PSiIc5Bx0lkNcM1pg4nQ3UGROOoHeKYkpgGGyANkMLa5jfEUpPHu7hbsACboW987xJz92dtuNLdk
HthPTdFeOdHVpw6Ms77tnZzOHMmYXLfZVbYRyyS/xY+atfOQsI/V0G0tVkESsDmUwd8l+E0D4Z4M
hTYJqUmJl59OQhzAUOAt1XtVic6prDSdUegMqliQz4j95lJQjpzApgNz/QcDkaYpTiLjG6+PeR14
/gm9LHak8BpsCF3gygdIeu94nLAsY7yS7oUO93/ZHcPayCQH6gNdBqfIiwjcClQRDCC1sMgbCHDk
ZN3ILBXtgie7lJNt1SaCfepAKr+hXKLyrWUFrSv9PLzesB4zGVaQkt10j5T01us7SfpZI1qA7LB8
RwCKpt3x8NgDYunlacaBrhQmlIZQzxPVIAeCZ00eDqpKr2/MvuWbgPgKoeB12dclDsG0m7OPI1wI
BjNvZOV2aUOkQI6FlguckJ79dKIGfYRvE0YSlz0sV56BoVT1iaTDpVmMPpL+ptMvQdoAfpFEhsw1
ZGqikjBx0ja75bOVMVyDriHqTScZCYS7fLG2UTiRAAhJsAhPGIIL8RuJr9+5WmXvcazHZbR0VeJc
qiccfeQa0VI8K9ip3vDMymU4N8XCvooNzVCcMuW3ioMpeaU9m77Rnkn7pel09TtNBMjqIuTGcZn/
72ARPHqZpgbqPUNmKYQHy7hkqxxQFA/WN09ZhuhNuTLJBNh+5sGufChPz9O3bPDL9qtfyop3Q1IJ
DpDFGP9EvcURoyAnOGlPyL0+meyFZ2e1aNbs7ohP10ZJp2zN7tV0M6Tg+EN0wMoyGcgRLgUs7h1L
4SYtY9oLge/wfJYOFdfpHQcDtCT+npXe/mkUAnPygb4GQ191C4rQe1Mj/s4LRGuYq/v6Zcigg0ZT
0L6aZaw9UIBXM/325pUkLg6a/Wm0UAoeWysiZNvU4Dt2m7uY0zbNJkxKRHasVG+X0jxNOdlHBoDG
JQt/T0JTuHGeBCYq4Cm486PiaR7dlqpyEMgJDqPwcLrUKePmQ+qP6ylBfb2hyd2sVIEwCBhEfS6/
+/47bafueXE3FZ1D8osDAAjVCpYG/yDn65yolS/qv21tyaWRDFjC2SUaThx9G5gbbg8035sy5VMO
3RcGyTNZw3x7PiOyGTeIDwaEqPNCqxWjndzL25biys9RyLCqndfuPnniMi5TixLQX5KUAtXi2zL6
lWQGRY4YhroC9twaJpkkslR+xITGj5faAOtZzA/0ch3n2WWJ0cd7CGGbL+jyhClqxHnGmCK/yYPN
EIVGqeXjonMFfsbaLObVMOg/06sgYK4AChgbGunrn5OLFsnQNzcH3G22j7HJBpsd+SE5cnhM160R
DVFIwb/+I7FHJA+3oeYBaf9qoIbnmQ/DSbtBqCpNcP2suHMBJkjDstiGpgjf36MVOvB9TEyLqy5H
s/IyhMmdcFBKviMNsixsoHLjQ7FYCQt3yQzUbbJHImJSjazToN9soy7DIRWJWV/Hr3zv9shbpMRb
P8gWl0gbGW6+QevHYXTQ6dfHkW6ig9w6x8Pc5/MbIdbpsy49VUgmxg/QvXkAlSfefSZuKdRPT5Hj
ak6jQavvnXXwKsJot97CbQscUFCb6NTSDhN/MVzg+WNDgRZmUP3JJ3JtNRqMjuApuB0nFNJjhs0i
kk+Q0cCdjPvZAfNMg4BL6cwFEERC8NqJc3RN+Tjs6x87a3NKGGgoIf9RBhGFJCl+tS7L+nFpeT5O
CMDXspLK4R+w6LLpejzGCPrGGUhcIXSrnYWv/8tLX/sx3IEraQT80m+k8lbnClabTWz4PVp1g5tN
0kR0BaH+vPUHCPNrdqiJPc+oIzkAvGR/76BGrceK1LmCAT2pWDCqim2pBfxMhVNht507AzrQa1X8
heprenjLU8tWiKbZ6WZPXlNVl4rKtayQnOBlLwHJgoTCJ7GHH/qSJzODbJEpcz5U3/gIPO4ShRRx
Hh3J5bl22RE2Pefe5A689OfASrMDpHz7J37lACv0yQDSr3lc3UnzVHeGucm9w4WIYS9b3XAsXNtJ
q7p1p7OrFIbUb88RkZukCumDATScOHyLJCq82k1DlQkPTmjhfepEdteeTlposq+n3RDNapg1Ffbd
DFkajRM8X4mJ5h5dt5emz8oAjaSPQLffcIqBEFy1PeIBbl37Cckg9HwDIIZmVDuAiiN/OieuEJhc
zFCdeARhC/DrYD03oIl/GZi5QPconnFjb54FgvqG4kSTC1cjKGxum7l2H14K3iJSjjwsZb3m0EnO
TSrkimnEvmo1V2FWC0lxGM8TuZVdUJVC6qsqlwn0Zo/aae/IGkOhnsLRtXS/ZekNp1SsUMkDXbaL
kN0BxKjhSB85+Feg+JIOPGoAIYdfj54zEie9QU8sIhjGDwDLRcRSBekCn0HAYRkUXJEaM/0dbrOg
c6wA9whx3J5jEk51AEW0YIcAkirCvUW08DF6i5r/OH5eosKvwL/rJj5q4vSf5p0y0YWkZQ43qJyb
QYbi3X+B8Yc/r8UQF6WBx6SIjcGypJiROuBpcIbM8AvpqS0uE51cth8jdDs4gOyg5I04BTgBhFwp
d8Jm7dyK3FHcJqWdX1rOkkn20WTGL0TyQYkseCDtkYkbNBsyL401wyudNGR2w9R/ektPO9LShjhU
dPZPq5F5Vs2UzTJRo/4ofmlw4l0cvDCUmCQW0VCEz2DWb4Z/m0XmbtuWAa0HqFFAQzZ9tNR1wumW
8E5NeRx9caqspyOPeT5JHIiGliIsuk4zNl9ACnmnRdr/FyZopSLp8a9O4F+QJTk+g7dXSxrVWapd
0Edz2fnglw6YKufXJsG7abjt+ud6V7ijH40sNPJypO7FqDmgwEAU9uH0AbakWCn1H+u8SJAOsoTh
fRWrKbEGO9iHEEiH7AFAz9etGV+8uVERz/rk6brtfPcGBrL/Dtb7INEz8TaALssrRF12h3D2vwr0
z2ogHhV2AOqEINWoIvvhZmS6TeJaIICu+Uy1McblQEgBzGgg+/pxUukJznZPKOu8Ok0jkIX2zpTr
W2F7op4VrcjCT4JazBzrzIU5kMhRmZXpd7gQ1o60BSG7oO5ax0adK/DsPo2Fm9S3370b9BfNU2kA
67MYyTpxxSfYnmNPxgL+Igpl4e1F0NpbqS6P5Te7MPSJZ8njQVzBkQ6T9Xe4zJ+ITHF46tkpNOuB
qVjAmsRAQpU2T+ZcX/2aZKtGEnFNuCn/ihbL2PwL8Nbj6bYDrCdbm2pZnYN3h46UxUPZoi6Y7dU0
1XShsBQRW6BnmZmnZLAHDpZqy9J5jh/t0h9p0Fn4thbOGE1L2f26jEKG1OIIwt82B/fQMz+LhTQ+
4Do986M0eZs6meFPbbpJJOtxFNasm0KhlrvW4LiPwvrJN5NlQmqeSpx4gupIW+likDhNRb3lN+u6
mchUQlTmHRkKOQ94s4P1F3fDZLsiN335qRWWG5JbugJWZssruFFsRio3cDGSEkSJHeoSZ9aNe0Gt
G1ZcQc0ypdXc8CoN/6Mi94c8tvciAdU/Udaram/ydDECrJkkBDcBZMSAA2etTo6Bwk5K2gtW4BGX
k5w3lyWJMLIzpgVhxx/37bGRwTPLeLEs0IS1z+65c3BOV/l+A+LpNQWsJ/O33UYT9UDzBcWuNqyX
EQnkbrj/4aLF19625bLbOAojNzMJL3w6ByEjcqzZgAc8Br3wbkverS9GO/mavF4J9rahTshNnLRz
nJlq9SytladGO2sk8Tja0RvqA4CxrJ0dVmWr6ArUohQGRDy3XyOM7oTvvw3+KboCFaXvex89Ggdv
lwNP3MN0/aD5t3S9jKh7M+cXH/lytwCmzAchewpzPU/D8QkyRFStWNn/R+zhiJQlhITho09pmPVJ
2pzgr7LB7c7ujNC9YcAhl62Wpqvh6YH/jh/teeabOI2Ajc+bn4typ0ka8uPB7UdGwhNMNVbgxUk7
qv5hJ42E/ORu/6+YVXNISN9HJ1rY6bPWphDmcKj5T7JCZGgoq6iiEaP8uJQ+4/YJ7zlEM0ckSj/j
DxxSf2cumBMZcEJiwoIK02GU34BlN3mfIAEecn5i3yXolM5k2Vsl3PgUmkge9Akb5XdhD0CfAykA
af+yT7WDG67VO6nkRjCS0AIPP+FCcwIH9dMWl1mmU6tcrmAdoLLkA0vZJG3gcBcKZrLG/GuEaQIH
VFRhK7ZKxP8J5PAVMhUzl/hcoZ2b8tfV7bglF9BvRlVMckcl80ZfVz/Rs7HQjKrbU2R/q+Dk1y7j
AtjcPMLl1ftaQbN3OuVFeBB/raKbi+YjX//U8zyccgGkazzIr7c24eG2pTMkfjp19H3TCmPXAGNy
A7gA6oxadANhXrXBD7BQViWdF8uggx1Tn0IseYApnV9tndzpWsL6a0tBG8rDcjkdY5pp13EAn/0h
teZRWYry08aUtbKqhH86GMyWvnCsWF6eIlZ532DX17iEeorsol34A4XToB/PRBys7Kz0x2uXTdfb
1CT37302OduufkkkFFv4GsAHZ9IAGEGWevtR8REwaNYg/0suD4hBN17MlOUf3rjSwx7jKcSyzGAU
PKdrxvWM7bQ9D6pzI8DBFItXEIjEmG41kYDyXcgRySK1FwHS7fSNZCG5mc11D5yAtFdWylDDl4fL
zu4mUFp0YEZvnZc2pgfSvvx3dJeBuC+mhTqjkgA83l/1PeP0OeEP2buS7zYd7qVV2x2uorZZt+H8
3IFYfHPmsQ3kbJGXr8cLOxHAlCdRRp6F/Lud2wMBUVYuBbLZfxhVjp4jvHSY3z4sxl7tdbwsnioz
0sCqstzK33BjW12DqvXzSIlrCaBkshxMWMrJjMrvhDgDDxDa4pdvGHDGAgqDuA2RqXt6tn69iyPh
vRyn8hVOXGtKUjKc5G+9DbPHos8W/E11OkYs/etSVRrZ1+bFJGJ/t3QItTlbx0RKcgxVcb9CxPy+
ROiCvvqlEUyeVyqIfoHCnkyjUL53BjMwHpfSrlDtJhfIGBhEQE9CkiMofFNncKEsbZlULnt9tdTj
vbgBCr/JWsHdjRY66Gqj2rFKKs5EdJjru65v+jWwgPRNSpwDt03ATOc4djgZmXRqWTO7nH1V/nJ4
NxFJVLKJiEU/ITpdIUO0rgbw30M5Fpz4CGLvvmnk0wdpkHG4OnHyJmGhY5BwOtR6wzEDkTfx/EyB
kO2h03BYGNXJ5OpVwWvcwT+YrtLUm/9xuFXCSx9o/QMsU7ZobDg+FFqxInE+TmwkaVum0rnpCMAa
ZxJgLe4r9bIawmnyJqbJs230Wy//6UR+zamotzyjffhvIttxQltUCuTsJhnEq3JPZmngsdeXrHLg
ZdFEX5chZfN2ojqkeJyP3/tJ8gZwyLuZMPTbbkX6vwwIZUObFiFsMMg1bJvVYioUg8VjAnWcZJq/
ZvuIRYdT8m4J3Xxp8e3uNccopQzjOnuUKxmgOCd/rS/cWYMoiOv26Q+vGm/WizNh+qZG87jeoql3
z8BK25CqtL0ohuexSGoQ01dFMOyaFgIYXga3Jqu9jBA11z9tSDCLn/AoIpYgqakH2cq6ACESIKUC
fKuMv0GWFAP8+rqpIKEKu3ENCuV/polO+Hwu6I3Jt1VWWYnj05fwio3EwCf4vcOC12tFvB5R1wlQ
aXOSns+HaRqJyH61m+o7RxKxfCPeQ2o9xhx3Wyk5PTHjah0s0Op2dmOh5OpxIsMY4RPiY89/IxZW
lbNX6pcCXP6khT6ZWMJK1VizRHCkL5o98rGF0HwGgvDVrNG5iVQJXI3+049upTps3CGwZH+uCKWZ
jSlDXUlgkY1xeJ2bW98mftncDk7DcQNca39GPFt2qNAaJLo9WQSMoFTPByi85pQv1f9kpI4rV3iN
in0r7WKTEqvaWrxZB8fKd10IHUEctE/iojte+F75nFAVd43W0aU9EghT0vvtckK+gFL94ggvM8io
AV9bZUXqUjNvpa5w+HXZ27iKLZ5C5KlFMEdgLg88pJ3nHI+6vQ9TjP0EcHMV70KMDEM1lYdcu2ya
iNG1zojcgLeztn3v4CGe94xkXzwHuoiB07oS4WjSt+2wZav5IppuN9IUROavCGKwmSbr5vEPvr2S
9v7P3aMD9DB7yJPclecstH5FqVYmqmA2Ep9m+w2hcpyGMTrWTeibMNgihLbTzmAy7JyqaYxQL4Zs
Z7odOEY7teT3guCZeU5r26MRfsAPx+3NiUpe3o+/6Hhiz165U9OdNdY5ELPSJqSUxll2MlhfxwAr
8dwVqJaglD2QaugfJiH9YhCKKw4TZ1Iur/erkDv99/S6JnywAZlTnWikOfEW0iFVvNIm7SPAxpHK
1Td7KBK35EDApVyuiYW9XLHfNyJ7GriWkVWXQOJ31izl+I0wR12vtle5NDh21ihBVGmDWdhN3J3X
k6QqxNaKsZWRxINkHoojWa1EWwyyYmDygA6i8KQFLFX2haD17XHia0EGmIs3colgF6UXp25kAGm1
hDizpUk8vu9WpboMi622PQbEmHV6Aknw5BfaIdSQehiCeDEbSxA++4HMBnEFcfOgT4D6LRtZ+Biz
QMU5GWv5zcXHDQhIfwFIUxE1HajZKdGf/L9MNX8d0+cbfURf4+D9aM4DeSUuyS4tbA+aPoHmcdoB
qHjoDExAmJjMKbtqe4YxkVDiTvdtn/eSjlSz6S2obNAlmGbUk9xIGkXtdIBwtgrVlmKpkZfgs0zl
5Qeuul0X4UtTGPfJxa60i4l2HUBAa8NUOvWvtFwYR6Ljz/fmbE+hX5BiGnccuf6/ikOeALzQMZRC
OwuZ4NExG7txV/23QY8t9Msa+Q9RB6Nh+pkrQwziZy+bOZiJ4m70EWFk3kEYaCL7btLPa839mKrp
Y3BeZjdvPSHiAQ5zDA9TB2UBjfo4lRSajdUVVbmDrPFdvz79X3yqs7q9ewksmKzGVEi6Fp+6vtBe
V6yLW9wx3NoynjFAgO8aYajkjFn0EdXjg14b60LeFe79CLXTxJadlhLj5EjuHrnSndJYhCObhk1F
PFAsKfKphVBSRBZJC1aBm/BG8OIEWOkjAyKRVTmkcS/r85UlGjs1F/lP9Skgsl2oXJap4ko2rNGz
6BZbHnKu82psK6vAQogIDzuGAGYpvXY5Et62EaayUjor1XYUo+ffzEx8tXZXVde9UY6cXcQKe8YC
Pw+9/sJMCgI8B3OcmZzSGIAw4Jvtf/wAaJZPblBurt1rpN1VaWxFgsrgHjc4Vgcka9KA0ThxQYB4
cikWSQ4j6eWyurTzFVa4glQe1TH82duwFOlbwNhOoKigKdvfCWVTpjAG1rg7IDc5GYTLqtfb9enq
UDGXiCZTWrp28Spu/3v74yTBQpE06AlVJa9HxFY53rlnGucS4bwREOHmgQ+THPKX3TJaeAybH3xa
JTBMKZZyZOXTt0AjDjSsswkRDJpvYD3KAZasIbX3SzoVacADaO5BIlfZQ8ehND42NOZj7xd4+nXd
bfx850hcojNA0wZUNGnEeMwwxYhGiZOUR5gEuuZH1gNiD2ELae/2ZQYdkAIeLRZ9k6WLScKBt6ci
Io9GRsIvXx9lZenbkD8lEpn2Gz/yfiAM73ZejzTsfnv1StT4q1TlXWfbEGnCi8CQgHno0mwoxgj9
a/d0vwcd0aYqIfwpxVkYgQGyJC7kJF8Zchy+NRjVs2T5TLo02bvOgcnCqIiLNCk37S9Qrh666xwJ
hFBCUirwL3DS2ZD5Emhr3LRZVtpCUfvryPPVljGFFlC8Dfxnso4lg1r3VxDp7EN+xiXYXcbr8RFL
7t2QABvczxr0AVR+726roP3mtv8XhIJUAnLqHrJx0ENDBFFkrde4BIWUdy+hheNo6/ea5RXKBUYb
/ycAtZZ44lzde8gFqYYSUeer6mpcjrPRdhMVw0woiwBzLk31MPOF7Eir8GUrVT6XfH+xNWY2D8xa
VvzCZkSrZD5zlszVotTb4ItFIob9ANV9yjTsDgDi5bKYvStYBkENFSHi+hF0N6tFqKcyYV33qQrh
lgtvvMArfxPX9FadKfL7fdVrEOMASIQ/OfJ6TlO8YIRL+QUac48K1ksp3fSIGHKvbHppoFMP3A+A
NCCIOF9SuxRV1mdJVWWU8lc3M7AAxWWqhai4Z2z+xxvMSD52geQbP5dyIJiiXixkiCW87M2vgkqQ
cLiM+N492diVDDRs0sjvEKek6AX30aANE2PGH9TH8wmxvaddIfm+YNTJnmwWiQ+NYFih9nrTzVaX
eACC+H77+s4E+db/9/sB01VIyXpJjBOmId8BmNthQd1m2BpTDAL1i5I7vEy+tfxY5wsDgm9jVBIS
p57pndQ5QCP4sFsR/pJCO4/eF/k5ifyTVTJnaLW34BipNhh2adjgBKMU8J9Yugr+6TZc792Zse7N
ui0Si7Scifvh+FWLNsFYP6Sc1PV93PkHvu8OiOzh5kd0nxlsQJiHepZPgNyLS4SE4RmP7N5709Cm
jRR/iJI5yHB/hoGydnrf+tyn3E3wixA+NIewHnKPAqCcwkhXM3iRlIIZnUAoQRmrtpNz84RRpSR7
ByBHugE2vSMRKaeY/GAV/lwEFDDro1RRF+JTjkx5PNECNwth4pgHwBAtR34hyDa0uN+CvU2gMyC9
YqS8QYgEzhx7yRGnALtOOVOEomAxNiDW3gp0Ru3mzcO20QUMZVVhBrRz11OAlSPQBUSkGZfQiVBE
6ta/8Hki8zRGWgHeChtYOGgv/gJchlCT+xi2deko7MQh5BflPIwUadDacaZ8FqScrgjIXHeG2d6f
DbJjT0+5zEbM8yUtkI3u4PUaHuyKp46eSq3Nh0/pars4mRLOMJTzpIk6zPDgOt2oY0NQpjllY3u7
VBGgfe4evPhETtmAzgIosk/4f1RsJ9dCKuBTUw/Asd5dSX4Qy2lv+fgUa57+Y1XqVip7xajvP+iI
HPp3a9GlSmKzUnNRbDIt9D+r3f4MiO7DIpPy5OOPlsuge1YPYbZBsjSJYwj4HslV9K3y87/9rGKx
prB7saoBwWwrFeEn1yy4HpeQWvuiCiWkCPFN7d8L3rYqk5tIbcr2ZBmeHIna801RW5S1sv6GHgrg
fG2KtSaK27j/81o9tCkJn3HohO46zPybJajw7RJn1lZHSr0x2kN1JrPvGQMdB1Dl8JltqnOwJNGk
Z7FLqgk4Z+xi7+eveyQz86bybs6MJbJZ+UKQP2Xpl5qTgNbwWxAtKQNnzU54P+4wB1JgO9z+FmjY
KU2U05/zcrfO9iaTGLk5c5Jx3STTUWlzZaFPB/Ej0IVxH4+Nu62JgKAiEosa0+rOXjRvCnbpJybs
24sgm319WrqKl23bdpUGahB17w9i4aKZ4BuT/NHwBerS1ZVDENiXZQXcIB2SZNpTTz7Ha3Xdwldb
iOICPXX8puOokati216QgO073avpznpSiU1fmfBteTWqkOVsLQ2sg6066Chfp1PbplpWPMp8YaeO
2+ZunzTPjI0IlLlHXfyMs7HTv7hnKwTUMqt7X4Cr1QzFEY6+0UvUKeciNXTst7n8opZuW+GZ6QNv
Lw12DYCt5LbzUaeMpi5jB8jr3GVPQ5QTlA4OHGbpoFuPbnLc3U2zNyEH/ymU3OJRvbHIjfDIjlzk
ukvCn2We1MX2Fm9+TtzhqiP1/TJRxCFmxexATIgYOVMTUs2gYyDVGxjrC4CPU8BUpxjGwEkkgQoZ
AsPxokmvqT/I9FeffW8XSfwCekT1E6zd4w9j11uxm+3Wak/aVlnEcNSWyK0Af3U/93Buc8C4xENV
z3wOXLWqwhqocwLAQU12rnHte56TRE083m9TTh/r/Kw9UNgr7AcOzqCF2omfGHhjddeATN68tLdk
9pml6DO9pPfqmjPsG9nqci0gI8FV5z6kGWIaVtx5c5mPc0l1GD/3dIvgDsGu2wP9nBunQJPd8TAI
ys04Zl/lrOU00fWWVBrMgucMFw2UYn3R2G8IStT45yAVNovhHjUSxX8WHfZwe0qRTbzxJ5vhGt3G
dpqRCsTjeUJrhhfuCT88jnR6JKY7cFbHikfMlW3NoN4fzF0EjP7vGFjqIUFyInVZ7zOeltaf33jY
xWUwMUkkK1sJaV0QNg2+Sl/J/rZMPbMpYLkF1aLo1DtpXAziA7fsRJx66XdGUXW3+zM50XM7g8a6
H9OQaUXwYSTGg93h08h++eWXL9+SYn1MzgqgKLbit25q1TrFv8T0UvEwC7EFp57nSe37ebauv1SX
IM3kQqrvRxoT9jiIic6vQ5w/D+7YM0ydqjKiPzExq2JSp9G33Z77H9khkzTU43L9QJGYd4/2dWRF
PY9UDFzhuSytReyJjtVMy98xPRrq1N8VYg3vvQOJNEWherexxbv0g5hahe01EBjUwpxFTjXzLk3O
4DlWAXw3Dce4zrva+/plrdrBp7/4LDmXGPDzd3Y6VqhbomxACLyBEwjxPlwUGFqUCfH05YRhK4V6
DtzD2RQKZQy2KUbCBcmTwJG59hbExka4IffRTQB91SkBbgIge2rLCgrTG94P1Ev8cb8kpUkoQlb1
KRmbMyz+g5VRXICh2Amv16n9jA9DsGdChvlNcBKBfd6zn3B7KoiLaEUWbiqNgfZ/VZw5eKkjgDtQ
N3cDhKFEAHarqbPHJpQ2QEJK3O2mJgyA3RHrBsYUzCSoUY4sa9RhKMDUPDYHKLYt6XA29jeCnOB6
XGWcG3ikl5qwfeJy3FzSPpzlIFT4Qc4NbQjy9RZlYGKDFww/09Exw8O+QC+Zyzb2JVSO8jLY2c4a
ZKxKwqo5rNga8AYxkX8byebJRdE7vMpXD3iOKtD732V6qdFgAjeaAzk1kyyMPA2SE4qawzPb3jB3
RSX8TLDQFyKuRFFo7i9eeaWta6Iyc9nydvodELUG1RKCWSr9H17Su5Y+5claRh827m79kin7fwAk
mQyNEl9H9bZBm8ZrKF+qgEWCTNyI2Okkcraf5aX/+LEnH/IteTGbKTLTU+N75ks4CQ0nrq1bGVhb
c4VuPOLyAl7J+/GXaBFUafB+tiGh1z+DOzD7BmoYidopNW+VuIbTLoo7WTiXrToDlY05/l+2D0oO
PgcY/Lfu8mqVsX5kpoRZyau8IrehJTvFFepZbR52zbraeNmpMcyt/wOewXKex+TQwB2CLejjSXDq
GxTx+CPucJ4pQGwqhgkB7BJi33cAOyYzq18GkEpQONCmN592h7JSiBnpIEh1GSzuf7KJat82xwA4
fx16VLBpPJmILGRaiCJ2muZD8msDteiWyrZIjeG3BRWoVka0S1GOEUZCrvMSV9MkQGz5e7KDUzyb
GiPSIsaUPr8qxhzQkpg3waKv95f6nqM44TYK8tIgKnSigXYrFPoRxSY+23vhIvWiWCZd/jaqbnIR
KMailLSUqp956b1PDmsMZ+85Z2qDu+E/udbJsjFvebzflicY9kNUzvpsapX8KwKrKIRghtlKvEBR
8SWBEyafTUzXtVx6fw9GsuZUMz+42W8GoqqhzDLogYON5n/KcZ0AHr3dS7xIEBZPlMDB6M56Qs2N
UXCr7vtHV1EYwAe6WoaIgxvBTxE0UcNfnTzvYTQqGf6BRBzUygoLfiEQ5ugrJap81uyei53iXtFK
Qr6vl8guzWPw/SS8Q+HLdfmvqpkbKMKHOqi+hkC97JBANl1eyTljOFFDYhlxQ+//eEgq4Lxzi/Il
akulCGwsFJn5M8aAvkPrgxcMjfCTLqaGZT+p/CFdBwe8AYusH2tTiI9v8Qf22zpuw5xRfM4RRNs2
Pc5rQHVwcdAdShGKbfgp+R0Ev3s1JwHkV5JCce6N0fbSR7HmJ4Mf//2XmIDxIQqWeMbyaxyEJh9V
F23zoMoU9PyQJogBeUVZtEMfSMePsYTaZ+7KFnaTeUmKlxBlAHyboN3W+xYw7dV7us7fASdFfNhd
YdYuwKb5hJkIqby45cnYEBYgNz9tzPC/hUjCD1zueuJaQkIpmtMHuQXuHYhCFRzq64Cjbhkw6SKo
OUyGUQ+P7Rm7Xq1PLjBe5nkOR9OKObO64tdfwoR/nNJEVLP9qC2AV5edo9j4pphyAzwZxmomv9Kp
U/u/OWKC+LQ4u0BBd+ptpBnsjcpiGUfo16XrRYhV3yg6aLEWa5ZQ0jG6jEjEBCLs2Lyh8MRsU4Wd
JcHjJBjTJygkhfkzSinctVgstqB8XwiXliq/WxIs/10QZgHxaGyHUgaB3tTlTycqinZ+EFd8A+dK
GOCBKEMy7Lfi3yP/45FIWjZNdWdQoem1BGLMD3WJG1kec+slZaXTHesyIJQGM3OO8xv+aBmIx3mq
fNPm8VJknVrLdTP2gvlFuk30bG8HXzDawUuH+beUy0NCSr6zqbtMFmvu6Q3LxTlLLL06NxCCNP/F
uAA4SIERKGovUVpNgny3aLTyoJiovx+hyCyZB0EN5r8YDUYdaaBPgaa2tPayepz9ZaceihFyPBLC
vx4htpEaAa4p2KtVOA1TkdAmKM/ncMfYPTlPD3PyX7Mlum58PPrMg2hI4hASkWBiNXQ76Qtikk30
zVxfGu32YE+5AJZ3oJPxvyDVQ08qX6cB1JPBDxanRze+70wY/FICRqK0CCMkiQauUDUtlbSLJ6OY
FaT6RHevEgjpwQqBOIVABQDi2Pmq2Gstyyv+550kOTbE+JgJ6krWyUIyxh8QtqWFrqJR039BJgpZ
GBrgS7FmuHB3AS60nO4bVcPHnDaa+/ZpEJlVQSxTlAlf1n8E2itRQyVd8WSsLsDGrReotLqlUO/X
Dl+e+TuIxDQ8ZMVdbjy2R2Xfjz2skOxDhl4dlqvrt3mtOBYYs9+fEuj3VQvYMRgmumIi0KC0osPc
/9fbNOuuo71vDv0pLcTNSiFBaXNkNAsZmRDI7h/0zXvxp5Sy6Unjc3d/Qi6TChwj0SrHoCOezuYu
iMntmYiHpKtBADfs0zMtRFGfA4JaoaBhFdOARBowAreQpXOKFPlFlJxIBAiy2au4rn/HTGG8NEam
WPcXmQsveuujYmqImGjrMzv4vCHkDNpIgI732ETHvJxQswhrOOMDlHXTfErOqNEXKXPEH0kGjQ/u
jDPhiGwb0HIiB51OZQkYg9phGkXjWCC37kSZ+j4hB8HneSlWwaX/80qrFIpMRZVXKALXjZ3b2wqD
YSxMTUuIqU9yasSqG6z37q+WSeg6Eerfy+VwBydJV8fKJAkkPfz5qwBBLGYCm55pb6pxvm81COyP
gCB2Q+smogeWpg+vhAfPlPs7KdBtlGZS1JUWq83+9HfN9g39ShVr7aDHGaUoM8NIL70bUBzq4rQh
yaDLLm7CFQBT1/7VWPCLQNXwDxgvdaKzuR/Qi8OMukm0adfh3J4cyEzonL1b2NEQnxu4Wv2PYPna
VG4BnbwfcblVOFjqOtY75jYsqfITROxAzVQGn/AFUrEy1R72ocAfZWrTwNB/OxgtaaamB22qcMkP
5bnmi4qcCzse/2Mqh/V+cTVVEdjzXYtZVzl2gNtAU7pDJZee7zyJ7lRNDSyGRWp+lm9/KQYcG+IO
jEh8yTZOGrCdQjAXqYjxRkgFidLT3ZBb2Bxp2/7owTC1jP2nG/b42ZR1ZXJ0dBx5fSVUI4E4rnL8
JntMdTDeHeIYwVS5LobdnykTElEEkTIocuP+Ucg/asRevPgBDUEY2bORr1NJ9aI1X3xDdUAR1CPy
IUkTu6nReVKTqgoCwbYZDr1HX56wyxd53QHSL/Hr8SXp06mZG2ZZXQMdCXVk9TrdRKsknlodlE81
+T3ThA0zoc34CFd0szGwybF+kG4L8Xv2N6mPqVeEKkegT0KornnkwsrAnoxK8DZES8nyQMg9Ucxr
h3TIojSG2vssrgo7G0AH5F0wniANj8aQqa4e7TSXUe6xnXWYp/EHAXi3o/Y7LefAAMhgUCF7FbtX
464SW48mxxPBO5ZIOKnBwRBy3y3osUT7xWeRcJbVgkxS2v0DFg2ZvtCdxmXwYldH86/B++fUnjbG
CGX67Zs2j9WgrUJjsp6jUHrWeGb2s1fnibbfWTDKGA5ZQRnGk9n4z5ikTjX9Mx89DcogC5S6oNDV
0l7pBU4D5P6i2FQOqwMI/Ug1XOKP/2Hm3wE8VbJNh7dJ8QiSrb9o6jev59qHFPf/B4yZDMxKueIQ
xXbBK/6m538Kurlk3bvTORSp0yGkKNJC5jaj4Mt48V6PlBuUlj8+IRKOfONti80m0rKX5YHOvnAY
X5h6vov0p8B9e/D37/NAE1q53FwuoolAXJrkwzZuG0j9gvCUYvX8FHmAzMlBYQ71lrYErnCPgUJR
r2aQ08rAphWH/9Sptl4kRI0UbcuQx9IU5YMgPf+le4O8df+zmXRlj1utIpaWg4xlo2HAqxvXLG7q
h5Y5k0ZMohbJ0LlCABkd7o1Agjmh3P0kHfNbfHPhBQnkg7zVR7zpkpOeT3xtUW24zZVM2HIBIfLi
KDnlYOTfCd+HLwFVwiivtJyiCaR7RLNMiicAd+K88bp5CNSReL2ZA23Un4j/tWqHuEvzfQEV3oDt
iv3xNcy4j/54EmAqqC7knhHv7aQnBwY5c+CsL8WJnb750B/Ma1ZLQ5wVauMQGgAK4e8gpKGtYa00
JkmzcJrNQ9RV9mey+x2tlrsIAMNH2gHfPfYada0PH7sOAUXsTCyz6/GU+4vy1i0P31y+jfDrU9oG
+Uy5J9BYpsKnORaxxfYMh0F9iM0qKg2UpA24ZcUwJHGADgsLV+OjChyp7APmVyEOZPTDYiVDNJYY
+0YAcWW6l5WyRj7a856UZ8HvK+0rMOsqKshcFGj+xWxlQgewoM0OwH6urjOFELJoXvtuEBV4xZrn
O76V3C6FImFs6sfYnBUIBVWsymB7GqLBJNN/ctDOh+KvAhVNAtieI8Omyp5PkRAea1Hz4whPock5
k0CsR5wKUDMCzIfItFTOgnCWGyBVemA7Ds3TVhrQ6Zrg0KmSekB9PUlmRJxx7jJG28Bz2dgyQEfp
ShY62IsAnwuldNvhbV8ZjMB635f+sbdC4/pJscIvqhiWmvpDGde5KEvtW+gqa+/sO6lRSsum7EY1
VWV8zYn4QQM/VWLufdhDq76u5Ap4vuyhzT8z4u67gxN/HEoCOSuhTUPY7y5jGQvDvScyQ7k1CXOB
qTPGBd95aE7tGwCppnMdg2itVlDK7pM9r39qH3eP3N3kFeerR+Mr5atJDU8peGIK/KaAPaK+jMo4
sSBZnQzFiCyNyM+A7oUhAV7wCz/zgs9Sm49khWC16kbS92Zd70SRB4GD0FAq8aaR1kPkY43apABp
1iJMV6ahQjJAVeAk7QzwefrcSWtP0pR3cS0cGut/GK9VHZgJtZfqyaM3J3XFG6k3CEipwpMAIqi+
59KZkwONgP/UpMpngqfMkJnSYFG+T+K6kYtWV4fpwGTWey63coX7CUcTBoD5cvfSSFn7xv7DqhJb
v8DBAPyULYYIQ0Dt2iqiEL7X7lsdiwi96U1GfG4m3dGJuLPrBonUV4Ng0LKnFGmdfi13rpRyQ2/G
/+DE3vH9uA941UCXuWhM3tlG9BVCTUVWrbxTqWgBrvmkiPBsgbdrq5IbiztIOldJKn7GYU0KoQNV
U59JHmadk7vOYZF1Asma3Lfkxc/0Vp9b1+r0li3//OwOibgCUrvrDiQ+zGPYd1UXXYPCEGywPlOX
Os3vlJ6V/ERixfTgB2Z1AhKnpuwHrdC92OEiCChhnC09H054D/ePBYHRVrhjv1ldx3d+T69CVGHA
tNL/Hg8T8Qu5kLe6z4bQ2+lISEUt1qQydOC+GGQhR+aXIz4/Fb6EykKVmVIESgNLJkHNCQddCzeY
BNlcHKvXPBCQT1sIN/1TgJuoxfJqx40NugieSrsE0ydzfM+aGLu4x2hhpWqAyXinw6fMotrR4wDq
ccHKifHEK5T2hgPWWQ++jM4V1tNXQNPcmGy3oj/JbXHybaVPcJEs1Y0GM7l/zufuMWUkwRhmXdco
8QAjQ5bMtO6bu2Kayla5br2HsfC23DJa3tF99atHdAWlfh4p1gsqoddbWZwLqY/i36gL/1tn6E55
egUAATie9xb4Sphs3M/B6R4YezZoOWLN2ZZWnP1Dk/i8crezdeFJALe4EBWwtm//xeHiVVjPnAij
fPQfHbHhlVwdw74dv/wczROtM8PtL0DZxa9ryy/SO8dn8vUuxZGNROPds8A2Zb83EklPnap/xnQj
zLyY3Zx3Gno7LFrdNXDZ0pXSRARX2el3q44+4iYqpqp8iPjtWf3eeo8hrEJkzS8DAUzwY6QVKQQ3
9DiVXc+6yy58bJFXrIahO02svGdn5Onl/j7Tt/a1yiiHcmBkWdsOCzy0gXqK/sTEG1t0WZ5kqS/L
LrjvgW+BO0OwvMTR3UU9w91ylsUhMmvvpNybWXILuPlUDEZXAHz6/kycnYltN2Ue3NIvKUMimznW
D8gsffcAaQSclgsPY3hFx2FRtNj7u/t9/PAttDKX0OwvHIYDuG4HtBbPlw04CmseFfMd1UeIPT1s
ANmg+yDFy7uQhhv0dDHSOiUIge5bOONdMlOWXnnTuFfeTIeAWUmmHcm/7nWuDHKv8s8+zMfKnjDv
qKbGdS38o2hulON/NW7Ju3aq0TR0A2PWVHQzNCdCB/xjuK56eSN4EOfjiaKiAyYAfzOH7vHrIBoJ
hxmthJ3o+pFh5Is9jImMHulOBIcgHidoMdIw/ZHuiWI8zALIISKcc8Nc20Dlb0heCgByTwF80En0
j6ogA/rtuO2lfbzGEjlCGphoyxmYquOII62k88v256DGTwU/ELTe3Bhs7YliDgoKBiw3d65Ijasa
evi1fVyshPxUlRfTyEf1oYDUZ4GrQKg67CGpTwog7zigqxLc6e6Ml9PMBxv7VB+LqiT6U8aC/sbP
aSjNYxMlhml8ThXk4r73V0tFlTwREpHKLzB1H5UJlhIBSMrk1sGzFVJTze7vz90TMz3iM+P/QAg4
H6/HU7QewzHGFi/zzEidnUIkzPwp/ZAfV5rCYEe0QW05a9ij4sMdZwmuS0IiormfJINp89m9zmBV
ujDlux81IquU5wVVZJGDNqmW8qype681b13g24GX3yR3ZOt8RSqWbJywPGKJkWh1iCqZWc5pi44l
eE/UpVSlaWkNiiqvFlyoamdytWsJOMnlBKFiY0a6+Z6/0uXdA5uWLxjuRBejMM85LS7WLr8Pf+5E
SyjAg4NHWOLCWYWo2AdS6387HRdKXswYQlUTHlicCxokJr2loxTsSf6E0HzRK6eSnI4aDgRUkxxw
BjFU77fzsaTjqur3cPaO+QVcWo9LVxSRpJFkd0uCi6VMiyzxZBtdcyKIpwozbTtT0ECarnp0JYKU
DcaCBHWnQOQm8QPQQGoGkwnAIunj2f9kBUdp+lqNHOiIqRsMGUNAH2POEOes/Mj2wO0aOkaI0Ka0
wSy/ooSaO6xTdz/qFYEoXCINvBi0enkbXQ3U5g+pYlA+kTvzcw2OPbWdGZmdQWBYdA8ToZQKY686
yW3+4Ivn5cyVsM19MY5ZkuqGUYvi8grPRwdOwLqfsEOUil4LVZvz2xJBYDptl7us0orlIEzaW8BS
wtjR3GpMbQAzyV1YyobSkscbbUvvm2C3GgZvDNcNme6dvKro0b+I7y2lFLkNXzjFu6tGJA7FBL32
2N9wsHBYrWSMeOXci7pjQlAWFPhT5QHrr3s1spUmDNiFr14zPLClBYPaPVesne924e6JABzcqEuS
ZdJa6r/4Dmm6pT8jlZ1VRyDkMMYkhshej9OUfnfo+5Htw/8GCUMmaWRifeZcIt7rIeifOfQlK0bf
ue8iCbr93meEB+BNMjyXRRwwjhrQm3HoeDWPhV7i7RLkMWuU2d3unPXYWiJeKzlsjlpb5JsIY+VM
XfQRo0BIA2RBaPcr+Dg+C3HQS3zmf0IbHFK4g9he9QbSjiHHuVpNBywvSS2liccGFnQlpwT2p+Sa
BnrHaK5TskMddRh0Btz/iiVrVJa8Rs3HW5IOFFAjN4mTkahfDj/NBQt/2DoZ4k4Sqe+0HL1YJB8s
b1qKkorBxOg/ldKX34/J9ShNcAb/oR1NJdMLQ5qTDBGQJ+BKK+Wa400H4QRq/BKI2+H4WjAGIBDC
V3EIR/BTzjLAuLuX1WPykow4wzt6GqDezHBEIUaQSoqHlcmlV02OeQNfsua6JbUvIslbtvBEfPt4
fMkiDsON9iNbDc4qNgQi4+WS7izCqFAqQ+C1eEH8mrjQ2cFC0f4GuCgB19LrH+FoJZlZE9NqhTn5
WgCnyDlcwnVInkjFG8PlkDbzVWzMBX38inKt1PvdT0xPoLvfOBK1Aak3q50jHS5A3RBd8Y/0FD7l
brBS2rBZ/xEujfMKBVxYC8LYoAaB9ZEVqPPqzYa6z/UH4nBjU0D+7WwBImMtPVJESjGImuu0d2C5
7BJovswtRgDWZ5mm7Mlk+B8xXTZDlhE9iehp97UXvooiQdyAO8GToFLiiBdcO3v4boYMhHpubIxL
5U8TKDJv2duZVzQGaLOHxiG3ZfI5W/oX5yii6QxNoU0K5sVGjgB26H1+N5o1t39rctWNGQMxTaB/
6v2aI2+/br2gTtvEu/FDwXMyJCOzZp8nAyjNMlCD14eyh/Rg/jopKFPBEIldMTySWQyArzLhfShP
4I2791XD4lRvW98A+/W6LLSS+SCedWtTeDK9sOhsimSPla6dY4d5DwX/Qbapn1pKN3e9UiRZdqq6
CUCebpBFsBuj08GMj358v8ksn8/tE6HWXY+clT4EHZDdgKUmB1+8PvFeL5JkUxfCW7xa/KVII8sC
y/5mywsihMxUaDuq/CmBJPU9Hzvil+HrNMVE8Y6eb4O/f4iz3E0619Zs06f9v2ZVxkwILCV3hBa3
IQDiFZDlbFyDKWaIXsXxEanZ9L30RzcJdWwIRkEtCNRgMyuMQCA41YalgAVFWDrjT9WKkNf6XfWi
mnbMrTGmQMyDpeR06GetkIozGCxHnZ3cG5/uRJQIvtrIgoW0usvhsYkgCyDkVfE1wkSguYx+ST8T
A2FZzS0o2NyO3sF2PRlt2+hpJ8RK0OjZwoFO8tBM5l4E9RqjMBefBY5qJLP4wil938Qlbq0NVk3q
I9S7kkoPs/eFwVeUzZpqLhNZSWDkfR2wHqr+V/o7r3Crhe1SiYbNZO+/hKBpkWM733MLcIlbGTwz
yrknu8cNqDh0ZXpUz7QrnrbScA+RjuXvx0d98L4nzaWjDD8hyiLzdWdselPJdvLMZlIVDr+k/xh4
iXSCn8DvkqcqCltN2FTaFutvjjWYvHTuf5D+ZTwBHJAIeFzs/u2fa7f/1R1fprUlXtVicQkdmwhS
I8YVgag0tzHQz6k6iA44nhBXKNeY7aHzaidoMOypwKi7qMFDNXg4kI9tMFsAHEtTArRFylboJClE
kQn4yUGLUcrVmY5LfCdrteal3ry2YYYU/qnhhybEkkqHYDu3pk7s1rBcSVkaPGj9tbXcuhpvSgaF
yg5zlEHOUgJjaOfndAK5o6tMrzsnLURFUCL86S0imxE2UD5VUG8hJhXyuk3ZOPEd7pdAbGBWA4kT
PrXYrm8jpHIoZgXI+RMIRfN9SH+ahzeRWAlFlE1BAIwFEZHoJPU6qTOe+t06lEfEbok7ntjYD+L+
5eki+prgLqy7nASRP6qwlg0W9r/o0oplXelzg8y8WjxL1800arkMoTRUXpTaSbYhhyC0Ix7QaqKi
iX9N1Zd94E3/3SVBqO9xeXVV+0h+gZm3XK7jPdrJNN8metA9BM0Z03q7L9q6qfUpJBMZT9TwXF+a
TeCaYhTsGpi1sOa6+k6ro+vPbhGHKpPFr+ZAPfyzD4gU+r/6zb7+TG4sSzyJtYYgnbGrBGl33opO
4DUPsgejiRd93LxFMS4CeDI1Fs69sTfGkg7xEGKOi/zb1BhPSgZKxnqSImgcNPl+O8RDysfU1T3h
7JxVyb8CWDniyLq/gcOWGs12X5JeevCwY0r0MmIwuEKYvUD5KezLhw/9urTKVDhhg9SSpfJWyZNK
lwGZq34v1RaXRFwRCPfWS1Z611XswSh7hOW7No9HrJtVDzYPprhjiD1UTgOxwxIx9zQitnAJrGZt
SkdiKT7wfZxJHrrZSnVqK/h9XSIvJ0azFzzG6RRb+HFauM3JUVZEMIsKSQu5UNt4tziWdcBg32LQ
cqsgReXuySFwHxWJrdp6Kna0WmJhkaiPqW3Apc+SguqHroRC5UIOA5ccCEVtC1r2dzlvrPFJl9fe
TEzkxKZ9zJf4v58IyffUNK37tTQn9oAqusu1rtJfY1pByor5IGNTUXST7aP/8N+F8qJS8+r0/WS/
ZYcKplo+mRbQBsEkKCoLhy9eVAfZxR1It1hCQPwM73r5Gtm6je9Vit5OB75OPoXaU1BF1TcMEBEn
AoNqOs1jcZ9GG0kwzYhNL5Xv5+TiW2oBANBrmjGGvciUlJd1LOBf/6R+X5uzekoxLgwyLAWpGwBY
XBM5TvCnVSn7fm6NA8i5+mEKpc2LC6tdbsfctvSXjb5IAthGUxeF5ylFAAw0SRheek8vNhVr6Vfu
eD7NvkGUZLggKYs+P67HBNLPZH4B1bM41rm+ydTEGYG4vaqDdLge89MHEFiYMaOFYHiBsky5T/mF
Yp7dWz9D5n5Tywjq4ODDSmH/codCWFnXEvS+CfyLY55Z4Q2tCxBdTRIydAn7GL/xcd+AXpIGFFDV
Ih/jL9FLM90R4wMyrORYTF8uqNHT4kjjNcUmZ6daJUyKadxKRtuhc/WTRLAWjhWl1VHe6u65Cmzk
4XJLD/tOi3h3Y1eMs5iMCHvaERrc5P4/bJiuJgYH78lx6WX08Nxr46VQZlmE6t2yPbX56uSbuEKu
YlsMT3WbQRgJ9+373kgvWxguI2ND5By3FbnmCZLXF0XgJU2dOqtc1Sfpk3oZwFc6OKfRIuKDMhTA
T2XEypQ9vFRG4ucAADGh7qPRS/YjLUqk70sCt5DbUfptF/+sCmWFnoYhdK5reRszDmluAgANHT+6
HiJkpsCdOHiVOEEoLfQo4stEZX5OVPsKkpFPjF7Jca7+fSpnrun8PqcRBbVOMbpB3MqDVYKIEusc
GCU9ZFX9nQ4FL/PV1J34DulWi+/vUHfuxJVtU8S369OBI68lFlR3NQyBIPFMeOdz/vUUdhDAdINp
ohKyGIBTxDNER1XOwV6ZDd/Q1O7aeh/H5bSU61/BI1SvgThFxX40x1HQe1tyKkGiZikVRZsjvDW6
iUOX1WKqw6XDZy9chjtBJuDM0jPk03gcqho0aiWUCjAPBXZ34zTpeI7en9EF0Zdco+rN3YphyTlS
U0E8YNnEuBnATpfPDzJgMhZetqSg/KR99+dC0vI+WiQV1GiBzNXVDPJipgRzk2FBm+5NX2K8G428
CYFWPSImXPml8XZ3nJJ9uraxrmcK6qN/xcT55EOTSE41gYGG9nTVahm76LBwaFdhy7qnx+RJ9o40
A3wn3IigBwD1zwpCLhkia4WPlsDProIEDKVb53lF/CvMyXZMxug4ialpQFuUWPeROq1uxCIhAk4b
Ot5qPmUNqwj+PrqPBOBXPxH5earj2xYSXQEyd0GrUpEdPKVF6Nn3wBsxN2FGc+kJBBBflasyJUBk
A1nWljHyFvcaDPfkj3SDkjJoQsGe7gd/phDtJpx1jp4+do8NmSdOPW+eG/OI3GN7prtObSoNhq/f
u+tY+o3rYCcgs7Ea9IgjEEnhNqWKhptQxxHP3qZugezm0v2KKBnQWyvz+pjucesnW0xk860eu+Vx
SFA4gkYGhkTDyCt7ibtZoTOxT5yOydRYdPAfjDQK8kHeLWUmw2/PL7XB1nd52+gleGPP2tKML+LS
OEiTV32sgyB68zx8bOjx5hWWO6DFn+eCrD8fpke0DLFLwOxTHbc3yelncMO2/iYLbgCbg4nqqvAj
Ro1FeWbJm3tzuEMbSXyQzhE66qjf8KGnix51BgflmYB55c5/mgzq3JODiDa/GBqALywHOLegCfLS
4/6qJX1O16x27m6NlXOKiG+bL/R6pdfvS1WgT7iLvjPS07w8zSIf5btl/jNjIYpxfH/Y9x94Umir
E8IJaypiIaMzGuo+iai6Z0WiqsfIdVlehdE9afBX9T6zTzskYnwJQuNtvBuqGDZkLLGyssoLPX8A
c5EuYc3Ymq789y1pxfXVDxvNWMd8sSqYiN4HomxTE7H/jDZqebTf5OrEBAXayn7aUA1g/WDSYs56
oVN7aWOUNivhk8XrcrH/P4hCx4rCcMzIYKw5zGt9aYsZtg4sgnc/3y8zYPXj+pMurKNM6R3a8YQ9
NlTK2pFkPAsHI6gG1FokfdJ5tOtkLrrzlxchAiwNn7fMmwpZirQTiNMtbZjuGWA4FQKDN19pfAkn
RLdf8V1EHFnQC+g8ngr7uhpZL7oGGSbtBcKjgfgDXhzPxrrA/ZAky094NFJ+8G5RHsaGY0yevr8P
pvG4CR27NBz+gh3/B5kIvXgPnJX8zRk3fRndqH8T0gotA29HJ29eLLJ+qAFXLtF5myFbV5dXe5EL
FuJoM8LeZo2qhpE3o3AfMStqoOqgEi8tsPLTLMkvpSObbOHBPA5ufTH7c9lzyoeazh8KtVEZSF5n
IpkJVqUzFC7cbyXvAcLyMNBn4CPM8DpZp/fRdYbmZzW2a3eEyDSvrnrh/XQ94/WxIOzDYBpdSWw4
DhBMvdni7Z5JAoKjtMjS0wrcqTvR2j3lhuH505hodh0XLLwIsD4RuwpIrKU2Uc8hNv+9rVROe5iy
wiTzOcPr1Tt2Cz/i8NqFTxK2H5lQaMKiamXBjAq8n54cUFAOrGNAGEPMio3Rq8gQICh+R1KK9Par
DXVHZ5kK4iF7zb7gQW0x5Ej8BCtuQCmNNabOnSCmHVzRG+7iWgIhkQdpbR9LJA/Wn/ObG25XxdKh
nD5k4xBdVN+XI/V6ML/GlKeGYqMtqfvKDvdY5gAwkLfo0g9Gb6RnnDuP/xzDhU5NIEYa700wfMh8
e3hXo9ZIqSs5DvNbaUeqYt51VFFxg8EQt92+Q5STCsBvHmBtQbBow97krrU21BPZx1XkHSXSTOz1
rq/nNNpu1/lK/vKIeu3ZNHz8BgOFPvHbH0lfuJUlOdNzl06IzbYVFAc3vL8Z0q+Qmvb1hh2D4Pns
pqAx9O18xbB0rp5aIjzhOdAXi6RbE7fv4+kDwue2nomwMp3EBcZUkXUmiYCAOQzw9wWSR1EJDjw9
dSkwyhbxtXqcwqXbt0vEX/8X/2hJRJ8DrjI9yEvVsNlwR3tR5/GbXJV3NcG+gpRJhGcT9+Ukjcll
3+yqZEbxD1oDglOlWJdXz0X8eX9wrKuZYQ6WTeHQiwyXz30LcsQwI3hfbcrKii7jNI6GXLBEjMsa
CGt05ncZwbxexStrPIBwZZJFqMurUqMElQVMVFAg4k/CTZEn6wkCTfZB3dJalQLUfDo/A/ejsbNB
hXIWnWscmqwVVf3vKirNiKc2ew24bOzilwDSNdMJn1HQVuTKf2zLRfh0xk5ssJzXnB1FK//jLBZf
JHKpxh17A1QiYWRm1TUXyZVQxewXUMpLU5f5N2jmw7ntWTyZBEvm4Bmuy4rR1LOasHB3As2sdmW+
ixHgYT2iF82wNKysBzV/MzxthvVtV+v8VpychovZhIAn1u+VjS5f/yy7hyuI2NaOZey3sDYlQN2t
bkCut7YcQJU8x2dlibS3v4coEpTOqL5j19Jwoui0CSPGF2+YdAydvaZHxPZIYQQV6jLINqCt0Veb
Ie0OOXobt29x46A/y1E8+gij784dPcbYJUxwqWXEe1R2oKKA6/kVM3NeO25wSxe/Z9HJAR4heDWT
CJog5mPIorVytgOAzfOLIlHjh065XnQfZCaHsEM1hh3m5mCcjvK8FOPjxJS5J4ulx1AyATqBjAfc
4qtxrM1HFIkBiVU2nMsW1023nqS6WepMeDXGxtxR1gsoQVM1mwujd1cVVKntMt6OfbganTHMzBGm
sxXGh1D627TNfSdkfS5nqYGjYevhuyOXXD5Jy7v/u/YdkJlURm7Qzj/evJGP8QPPW6HKjuV2hYjo
98TYwLcbJHfoMUfcV7L33ZZ0trSt1LLj+gA1PlEHPRx+3GRQYt2POEIoqhZrWFfhYeQFCMea3rkt
4of45kQLJVjxQ9DcUPlHA5WF5p9xp+GzKrhIkIo0D8OlCM+mny3BvRMfyMq7e5ofIt5SdpWcnRdG
z1q0o5xmi4frvyDn1FQev1vncfjQv2h4uOnR+P7Ya4IyiMy4VOEoP0CDkVE3WXFCeYJn0DDDXNku
uY9ykr0Onx9Bv4oe2URVYPthhM7+k4L8RcHh+BqNZ4M7uowk/rtyhjMnMlv8pSRzrhGhtMI/xwLD
agqc33ssXxCz6LUiQ9I3L2TatSbtZOU/bNRez0+oxhMgIJWhBF6B0T1yXZeaPYa1IHz2R1RgOi96
NYLK9iH3A5UguBwLvCfGlsc6hMMZEvKmuSphs6I63dtPhje2jUUz/ziYK84IdAkELdSgVRWCYTWb
eO8O2fWCXgxuYiesiLYGzOa4le6FmDLjqQoRCvf/lruC192ShGd3DBr8XKfn2t7W0OGJ2b26MHy4
uOd6EnLyK8aSpZ8dxsahGFlQ5LAhdNDu5b7mvW24qa3ru1/gUYLQW8N3hD6ELf7xYyeyuCw2XmVl
UclGr8OHDHj3c4Lnu8oFhppVauJdkoz495DJTEc5G0T+C4B+kgq/p+yu565iIO5jN4ekZWYsWpQI
OWFvZRKy+pUUoii3a3y72do4fURTDY2TUzwD0v4v1sKlbsI7HSFXOr3Whxf6pxFbyqgIQktaJnFo
B2do6g45HvZ8KQKBzRc91ikUVgdX7g7KmhZF2X80oQIO1kOKglfBwj6/NYe2fM1kdLRj+REWLuKR
YF4KrsaiEOc+VubawrBzyuk/IY06nyQdx32fcjIvT07UxlMy7D2J5Ld6OkUTste0ONCsjA24Hmnu
p4xZsxlC91FDYy4gnVC/pL+cbMKprNTjVlfPVJAoMOnKQ09slyF/U1HiXmwqGADm7LlrwQgpiZCy
DwLk5BLyCM4dn5qtRgadXCl5XpnEFp/4NuUXb7x/YGEW9d5k2EUlR4PfMF+twaP9txkQ1lLAQ5e6
b+jsxPHyuWy34eIuAaQXj2S+A2eQzJOamJQLvPPVnHIJP0Vzmm1XyWRlbt7NdeMXT543u7cJukn+
AIqxZL0fUqgby+R6rjpacqOA7MaAmcBxssKkZSxtuw5R8BZNwgAaqxhtf7Nh+AkUKiFykanXB7j+
DK2HsaEnj1BvAoadc9xkuUHTSVRLG99mY6KRk+Q4z9KASEUxBVuwCeT/HtEcmQa7dTH9my4hAuVC
7v7adlGQae4rDOg0iLVubWYU7x1u5rgvxXADpjZj8FZEav3K0EnjRM3vqqYhQAPViesC6MYvW3jX
TmWqSvwjnXHeCT18vE1OZU5uPDfJWk7FegcbK+e7FmEp+w9Tf6WuEPiBXxXMghf3dIwE2WfbiFEQ
Rz6ppEZ4zqqZxN+RBEteFFnbKxOqGb+i8EIRNYrLOAb6xpBiNdDFbKX4ajF/EHc2pxN9S5PuKVjB
3O06o3zyazOxzhE+QJDviTiVOyX8mmb5Ocj9Ix1PPGQVIJETiHL7qOuzgi9QCpWy6VPfa68MQ/mt
CPBtAt32gODVkVeu0CtmYrABy8x8k1CytoB+EcohcFZSay31HKcCCVS8y33XmcZ6yUEIEF2V3qRw
0RIz8yjT6Wi/Qa0p3ciYKBMe54c0GQoJfLw5tWx3KcCJoANjaaSGBucnj0HF1a/QehtiFp1xzBGm
WQlLY5rqwXYKjiVNQUO5L8cUioSXnVK8ANQSJmU7GQP1uZpJt0A3BvYT4DMXRPWS3Y9Bd2Fdt0NQ
LznNXUVsMhKUKgsz8OHj5MZdRUQFZhOuZQxnIs/TFGVnEUK1ek+u6vk3uGaV4yRRXBiG60/P9Kqu
mqGpBle1dXzeHgh+t9quE3We5PqG6Gs0NIBgbngI49Hgek70lD8voGAFekSPTDvvijRSn4YSUci7
BrBF48XuqeITXjWbOitEiHauaKa8lyENwKuk2H4S9frjoo8RDzEZR7engmzdXbSem3QcsclHr1Yu
bHFtbWQq0P5QmET1z/5gDb9zyzUx4THESJIJto76LOLiXTwM3NBTMwAA2vbd0qF63AoxXJC7bDiv
OKhI/v4tD6yQomw8fJ6RehSPkb0Mxx7K0+i3R7EdYSR5qQgfkmNJtU4g04CId3VnwoinCo60ajOq
q18Ou+pGlrB+aASmiw9mgVLSSNPAwSIhwNfc+OspHwyKncKMpLOgAi8TMRLz5CID+xX5PIlKKPNH
aQsvl/7Yv7EtQpgDSBEzftEql2WiRp2p6hIlU4fxIBTr65GXK4jCdBJbh0n/7Binhgol8GUIfQb+
A3g76D6XodFcg4M7korvWXMCUj+9rhJIiJPn9fFExU44QzC5yArpOKly2YqxyTETnk7fJMK+lztf
BPO8T6WQ4l5+Grql+e7jTPJReOT8v5xseF3FrxaHeXWd3lKDW7ITZk1HW1ll/kZ/USkAll1tgJ/K
tdYrI5GusOjOy4iUL7l/H1l0+qH4MX+bEpenTT85kf+4eQegviLI7wERQhi7uughl95vWM+jaE3j
IBqE2H4KjTkBAssQPeEAlwlLtEV4h9y1FE3LaHqdGpbnEgAHGQAr89O+w70yjzOaFh+T9FWheUNq
XovKbAC5OFn1DINWYG3O7pegh2bgWL8qnG0p6wD/qt59NbqexHMHGycwUEjOqPTEIs8vUjnMCmId
kgRzhgnf3C4SIwxEg/NncCuHwOiPY+l3utZDSvC0WHSsC9E52CzSNuFnTm0DkNrdjzJhILhGEZcF
rxXhFOShtSK32jG0mDTGUduPNndXjEWWuqPfXzm23hONSPRxKQpyThhsgMy5X/yQYU0jQC2Uy1AH
Zkw5zzP3m9+9ofhJ4IkNPM+nBZoAUIi7hXKlSfqxpqEpuQGzea2h6KzGK8cMUmLwQIPiLnvlpvTx
8wq64haWWejAXjDQTzbQzkU+sGZoPPlEkXmkoA2IU32FluAAZxIZXkAZ0KFc7jOg2R9msRTTVMXz
MOsrady6c68xgRC+iFccCxekQfVSJ2yXAosisXM0I19zjp+sNbse9iDMt1Dy/8Kb8fbjlEObBOcv
qBMSH9NGkZlTrmwvGzBnJ8Dld+fbZWJK6PPM2e7HbZv2NMBjAxfrx16bWlaoAFuMkyj+DP07qaYw
//IU/dV3EP+NHEIENXvSCDc4ERhKITngGd1JydJI4goKp/uzXqMxz3VrFoTGVOSHgnstNsh0t/xJ
8RVWHfufOumeW4zMr+u04T76ivajpxOh7a/DtDJV/lESot61GrSNxH3yc9PhSvNAYKb9JaDMnxIG
iOqCsRD580D+fa9Q6ptSvlEEAzf5Q+nLxALZd31EgQmp5fOsPHUJDQwhjBJ/G//NF2/QfyZNM9mk
+8AYtF1tpvM2MsH7Gv3u44x1WP5N/3PFqdUQjfYb468DpIpuyBRQPmy0p1Vk7ws+h+GoSYsiA/UU
tmH6I5UGtgi2i2+EBppiR+NszKOjBti0Me2J95BvS4RLpoPznSAEqg8yK0r6GMmlty0d+Px5vDsm
BNgQNSS3voJzYsaO82/2czSSs3krfqr9vR17GDW4RJA+32Rmubz759pK8dvBIG7XHOmU78V+zHpz
02hFLIYP+zDZWeZdvIT0n5MtTwdcNxTQao9y2cZno/QDikTKdnRPqzQ25bHbu7DoBvJXAwRsi6XG
1d5DbV7SLDvcdGa90po/U9FwJnlzIdegH+ggYYOOy3IP12fcjNZRhsbPw5xfeAa8QwW/YedlhuuB
5hZ8n4sfqc2L8BCV3ZMCL3nh0mFH0eXj9inrADF/MoBT7FxhCHgt4lzAaF48ywZ0OBas0fpU55zF
HK3V9bA3zNFzKKZ2bvm8yedNdj2OL1m96XR2aDIPSA55kFMfD6LqcKYVT6pRJUpymtBWfbcXda+b
evKNAmfLDja69r8jr4IGby0uxskp4M8Dl9ucXLAmblp3lzGGkNog11G7UFTSSE1HMlrRxoI/GoU8
iYWKKgyzEK6jwp9uxiANtABKUIplRWzs2SxflOT1Gtu1zlWjdf1RNwu8LZkQFoPhLTnjetqdsDf6
jjUmej3Q2q9D8ptbw2oJSsL0wKU0y4VttvzR0g1cSfnK60HAlnmYe3aljX0f51xsAHDKKVZoZHd6
/Eqzrt+YheTfbi308O05gv/kLSg+Nn9q6ReDStXKszVhZJESmbA4JuY1eCe+ReDbOy+FYRq99Yeh
YRB/rrx3HqcC3KYSYcgz3D1I6+O0HFZoJkKnevCL++gBoZyq/zC2s4O90m9363RyO6mHcwxsj9wf
uyh6kF+PrAxzAj4VvaKKntnCKEG+K1EvLjJ3QLyACuQOa33leIX6Xh/pc0fgblbr2S5nAETz/Jsi
ZWL/pA02qB6LrjlV5YhSU28gS9EC0bTmx34A57oCIucT0lwUMKLA1DM+x2j+Sf7/RmjNM1PjD9nx
pSo8NkCPQbaVnAMB7HvthzSqH099usxbJqvHisn12L5mUgBD2e2QzxUdXRpM/1lcfEJiC3vXZcXU
1TCDElAgKvwjQH4MJrlLL4xWyYpgZC7UPvR8pNPOAybkIKMXVM9wGZF5JbQRswLlPWUp3+fjxm6l
bYUXhe/374BxhRtQWM9GBumQiX1odYdPXHARrid9Qd7irCKZZGgEnp/mrlQ6ibDXFSwGUQ1j0pde
WWGiuIGxGEJ95aH6NHNx3R5dyOZuk8gMevj67vzh3ftWQdwy7ldVYcxCC0t8xQpvwZDAR9+XaEqZ
e45S3SQzGCNwYigOI5eam/57FSpTsDbKC8OlsZnNzGdXaWqlg9O/ridx82bOKobrVWuBtLVyEfzu
Gn3k/da1UreHgNAc67cPxUdV/+7Vmp0ihaxttlB/zWy/USei6GHmfv2zlGWLgxWZpbrO265Zsovp
62fM81uZ38gkbuOXFVogZ2bEeX4lYXqwuJupW3dJBUJyIZLZuXeKG44kwuUTJ8cUNDLKQ0u4SZKz
+Llutx0VLl2uQ5QPQ6d7G7LGZSUlOIJk8XKEAAvYsqBW1D2ducOJu+LRHCfvQxP1eaHtkMKIn+Ys
yHfbAR5vzTWJ998SelhIQhy/VNA5hxXbgke0tGYtdtzAGbsqtCm52EipvwC+02zvnNuXESD6Kbiq
1RrMYExyu+jMaxAe2FVPI9k8+xlRJX6WL+r/8RC2HegRkduTegzCa0aO6Qqq6TV0S7Yaf9H/eVas
+B96UjwcTRBgOrIUzBZBakvjUdhDFZYAXYoa9WQw3/FA2O9ui9x9m2Dh4BaxCGXJQ65J+fcFFpt2
jzUOBA8lJZF+3pAvYc+1pql4XWZUyQ1fsEAmSw/CGNJycqxV+8RxGlU1D3ZGt4HygriJa2F+GkGI
Knx/wGXdENW4sjR3NN0Pnezb9js9FU9ejbT9H8H85wZT4Z198A+foRrEY2ISI9pDHjHuATo6tDVG
sA3bUV4WE+vFgU+Vhle1PSbEiWwdUBkkzYTela9tYiVYYD29bN8Fk6Q1DFwsOP4Vpu5xZbeJFe1U
1WDLQN/zbGwaN7Yh0zjPElQa2KSQLENdrqSsy5J6FH/JWzro3KT7wbcPQMRVMreJ29hMHh4vEiyg
IVRvgJJqrqC/TCNQC81q9lqh1dc/MEvBhKIk1Ls3KYMPBbuhgClS3KujFoP5275vRbXFoCw8+EGi
LL+1G8b0ZMfSY7UaPD1jm1BrtlKKNuNy/CTQTNb8rNt/AHNTyKRmg8pZxdecB6/7Xg6jA+AGTgDy
tb0Jy4OSqyGVyl0ZXE/0nDZmwumPiTb1y6yFYDmKX3B5OBTRnTjU8SwhexqtC/R8q3WkLrjRiS7y
a09iz0vRyvOHLMhLKagum6PaJFNg3q5GAuBZCH2cjVN7yD/FMPuk8z3TDbvqzikT0wT2S/bn4QF0
9Jc5335KbB9ezZvnQPzW05vsuNMzGKrXVkTtkIcJSsf986EKZ8cj8JpNqEqgmOz77lg9+ydiDKw7
RBW8/uOQhqkCkOo1lFYsS9OzOk7YVV2j02ZWAME5PlOs0SIc3F2JIXqmxqS8BWv7FLCSzwR7amIQ
1JsbYz0AFVCfrKbdWVzNy+1hG+QywPogeV3g/khcdqRSgaPrFpI86heACfJu7K16lEN6adHPUnLE
kEA5vgrDh63E3wtPo9JgO13gu+ctbfYCx7VCcrUZHdFI5/kShVH2Qva4vl+Q5ocELeb8IZ8jRa7O
HPhoWPMF20iMwwweSHQM/lN9GFsuNXFq/OlXhdXuPJlw9Pfzoc93GASFVvObq2yeAAY+mxwXKdb4
VwAFPXYm2buFDaunB81LoVcANzuPdZTQ7UNaEqMjecyrQFP3EmfQ8Qf/6bb0yQfuRfNRxjaXEbA1
wUiz2gB3HH5xEPLJkK/XOD5GI288cuWve50WMQ8mwZthiyi6hAwqPoKXcbA2Yp8afeKplg8Qa325
/qx14ECb+dzmRqMP5eQuUGFB0p0V6dTs74KOf07PFog/Fd1uNabfWpeMkdKIAuYDUhM2uAUsw+mx
nDEqmu1FoMlGT0v0CRz2kibp2WG+2nOEbfe8X63gadLgzHSg4kgCuYite7XX0UjuiTq89Jxz3HMK
1Fr6t3D5Y/7/YM45vsDIpII8/W8HxZQeuefj5U29CMtsbswodJw8/tdMP/uZJNSpIh5bvV3VQUoQ
55DRsp9sDSTGlC8gwNxk1Xnm8bCHpA9ARPs8RzRFlB2dDq+jqc435g/XpPK5yr5Ca8MtORt3xNYW
uCjCtvYVm9ShBj1rq2G1R0RW2v0U/fhIlt76dTGI3AIWn2PUwGlD/FpO0SU/7dkrGJEvJtHOA86m
bCpthURhW2KdSOVSqbl2zNJ0dSdsDmLYZVGyiL2qZlllZ7SxCfN0inrQY5amjqxohcMZn7uIH6Le
SdwdaOF3m5xtRcGB75UjE2tNaYJREnOaJydsLr9Vw6sFbRUB1j8tAFEu8nEdZ3a/vaJ75iub3mSC
BEG86zyiKtqU+tgmr9KXqfkr/9bMRrSXeWEFwFaGUMk7xm7wBtZ6y/3Gyy3YbbQDWSHxre/PYOf9
VqLMK5Q9P928p/djjRTGRea8ccR7+7mwXc9rVYznYttHinX4ZTCroKwSSmNvO25TyK+/9ECBn7Wd
qGC4BKA8T//ZIGZDo4GmXOpmaDlNxUp/y2CjKTBKK53u3qszWu5YdJR/ZukjiqwGRoJd0VtpOpvg
pO59PU/pCs1F+1wBu1pGB0/jwS10Q7jJUNddqhZuWcY5sIRunIAjb1/uMKWI45vqgDqgy6BBimha
pOjQEd3MYFpE5GRaB+6HiKur5qQZG7k3d95deSkUerP903tiPf89Vf0JVPR0zZjx7Ug1ENgJHoUk
xkdvEuVR06WFY76c132sfRvIgViTYOfr8JKfEtXrV2yAPNUMEBVeKuuwJ1ngltO4rhsO5kTzDQvZ
rKS3a0e8XbDmtZ5kzYwdcqE+/PkVA/Npo/6mt1o2a+HGeMuEOpZcTxyaJX11bPg7AIwq9fub5Y6L
FoXIqYqE0o0KVo8pBab35acHaVZG++LHHHWD9KE0ZZ5xNmf+qUVhk2AGrQZ/JUWGklIuUDXaVVb+
CNFYjOMvUj/dERcQlLDxEdTddfJrt86nm7VZMQqwa9c5sh2U5qN7YmnUOuQUlcXa/pCHPo7l485r
d4+ch3Yd+0LkYIetYQImRokrojmjDEMqF8r+Zb5oSvZqdQxf7NZeHaeqspao0g9wj2YxKrJunp8j
Fs3LwD81wilDcGc77bWHk07liSPgqK0eTJ7rmzZlJjrfaxPvwGEhA2Wjq+NS0UM3cYMegjBLb39S
Qo6Y3Hp2rPoo1gj0yKQAlYAie8uSSTRK+8Om0/NlnBddYO7IEkVRMZNLqbQfUK8Fa6FE/HLPL6bn
jLPvlKstfWkMOaEOPvfhHCeNQBVl/lutm4R7jv+9R/QIhXRqBgI5J+VHb76IJloaNjGHlgOq+X7U
HgWh+0GgCl+b2fsN4WILPy96AwYSSBNPc10fMiHJwrfHzbRneIkMk7xuKAZnm2gam5sTGukxrWO3
UcW87XT+jqNwsaaQqylaxIA67yks+qC0suoMfsxQOaPkodYDZ7ObHWGmb59zhkIwjJaOOpYPPbjZ
C64YtoLMxv1rCs0LM+Y3eWz0PCwXY+8k/qxMVmoRpq8al6QHhY0WdmiqXVxHel3HMZ3mPh3jdJyC
YDwYPHGR7ptC2ll9R/pGxS3qvNqNHF5GNTScaIxbGgTTgR53OloWhFf44uE+BhZ9QG4ZvglALOc6
P+k7wFfPpR46r5r/qVdhx3gLkoimSyt185Leb2eD/YPZ7aqNOe3Lqgx7NOhAaV5SnwurkavGKjdL
eRbe6X9GCPIkjL89w2ZnMbr3EmUcQQZdlCdGU1PD/E5AgCZ1QAarr9rZqQPxXG9BxO+wxXjZ3mF9
W/3qh7yYbB4kZnNPuJ4TSa7bLJREv+Cect8+zGuKuj7dmiBwOct8DTEGBhlYDLubtxxh3qlLjR43
CjFecQauTiF61X/TNTK7lnt2Br4BVu9u3xvRkZOCfHt8FOvYZYbhIaorAmEA15+klUUMVaRp10hZ
jrISi6u936wn0DmrLVqwwq9PWb5G5jkcaJuCFYiWcjlMXSb1PCCU17/kUQaQhynTEq9GY26UBE5O
ERW+f1SFAzPEinuJc3SIM6SnusLVfsj4erpjeBV6akMTwhovULxHow+iBIDp68DWRZEtAplmuls4
vS+m1GIxowQmUrjm2lGlcxXlw7237MWnMO0BrALUBFiXojTm/i15bhUJiNtn+trBXM3aLTgtzbxR
rjvhjs2uVq1fvJRdaRTAgboV5S/cFKujKtc5tt6g5cHxG+BAkX/AJVAzBwzNCCLHL2QzBCvcsH+k
v+wDzbYlinJS9eaKQ9U/0CZGGVrWqP3KXpladGEthFQP14OzWy2rykBX17KO8heV0KEd4IknxRyI
ahuDeqg1XCOvlobsOi+1Lre3uanpkX/lqoIXVJmobx+U9ZG44kV9hagyfZZFBnhb42au/fVbbo8z
4qivF47p8wmdnDnINF6Be01nyR1myJiUUe1kbrNDgwObFqJVxnY5Tk/teI064Hd614aPEPAbIkyY
R5QmcG4sxuSz/M56Z3xR3oIoeJpPrZRWCbFzssuFFZLVz3ozshc/y4ynbkV5XZiOWOKHVqaPNCNW
VmGzckcDOo8LUT610uCosSxrCKszqLNRAh8onCa9+hZBG2xNLiqhulB64eQOjrAB6kqRfLKhlo/u
V+GuoTJI2cYao71yA8+K74xedOZrmB0uMivKfc7zVcgomTbbFaeQM501XvDeS2yzgb2eJC75wnP9
xqOVx/KC2g+oA6qpmjx604Vcp3fca+7gZ2EX0JoVJDhxb4v28qRFlRU47QhLokYbZHsJhWR0LIb8
JwkDIPVQyv2dFg/mxX8vv6guw2/LbCb27y1VXUYIwNVu+B7doax5SfFf+EPqFTuwzHZjCsvi/dzR
w7OIA3z9hMyc1Cr0DiGOUlZlLI0Z0N9ozX8WOQg9cAwxt9opmLaXv58OptKBmLGkLoWQaO7e6/44
vmEXaMGYWKxi5IaPMwfZCgdKxqhHS46XB66ucQbf30ctlfqLQtDj0avPnz291OK5RNXnFVY819Fe
0tGj5YioDuKG2fFnCyLsvLM++bs8aQ5AC1OnpzaKgEoA5AIRKRmZvtV4n+dPvMYcNqLnCmU/HI7F
DQXw4+zTcslYw/4NnHK1lE0+0seGrj2bOAAUX/y7bo4ZtHmsDLoiRip8JCRlJDA/AtZMWH8GnHxw
cyurZ+bw2AbCSnP6N8dlvQQG3KFaHVK+SXnMna2pdvxMYkCQndetUOO6LW0GtTk2F/eKzwVl5JxP
m2oQ83EXMBDv+Uy2WYEO+JPD9ULuMiGjK1Kzut02w2/a8UgTTVO71ObLgRBUmxwOIQ5SC1EiUGmp
IFa3sTA4vOacI9bFzyC8uuoX1I/Q58Ijkgkv8WSKN74woCoV3O6A2sntpgoZfnCAa8DXmlj/i5Sl
EWgtQvZ7Xiv/fuwvMKderrbLv18PiwSWRo5D05WiHbiPdV/rSRK+7rTdCJ/ujn9sNacugc1PY/IX
12+anvHcuB5J5BkKi8s7vD67m/SxiXd+4ogbkKraIhvKsHqfzQgMCAIHlUFbJW8ZLegrKfCose+c
2fPpvcw2PQKRESR68mkVsPpNGAbd9bLuOXTBGExNtLtwf0ACFm4YDhPUXMbNuXJH+yGIPNNutgUD
MNnXeIA+hMQB1PdeGtmZXAjAt2PSQwSMDSQGYTwQTcqZenQqReAFTrWNQIeQAcdCgmfG7X/CqhTO
Nj5xlawnYjBlG6sURbrfA0Wqto7cp0SYh2PkobDnlkY5ZBlJNirUjcNLxRTIhIoT8lTzH9NxyGiu
qhaQJi4RGqgS43kfDv4gALQy5XMAMD80O0yNyvhThEIdLos+gj1/RhquFiNyOheTG9Akn4ZLHoMQ
F2V15iMGJMlTBMxaMlqDoBmw5VW/1PscQs6/hLh7w8IJUUTMEkmLArRfEDVLoMuZj+cypWP+7eSe
5JkDhtZyr6XIHEHLELm6uA6J06nWVLKd7A91VPF3npnXTDMO+wMD1v0gBQHqwqe7Y90JKbxVv/4h
rsLZZ/ZTsp3ge1wB3R0Z/WjpgQHTloxXYnpbuLdkNlxYPSFFc4Qz9x8C8/NA8d1Im8oPRWpiqETQ
XhDQSNPFZ24cmoUI5Q4f0l/b31tIrmI08onWazlGItt0t+0wsJ5g4DdJURjOTFidP4B1w3z9BIbC
EYZ16xa09qUJ9oGK5+WNeL2oZSNN3FAO7SLrLp/j21ZZsNuMkKZXAgdt+X4jIra5+6VSx++iPhxb
Tj70bKomeKFmQ0Z8qM/IFvBGnMFmXkkbt7tEVuDKSiNfgAfmNGGi7nELkE8iNdXjtJLj8jKgMYvH
c35YVaN1xce+uRZaOP7dY1NDjueungyYh794GsDt2DpnMlUSITYtjKpHVK+b7M4NKuJIh3oxwCQN
n048bYyxzrbk/TLsqUEJzL7exg4x5fplBsDE/8SkHcDR3U0k7GiKPFRd7cT8qCd0jH6/dWUOhPW1
ikXDodI+m9pXZHV8jkUP8J2kb/YmANs10/cUwdH4UY5Zey8v43RUjvBYcSclGstvhNAjwsdAToYF
X9h27ajFPaawEye1bfe+MnGwpxle5215kezIBS+E3Q0ba22tObOmzyQYYW5CtIpjFY+PJR61GMMT
anPqnxrYF0SEgR4E7YJfnoxnprdlqA+/3YothSoxOIp/ApA5G6k+I5WbJUAAtIzG5oq9FsVzsYVw
RZm3JaFuj4PHaijgvcHiX5uK99Ul/V9+Hx072EgVOvd4x+yDLk6ohqBz3EjmnkqJjowrweagktFm
I1zogdEwr2T4P2qy9ypoROieL9iFgW+r2YR6ZWWUXQO8p9VxjJMsb1xxzBuLqcUicLJAG8R/9Ael
5ilkg6J8/ltbn2YO1dKYsm1iSftj7LFidWrv17uh7hIE5u0n8wJf3izaq+aPM/K/jBiz93CB9LdO
Su7lDJwpo70jcUJ9iYkMugnO8Fk34vMAFvW3Zwlr9JfZpdRLXIn69TgoyAEfBPs2+EFgV/ZwNYvu
3HLe1QIzT2didIArLer3Igs8UIhWXcXHcKQ9mvw24jBWT/Baq2+cbPtuTClfYM0EVTrNnP3y5g52
4nhUfAbvmIsoIJB0n4PGPkXdzG7H7q4ldACT0KZC35l9XVXHlwX3FlO1R+qvFLh836OjKUe7g1Mx
nLcS7vRyBf7/JgdLtCvz9EGR/0w9ijd0KNGktMc5s5hb7F0PD0RwT8FMg4/jI2dlcrM+jj5+qaEO
AoZ6g25NWBivpgX4NVdo+0N/fHnxJkZCWir9+daKQM8Ye7i7pZFLjTbodAAx9JTKJ9HX9vtO8WDr
7I+3tNKKI5X/Fp4NfivIstSAE9BYLETfxF8cH33lrq/oG3X6cn5v7JLEYQ7zNHPQ0hENkYSwNS0c
7E4l3zL1gwH3cLZ+DQi8Wvl7rVlHdLrZLTKhYKmmpH9DyeHNAslg2h8SFLFhA79PhzpWJMSUVJ5d
XDdPJCii7pJ0PbpyWvEzkaFaeuyVNiRRVmcOQoPaOaO1niEf3bWGNBb7uQZuJ4aKb2IwiWWhfzRy
S0vrE5JROC0xiNp7CoxOBwp5o5LtBUb/Id08M1VxSaqkrPmCmi4lJUpmjx7+PUAeOSkTI7sK1UVA
QdBcWgVmrQVul8QitVZ5IBMfbVrNEXjnGPNA6pG5Vgfa6YwNsma71MgsIIgoWs4kt7j8biEqMiEt
pe4MSK1AlP43uw51Bb6JVp7MDSEER+D3q+yYhGeqPKnMLGor0YBGxeAgqXYBHWIT70YHeuPhaNTN
nzq7kjlo0ytnrjgB48UmT9Gn8zOylURcGs7mZ3f6xaod6z4/gPfE70fCZQZZ/2DPxu8tZ3MsqQHH
IjvKf8VU7f17FCVmygFlxSvsC9oTRy/53qQyXeVYQDOpqItCmQWXGfoy3NRHLIAaQm7fh9oGVZnE
dPhGmIsW2v+wLbqOVNRxIh9Fsk5Gp3VnQsalO5GWYQuJg9pIxMXMBPphM9SEubxcy+vBY6hjPWCn
yDOFS3edy0Zqh2FUgY3NrDpL0gx/iCqWG0yKJvvgjJbswVWwR8czCg0jx8lw/kNKV++q8r25GkKq
D/y5epRH2b0v4M4yp8wWosSOxKdWsyhpdFku9XM1YmCsq4fD3254O47R9EB3ayfwx2YwGkMsBIFP
IWhYk00uMC14ZuFLyhfxqyAa+xwPgtSDZnzGtI61BsCv5eD6jlzX8gPOlDr006x/dRjLhe3clEoW
7uDwLLtB3Lzuu281mQx9PvfoZgzvM5arGGU6OPYzDjalhaaNkMoI8lLjezvieTGQEHD/54tbrRkx
36I60Geh5PigN9+uHWvj6OJJ54ktHRJtNrpH3QG9XlKGaBwOm+b1UwZLCReO6lPMMUoxfHCcJehl
hu6eDV8tdcWpBRIw4Rd7VV6SIhjwGz9VgJRsBbm+phn+A+jZxUPAZT0xekGWgHQC2RasgCT6lGSk
xKGvXHZU8mjJl/EhIHQAXjgNDmSB6NnqVCKNbjodE7+qrpdgFXxJx5b/sl0dMDkJQ5aV/Ft6Xuff
mYLoN9JjtS5hpaAbmdFwLcRPfdgPmFCdCqGbVAhT+dOz+cvRWymiflKOnHqP+tVgn+b/o2UlaXi4
hANwYXCcCGcc9ruNqzSTcRFCZdbqcTS3E6KtVmoFfJn3dFYwAm0yCgw9+8qoxA4lFhYp/sctvdf1
T2TbBLmiFNm937IRdwtqLzrwSSIezsmTESwDDDeXziwKRkkU2IVNixXHhtKki5SpH7RDRVc7epl7
/0pwP41HY0ehN/fcm6qocRj/N6lsWglODFVklH+UxtG5WzYUiAW6dmJlNIPW2OkOr3TOz9sbfk/N
/N1r48qLLCK2asjS1nj3JEF/yJVAgc3lIh0t81y0EmHisRI05eM2wt5/YkdBqqAZMbIHQVGmkD9/
Br5n5OoMeiIQtJ0WfyAo//xFDx/ifboYevI1E7w/n5dzl/h4TA1I9cMxn2EYrUG6zQnQduQ3gkP+
6BwMJ2ZByvQ/3EeV6vfWCP+7nuSu+WC8Gr8U9rizsI87mLHrWvMaOOZx9jl+z5FGXhgLrRA0bX94
HeHuRw7apSeoxI1St+ceptPaULkfd4dyOK7t9gIYcn67lRsGAcn40+sFrFs3j9KwMA+aKtK++3Ob
4pEiHFmPr0sL14G1EE+2RInsGO5cDK4LXksbGefraEZRtT98sqy/WW+MjGpjHPqTe9GZ5UA13Ov8
c5tQkP7HN8AvnwB70C4yuG1zTKsgbvorSVWuPcOJyWYrYnA20q7vYRNlETugRH06geZvtHEafRp1
G25CpR2fkU+1rm8mr52GSsXCh+nlDARDnaVjWTavz3mPY7iYkV9hxJHZAXRv2R16XU6rPUFVjA0/
VOgSv219M5hXb1cuCkOm3A2vyrIvbawInvYlry3t8ti0UpV7MTyTqkUDwj/ZMVSRJXB6/70pL2CF
40dJVgcdOZnV/v7hNkkAZD/8JWIvHjxXCdOn9PzrRbUYFRvdKeQ/6VBYuAXNcsRIO2DVEQhnUpXl
tHz3/mMZzSaCjdpesLa3QNQlUIKVa7sKVAq0e4c8kLFTITuYM8jdOU1ge4MFgUEAPdYoDVwU9dXM
NyQt7jGgtl8GTI6QirThoJNB7w0TxADvW+ETPxTFLD8XH7Oqz0V6DnIoOV+syDbJKf8aFt+XFf7x
QYlBVi/lYk/rQEgzq7XZShHpvDPq/ma2ZpbUxN/5pN3BJXcBTLNR0PCj1qYsZ596rh8GF8rtlVEK
gvGGI4Vu2GlV9EgsfT/56f9DtvsTPVdDMhPfQ81Gw7g2ct3aWlneF2iMegZzYBmnSs8gtJjkOUyu
C5C95LLJrUwawZ3GzmFJDsecqHdQ/9ccp5rhhxbHZNwdcrglseut0wvaBe/IIA3B3q+aGL2CP6zK
RHfPX0CDDv4sBJqNEFS/j0wJpqm9cquBXTxupGruvoS3WCQD/jpOQYKC81zm21VacuqTEe3NP0ZM
LOLXwQeqEJZcCL76/y4b7PhRIf0L0xHKzREWtzw5jMeeUvQO7e0l854CiEg/2iucd16IcFCZIGcB
hEWeU6JtlxaEKTOE8jWp7uVjTGSwRb6rif/npLc/UL6ey1fTXJwlAS2nmR7PGSTncsIboMkziAWl
W6985DPOiR2j+Ry/iqxl8ubpSbb+3zGG2W99JDWRiaKfOFQ3EnlhXXi2Jtm4RhVZLgJhi5km1Or9
5aYNuXVA8yrmSQOKeOPzXqyRGs+3DOolkDxKqOkYfWjvzZ/l7KYyNRPzh3X818hUMXEoXu6ghRoo
N5fIIhGCawLF09s8IYB7X93zMhh6yMFD2u+L40AEFNCvvf4smShVoWlsv92JXI9Opfm+NZZYiWia
AdkPVKdNckCCsmeQPv+GrFl6gtWPbzjo/rVQJUXB11mAFJYAudAgNQAMifDn808Ei3Hi+vS0ZePK
Pr+3ooa0TdN/rTee2i0Xc+fI62S9abT8HtnPYiwxO/GQwa0saz9G7t3BUBSE6OGepiXq8x3GhpiB
M1zHSqE6rwUtUnBC0M/o79/RBtImcyL67tSqQ3vAXA9fbjeXF1JFtQmB/XVKG75t8aEr2Iw+s9cf
R//MUHIcEfxoBhjRfnSd6rUGaMs/UbThKEslWDxfAyFUpokmvIJYxKI6tSeMbnz5kPGvt2rrmd1R
q4jBF9JXfEGWHj8kLXHloD3woNPewCcZcyHpOx4nhkTlMUQHdh2uRAh59I++v7TFRveRJS5RmiQs
Pz2xNYH8VWlsBe1XprDN/sau+wp6QJGHgHcP35i4mtlmAaT5KG7OAtrLpzh/XKCw/l//JNjypfRj
dqUv6EkiR3CG8raTM/peiHBFZ5sczrWQ1+HQpZcd9t7YjlnbCVOJPQ3dPygu5QMQr8hDJ4yYZpH7
smDVFdrmocCsq7pzpvr8WVjp0OJLFBus0LJhV3ZEI8cE58F2Ke14alHFocIYYzm2hfXt6/wvTtRb
dBnVqsJKk6rwz0u1Q/+ODHIUoAQEvoTp3BK8jYzq7i9ZgXQV2m0ORUMxIfxHoGCwJKULQSK/2i+S
YnAZzCiCVhixp0ABCa3KXJjoO/eNGhDIBnqOEXD3OSGcI0VD8CaTaL1hmxe4r45demzUvui7a2VJ
enbqlO9tR2krsC24PSz3Dn8P+WDC9YqgMSAIKWr+0oNKVyUDlCAqZIUyl0LjTOScOWsWCth7ae0y
NHWcOBWcNhina2rG/OAjwCoLBa1edjA1cLMbKx+/7je8gwA2opvoq4EAxQyd83S1BcU8KaBfpYak
ssIny/a+kSEngLGkyWPGRJPaRfz6iOa+ic0cVbLFFJPKhHQSJfPh9nKS3a0o/vWwv+YBHzTt4nfD
cPNAn+7loFeAfy0ltQ5q6yuR6S24c/v9W7UvBuvmjGYR/qH4S7/eyWjWwL8OnjKxvR+kJXFTTpIC
g346HeYiKrE9rrlGpgRGLW/J6h9y+scXL8/4Osg+ALZhJ3tsTohJE52OK0BMvNKYgPo5L+1A2GBV
v6jGe4as1Jz7jzwqV4KrR5h4KjIV+Ub8eja2OlfXriGNBROq4BzbdqInkuh2Fx2xZKEcvnlvSzOa
71M7q6HR3IU8oMawXmY2OlM4IbWnuioBOiJuFanEsh9ivlfe2UGeE/ui4ASytYdUC8ilmqRP+kp9
ZXeAzeXwlNfZLftUUMwsTMMoBifSD8o+uv3VqwMfT9X407E9g2wEI5NPHbHs7kFeD/LnYtiyWm92
yGMOoewDx7Kk9KxCOYcuSxLXPTwNyJzrpjLOHhHADRWlOvkLBKRATiKs4V+EFSmMdDQQO0Q+oXtE
g4yOHFlMxx3Bd0qKf5BAOAFsvMASS2/ptLzrWlFIhlMtnhuVZoKmKDfJ9ieq+BO3C6FwNufkyDWT
kSaFarVJXF+Zoi3oxtrYp5+13sq+4JU80HIO2voIZuEoypNx3CDqMNckUx2s8NlYe0iS9vpGnAAv
48YV+VXjQy7UUr199L1qyK+vLHVt3j5NEUUePVWRwhvYgfMgeCw11QfprmgykXCR/Yvwy5tf8Vrp
hRerz6g9OpsBZepmf/FgJJ4nIXcTeXvnk04fe7xF4Zy71OJ0Mu9Gl363Rm9ErfrEAnH29J4dHENk
uC/2/G9NPOLwA0c42g7ZE2jaCfO+JvHKMMJKEJWlf7CHFpu+E5oaRXhjFea1i+dqEgPgYzypN79N
XFj8dQXdndDHcHja8GzDaqEMA1cZmvgJb+5TtTYto4wiw9ZXXYABSeeqJPTQWCO535UtgwsAkOew
dL2KuSUnphnm46OEq2IX6I4DQFl5Ft5IIw74VOzIpZaA6MN4FZEcGZkSamksWutk2qoRFStSsZF6
ETYAc3FAF4H6/PunWVBgCoZcugySYqvLaTFUFN8VlyE4HvRi8T28eWqydGqiKcYMUoNO5jhK+Tiq
4/b+aS7YE4jQp9YvQ0TKrdKZdCdo/mkjFuHu0HiFqydSslAXn9XZLfYL5q9q8Ozdhf6Bv51g9+MG
quWkCKEy4SPCBV+QMljJmd3pIj54ZiesGoh4H0Mhf3DHbSNzDpYIAdzf9jzAMyOdrr7Zb3gIGg+y
Rpd1zBpwW1SA/cBzSZ1YfD5FDGr/Y/NczYM+oYCbwVLkYljdWqWiI18f/BXgb+s4eQS993WotES3
z7MbsmP//gP/aAgZcbJrBWGq4zQFUQUA8q+eOUgNxqjC+Ps1EgbRpTt4nZqI3rcTs33nxJrfqd/+
uhUmY5smWmvj4Az92ZcfA4cSOMQU7/zyua+ulYqemD4PrO3Rr5BqjDEzBU3I7zdOh6remfdIVgaw
prsIli2Ij11cnIbPBSnhkQL2NtXTapRU2fb+7Q5BJBWTLkpvbBM6sEZXazmHfOJgUrY9zVpNPblR
3WHlf20V8rEM6qCSp92hQRYxLWkAHIyEfb0hKv56xzVAVh5V3g7diTuuBRAHcPRku8xbt2qJuLrl
QNpyTNEc4ZnH0mFw3fuy59MT7LPFtFMr5pD2eVMr3KnG7NTqaT9Jo4iyGv5qvjHdJsh4p4XakZMW
3zTeJss2OsYM60T+BdTcL/7KiZ66NGtde8nDFqN9xCTDaD3O6z6QqOyOihAvtuTzuy5vdrnViudp
CZQ2sMosDdcFP07x6RF/6kdMG6pveLumSlwBcPWlaaVUDcHnV2ekKCd+wy2nNcXSxa24E8B+tdaz
B/gCdHhMy2rB6r1yNLrpd8+dBcW4wQkphe8UxWSyxqcLczJEyFYrw8dFCpKsjl7RbuFGYeq6vGDP
VsNcLkFHZlKfivec/HLAC+YuYBKY+LPUqUY07ZuiBhMzim7jKCD4IMnCg5U6vn2gcBz/YlUkD5l4
cRRkn5KgPH6XYcicnjaoiC4qOfyyxwRj1fPiOojshCG69w0b1rDoLcOS6xXyyNgI+uailk8m1Yre
/zDLhXQbpIUzzS8lAFv+79HDKgNVJ4+DhpCFt/pDkY4Mkm0gD/g+SUaIS0SXCMJ7D6TyHIsF1FdT
s8PZPzhdPcsXy3/THGNvq9BWXss9f10ebEIUDq3dwpQP/G3tBkAdA9FJbrT3PdNpXdF3ET1nW3Eq
2Ibm0xFP43ASUrPol/gIutTs2MTp5XH2NKZcNPrjBCEzE3bEv0jMmTkxSua7oQ0nmg3PXe85KVGV
SqZUvh9/h3DOHQdNDvjwf+w5uKGeGFKG2uCGP+XcuAg8EikTXdvOO8CmLkokGnehnG3h0xhgdZtM
/9a3avKWAY3MPpue3PAh1jyR8r6S7FUKJM2CbsTFAKotEGq+awyTffyWgvetejRVaHeLVyCR3J+x
5x3lThqCXNgj04oKAJdPeEugldulSnWNSMFoGt6O70iDvFftln+Ik9zkuwWPGeKdIcc09d4KSwvb
/SbuMUBtUvrPPYyL3JOctD1WY/ucLPy7Gbj/net0rzeNiD13FVIS5gwCsncM9xx/MsWo+6mGzYcd
+Zu8i+0onlME8tpdjXwepV+Trec1SetwO05XIIwUQPJewoATjQa9xq81pQkRk4OTZwNt0g4pLSKc
i/0IpjM+rCwEe0qaY8qnUn/F6NNK4N9LxIYGTywkKGBxgrqWEpy0NdRpG5PZaJj4GmAY8Bdh3UxY
q4qXWnnsiUIxhR08qETmetmTO6eFjmbEZEGUfC+HOOO8MU6zVkd11z/P+u+WxPoFCIpXI6NERmzC
n3O4HXZxFDKQlAWpa+lLlBVmLwvLTPn7qORcfxBZoJac9VuI/GClw1BHubCm15mGND3z6hoa8JOo
UPXgIBeLgfIJSTt76LKSZJpkzB6GYxn+kCiS3N61i3bjQ45xRmJzNc0/MnIoPtm+S2ID/b0pZepc
CQddrFhwM/4YirfYCDjQdjD8lMvQDnWAtBhC9nPMDoIDL8YdFP+SCY3SIS7hP6FqumKoq95Kp0TB
yAa2hWmjCq1gUpEmjC5zHWjMNcG2E911M5It2UJrLpTMZzoYM6orHLFLa1nU6PDTZ4zB/Cy9GHaT
YW1KoFaWUsYjqgfVhzZ+1iXS4LZkqVBOUUy8dG7dkZBbH1QZBOK7nPM0nAlMt6QdSP/AWTtecxgx
CJ+rr+705buPoKBHHuCPxa6Zj68BwPlFvgHfQWDFdxCd0rfXexo3dhSVaTQNosFHPc2Smy9mOEcK
W5h43MgXoonpr0xyElPpofJ69mhVnETxHQxaMpZELl+F7DLPtPJIXIgs+nOls7cf8srbkumh0vDJ
yNb0emrLCXd2JrtvdM+EPHU6ZvKRKC7WdVrizsk4jm5GOhe0cnk3Ny+nOZBGEd4uryNzoJrKDTmF
vMIJ3RHtKb2djGhCRx/xGFu9vUEDSYBlRLi0vOCJS/nBSimoh+xErnS4rbGWbL376iLjddeKb95g
Qf/77OpH3+nZ5xtJdhtQCw1uYCNcoQRBjnES2IRE0NfwukEELXXnP/MMD/c8LzF/xEecsfVCT57L
KKpunnR9ysK/eigTPh3Bx0USUCFQZFt26blRsx/R0eS3Y2x/8pqX9xdbNv4c3VS7z2JVIGpnL/Un
ypAyj5tdgHcwbXxm3gWz49tN35hc4Nw99VyRUVuax5nLgskc8kTddiKVt6nLJjbAU+7x56y2GnYL
ni/iBTL3K89atyElD5M0GlyAxtORovPZ0JMXarGQhFclquY7v5+9OfMdRoatjn3vcsXBZ1pRNgm/
8GuOHbl1M8CC/ALRIiKEnGsp++5cQKBy6cdbRhZzhRAdsnC/SpOl8yzZSiQAyreCO6jiQjBJ0k30
oY992d0lKYDi+UDj94sMGarzhnpjKMICk000TGuuJR1x5LgKttU2dI8eDUiKWF9INd9A403mtL8B
CJfue/evwnjiE2EeCnokVfgmEcUNqnZcIqiRjNIH6sL9kjUE2X9rXjMPAYyheY/57Yh9ISwYUnGj
8X3nB3YKvWzoot1WlBrDDPJztb8JZ/4VxORnCDqzwX9u9yIewWY2aBm1lV08RPEhfxWo3/AOxt0B
poBhSwi3EMeF2JlvDziC8Ua+e8GOmzO6mmh+PGPEoCjs0wQkCSud6NPUnyaT9SNmiwsEFXUNXFqM
Zfu1uax/ejaiEQ67OkSiEUAE+Sgcl8VEYUFxmo94iq4kaKsZzWpSlHOB9KI9QTP+3ch62IOgG0k7
WxDMM6w8S/i0KWvhe59zUcIXe3aS2MBcldn41t64KahXpXtBHmtd6YDY6q9XOg03ow5750jTfbz2
3/+l9AGJsb+YgbiT9qFX6eClvrXEgdAaAxeAEZKvP+kL0qNfeV6crJ4gxei3wJhgScOl74T5IT8M
fkzRe518k8t/BGz6lX5yig/jFWn7QGgdBOLD0/GKERtZLJLA9Dz1zwB7U29W0Rs1479qKViAnYcb
+aSm3JD1XeN124RwlDL3Fse55xzFheqZsp5Hf6HdygPCE8X50m54r43ylI6dc5u8NXCtNApO/3B8
Q276d3z1Q8Aa6sJ3h5WMcEGWSKUoPb1WjDksONalnV8maCaVmse+yp65Zuuip/n9wNgzjtOuceKD
eBFECe2SeXexRDUdWnkUfGRsFbwtT6w11+eWVM8KmVDQg0swhCzh1UkuX54aiHJ4Zb35CJOteDac
S4ggsfScoCdYDTZboU15tAJ2/f+57yxND/oxyew7JkPhPgVlDQ29/+zbewNXpxLyx+KQDSswqd9W
s/ruDMAtjD4MgPNGB/lBuuBy7Pc5J/q4xT3zIyBXgJByWgZ1mwM0LULxlvF32tjlixBSUJ8RCyjU
hI7h2UL28JSJ7OZNfwIeq3hRrnYIdtPdGCWX9oYKlJn9wjf9fITmfSF46Dp9iViWp/HyfyKtGyzB
XE0MBR2XyfA86gdbGm8+dDW9TIcHqRrijIEBMm22rAjKIKC5EboLfmSyB3Xj7kHXOMSGsRmzaPXs
Qtw54KhwKQnMTeTNIq0SeqfNmkTAvdpvs6zAfgyDpP4YTlzrzoWotG4RvlQASj+nAvQ78TZ1SIdT
Ak/Suvn5cM629oXxqIqLQVdTKxYdpjbWabIbheqrHqDND5oGWcmMPe3BcxPJSKsVFMsrPerqSN16
w00Oq1l1+T88e3iZ17rjxKYa1iVdbM++S46UU2SD/H0gB5abd3jTUkEqGGPL3kj2stTVdX1hnQJP
h7iiuUi7EwywoEMeQ+XsjRwT0lPifNbAY6eNCibk30Doh1jwaq7sQR+BXZbM3L/qBWs0gu1lGPuY
RIMWkJdQyI8x8W8xJoGxMZ+WX/OzHUEvSMyx3DSZU/JWh3Dct/38QJ4hp8KZrj6gcQ4E5yB2m5md
uF0wYHcbiidp9nXqjpL2SET4sNrkGbXGE5Yx13f7Gz4wrTGTyT+tmPvcCTuH9ravwt1dK5Y64Zfj
Qhz4JQbm7JtCtTD8PwoPOWjQ8RvoEHyi65A7jRl/T73XbN0KAq4nLDczTFbMHx6lFaDsjfq2bYmC
STzs55wNrmPfh6xoN1Wr0Iz4sqDBODsnxaD0KOVWVupUmNVHdNsLX/w9jJbKZBp+rsJ7t6ptafcu
XL/lrcL83+29dvvvx315/IaDjxIPntuYBq/UoBWgQq2LfWtTw1cSlCLgSfRi0tR73GVEnWTzoFkU
9dvRTZDDpNWCuqFwC8SGb4TZarr76O/QrlUqSfZcUMAovWySR9XPJuZi2JibGy5Na8LiH1Kelwxe
hwx9l0ycm2TB8QIVNMpO5zSiruYmPYud/pCGIuQeNvEM9SookogXDFiZR193A0lyLjIGjQXcbPHT
o5KT8/B0B2nzRADvClxbb9j/VRhy5hhGzm/hCev275xEj4ICT6K2mB0mZ3db+UXgK9mY02HiUnnN
S8IMou771lrmujfHGP/8Q5IpgokwkDJLJ0V2b98EDWvdxyhhXHEa/Iq8GsgOr5jg+VOlGbgecPyS
7ugRQiAaLM+coG/iVKtBSn+vLV0exJMj1DU38zEZN6NfIrRb0K2iZ2dGClPrMqUqXhQDfXbYsUEO
8vgxZVEuVRrtqzFSxuCUYDrVYmnrq4P555U7GPGPdZfpizOni5SY2yl5HtwXY9L9+VfLSBVruYtw
CsciCXr/XqVR8OaI/RGbfo7aXbMM3URMpTGszYAVZe+himlcLnF+ExpEFhsGCtGTPQLQ9w/oIeEB
xt7aSK4cvq3CZb8C4fFnU3JX94Vc6ROhYKIv/FfQ6LvmNEsRGkpkt3XjNNN53xQLUdoL9FMFQ7ZK
lFaENcHhLwpVenij1xrKZP1TVH+KjyeMv5zQJih8wYBCkGggSnucPbYSe87DQl5SBP1qHk4dQSSq
ZmdftnkoxKpSdaUfebqV41z5EtpBzfMGhKegPDUr2voAKJOMXs3IahLfqx4UxQWEzNtZ0KpPCkuK
HxV+ZfCqMMkQQqEJMfAFbgOHO4XtrbwWlCIgK5wgK67GfVRj0JEVshGtQJu2Gek574joOL/qWq+D
F+KxvH/DJ9ciYuPlWNwP5KRadBm+DDGQpi2P0pvoDX70nW1ihr1uZmQ55OxnNLwYF9ZInBdWv0iu
XWOIBk9IRYGB1KQrJ3tw+zvC+DFrDTG9HvRti3oDhgY/gsyzfYRisl5ZlSORj11ISINAZxW+tPbz
cpZVighcCAbYr1dQYNCnhhg32ZXgBn+D+Z3hSGMa+o7RrQJ5c2qyhFPxu0lR/J/vnilnjNHqpatu
Px2MrY+WlXozqCk8554tVd5BKmRNywJNCkyr2sEqhhG5gS89Gu8hD2CLO51DiEQ71q60anir8y5s
uD9CIpIf4bUpLXG4cB1T38lat7QhMKd4YGiBUhs2kTeKN2diLhhdF6/H0cHJFQ255TIuyszbAjNw
3lpHGcXnIWj+9tsuUSNGH9+EUrUSC3G6awJ3Hsdk7+2jaffNlux8ZwHokOveZtAOojCw7/TEZnR5
AeBeySKUCEsw9HSGl/ygigtqEF70QPuQTKTI6eV8XYphaAqll2XCxxSJJYmkGFQ5wXXGlmkntVsu
reKFwaJPGM6t+kmb5QPM9U1YdUEjDUtMibNy7xHQnzXZGHn7qknZ8a1IHEnmuVNY8hCpTAm7EV/e
I/DIQUvOrHCM4LjbGM702fSkIYbjPPTKkGLOjhP9CZje+dA/IVutr/6vkizOTpn6jJO0z7H+Ss9a
LD2zk4LZydd+9Hupo2cXYaKvCiedTjdQg2loatQfpaDBet+ZMWV5HymeXkhudIeLnG0UflJsOl5w
ueDX2MB7rYSeozsdMS+bRTtW3E/CpvDNOMkfkzFltVPYt3+EQaU0WdPkWpF/BFd3kbOsg5bbI9YM
SG3EYEwklapSz3e6KsaIQ41JAOhVQL4e5KyqAT85lSdzfI/D32XOE5agxHhRoAwCbx56qHBUmyrT
VkNJh9hpydUyT0NuCuKHukadFQgHe5y8pua/PADcbymrovmXB7yAjU/LH4oWRRU/Uw9ENSatkKZN
Em/kfHL1NbX811Bn18maCui67t0K6DkRrPKv6c3/NzQ0SZIf3iUA5FFEapWbQDSRxkNl6BeZ7El6
jZCr5GOX/uS0peZ7pm/a8vhQKKR+Cwa+nR/9ipXvrb50YAbZMmTrXr1ub8Pc2jRLHSd3wGYUIWZZ
PRquzJQ6alXtx2iRStV89PJZba+F2sj+6YWSDyW17Ml0vfvD3MMPlE3ALHlskxtQrBfeFXi4AeIW
gz2urikLvTV0pfS6t4ECfkMt2l0GOeFkdWXHDhEdHSx8icaDPDHg7qVvGLERGSmmBGdUHAfrxELD
v9nmA+6o0DI4eAJaPRE+Q8EdMkkki07Upblg+GtD2X9TM0A1L6/mukR4syy+1kRZIj9DT9qPSa2O
TIM1IAiZNF7OH0AkJY8stumWsrS85X+vyJ1pkAAbhrPDVmP+K2cMOJ0KN70sJLpUlewRdr50fFu2
6BLGASoc3HYgRliz5mK2i5FFzeSIE6Gh/CNHrr3QUC1Tbn93jAg1rXCfpkNjSJkmcHAbR5JWvEcp
YQDGWy/BxPHcqM0n1YfTMAkQhtuTfiGxEGCQCMV6kgt8Dbldek6vRebu0PhdzJ9Dv1nzj8RJtZFg
rnhfGLQ+R9Jd0SvfPsJIGcoyIFp2zTTp4UooyopcnQteBYGQ0PNppbCw+eIJvaaBXAKHrPxIDIM0
lOdxFN6mLhL70Bm8qniWvJH9Er33qlVoxuHZ3KRy0PYAOz2qSXR09Bx687GE5k1Y2+B4/zyRPfwc
vRGuRi7wV4741cJz46n9XV8CMVBTTx0SShwpY3veEdYBq2UxRGxXYldeon79GGQBUCoTvup/G+OP
UU+wb8tIaGNNhEpEfSg6EqLLAVOttu3Tjf0krlB/a2yTKbuChyr0YpsSp3j6P5uRVYiWYxvlriCB
19uprZ4zAClXD4qiWuzhgOqriDghDfr1cgVE5JglDEJp+8cUCR9iw0zx6re6mxTXMeE515VbPWXU
+whpp+Qx55Hm4qhipaW9jcvzho1fns7nU8UwNDzN0+ucXfj2v1EXkjUGn08Gbh3fswzxBRQUyMDF
qkgAKioL0dnK9oV4llkxmHxQpvueqawFxuSZRskKIzIIQnAjpJhCb4YZmcbfHs8YZ5Cy6EB/tJM0
9BHCp9lHSY1y91PWHd8S6uQfyehRLFspRhS9+iBGzDYZes9Cq+E4Jd4UPB0yBQmbRCCVT50GcMGg
LEC4jwaSxRRnMJx+o2p7WO0N0suCVTu0RcjuCMeiViB2y83sr//enWxGQ//GsKMAO+fpS+MwSzGi
nh9PuOxRMizU9qp7h5pVwzvIz21h1jZtw+sRBtkmF3J1pHXQSDOpTjbcbgnTOM54O96fte3BFzRU
hHMsIveDd9DZI0/J36mPvKIOxaKgplPSAAjoMOtYtL1m+NZCWOXVuvYTKKd0b6Cyz9ya7GBzc5IJ
sTAkPPgGsXmAuAEPiQnp3mpOI5SmOjnJstif2ztQh6ne27dDPhPtQ3Cd43HBz/BKH/00nuRXdsGn
EU9vglg7YUk94mjXK4pshTpgHB2Q9FoEHrNZ7pbb3KZ9vvTQI10p49N7kZShtXfccRXVFwmvNgju
r1rbde10lPUmBZRG7iMf1pDUXzlUV0DqJ5/bugvCenexs2l3mPRCs0frZd/oOf2U9lW74Cl6/yXi
gafTENZSs6EH/AaRY4qUxAWwPBoS9BchIAMzzaFu/F047gtEZqL9+LeS1g3k3EAC2dDaVrT3DA00
v3xlK+QcTMVHsl3rsGrDRtgKWzBee01QUzFButZCTuQxiQFR3mf94uUKlLOYsIg6jRSqV0SbYfqo
r2DU7zAnG8q3BqzJnJolcNAiYRx9uuJytNo0d8EcERGyY33xJgHL6A2qdgN+SWMPtDMPL8oNJn5f
+s/yzBk5hkOPOhdP2D5ud+dxP5AXd/UrJkVlfp28eGTxmVxkdqP4QMwBa3q+Eu1KNQJxf40PyXBt
ooCOv4wCJAJMsFI0B6MOngmzk+FOTB/DWIvenYh3i8fpblVhvOrN4ar34NtZxUXzreEaA8pmTBe6
NcRIVf1h6zkACgieYFzUUcF3+4gQrrnRZXIWS+MUVtiKGqe1x7nCdez5JcG8fLanbDavg0V38W1Z
W3G4ZXDGM3gHwXssKtgx0Gi9EREj/SV9+RmaWqTOg3ECNGHzNhoKc9aBbjEhwzUeiVP9BJRpYR5L
gk1PQ/eeE9GYVHNw2vjJIJqXtN4bF0O9G9paSlOeCefhrr4FKIZSW+aujWjU6XsJdpsP8OQnLNB/
fsPPoiXjuNSiyaF2lJeNrxrfsY4q11ANl1v/BrUtOp5LF/YBXLmUFv77sr7YxZQ4IO/rgM7HtWeZ
swjLx8xsBbS2MJEiPXEBZ2YGYMljytiA/lKYL6S+rRPq0jkboo3Jr2vKOARf7CY4OBMfitt8I7DF
ciTsx1Dnl5HmUepxJwAKr1CSXg0azws03C9y58qIUJTGBXXmMP0w0vq7fMkuS9tR4ziqCbFvxFxq
MBo78paFELKvQfLP88lxJEfVJi/JjrUuAVXIxm9p1xK0djM8JBtGozWj01HNLmqwvtxqtZrRgW4K
ZTnOybypPAwgr8pk3d3hzq0EbGd66rlYEnFG6dTQLwDEygpOmRuY2sLzeTQH0GhvUtGJ6IpnhFDo
/iRyVdcgufinoXDuxoWkBy8MH3vGLCo4SDZ7edVnNN4uIzE9wEwKnPL3qzTsoInT/F4W9cVoSztA
ha7pQSPGgzRucjm4lPEDGLCByNKG+lIG0laWcYkcyW4hbbAJVGDuxoZ56XsOpsNFz/YnVwZnBfb+
4B35ddDk/74oA+QOLr+ob1X5GNZWUtYG9yUtdtiVHj7XPX2GJ8PAy6IugWIY7OKTG+N1p61lSkWu
iZ7JWHs0GR5lw2fsT0Y+oOJ8DDz2X5KefK7Up3d+iC6lLrak/y5hF0sYlIk74FK7N4d0I19KLMVB
kVRJvKNOECv1KStombjRvJb1PvqExaa3xXz0mtDpLDJteT591BqMhG7IkziFdlBRE960lHqS1rjU
WHCYX7ejhdM4l6LbJwUgOQTog6yhjlcr/GkPvFLxVzyNM1P95B4SWYeiRHhAcauWm12LdLN6kD/9
cg6yfNqa5cW3vo+ROXIFCsY9jxsh0HRghRoiJllzgAH4+twDrKfqAXaDHZhpCY+lMYEzy00u8WcF
KUPHdbVyqkyBJbnA3tvzzSKlT6X5Aad0zALf3g2DgTyiiqdTaFyAim9NBMmieU69gRB8qmqNiBfE
bOqkK3JoRWAj0sgYwKoBCywQjJFDj5qqcS1VvnGf6ymbgVphoxfyAlsmMx2hVLzBpVNBwOj1smSS
3EHAI/X4ltcKt4Jp1mPWvUBB/IR582UoWdKZXQipHmSTcoYwW0ETo4FNf+KMcbEdm7+eSjU17/BH
VpODXhQrA8FyUqL+8Gc1IZ2/L7iBdx9U1rp8p/zdZ6qLonT1SXiWk/1S2JYzx91a6hitjoU7Ysas
cRE4sdarvzklOJhWRONl/CcG+Y2MsVUOZM40ZAucwuRmBKPsr6WbQTfeDp1jhUS7dKagfXIW/eIm
MoERXuTR8PFpSxZgSXNgUXoXU7tjVaYvUCFpCdPlZprGQ2jfVvQyAVLdQgIjRUzwK+vIH+Rr9mDV
iGZVfYco6A1l/eOQ1eH4HkcUdsY31OnNIg63HUux+OzgxjbdXOlvifoRO0NRVPD7ZdH/Deo4axy+
e4zyRXsbxoNOCPW4CbWE12BSUALtIRiGIGTbtc8CdDqYiBJKNHZE180nEFOrtLZf/ize9V0LsX7t
9S9kfTTbVqlQBIpSdOIVOxOqApthajFovrvhDHD3pF2AY7xKty6kHJ+NOteTW8w29/oBfQhIT7gX
OIMKWcGmm4awPvWCsYn6BG5KAstnc7A8If+6kq3Gd9sAaqUBv5tbK0LgcbdHliPQyRS7kfd6RuDY
QTVyQDXbvn+/8F+pjzZEGX2lFcCDFPcGRWrb1COh+GJd8SqgB++Q9Rr376tzjHbbaONwvV6KIcax
MELVkpZiImdrza8LglUwo85jWdUnpEWFgXiutxwUjeSye96pZnOx2DGJ9sqOrzMp7jBIm4k1kSrc
ZMm9ldy9+yBCjVR0Qo0ThtlH9whxf87QceCfIEQMebVL8W+3wP/IAGXqdN1Pxyscrwc+uAidC7Hy
w+xYt8r8Q54PlFA8dvoYSiK4MvfeA92KQYP9ZB+x97h0A6s6/yfTzqeFZAGj7qr2C2J1SotOBhyU
Fn1AY3puStFO/UwynKTGNf4W0VvlCf5FNvPN8hQINx23vW1FrG5PRdHJv/CScVNXggMkUlSOP5ES
QGCn0EtyrhVo0WjhqjtZsZ4PcAM71aFdc4d0rR46B47f610mv1itIRAenwbYOEIzGe+pTbknbouC
8wb6Umn+l+vyJzLy6d8e2VDb0zqHPGeb9K3aiGdocNV3GDZiOeYKtx2mJNmFzMVhSbtcGZ27ArLb
m0y4C7FydNqYwIEZsDfrO0F2K3J6/nvnbOUfsO5wY+/cPCa4J9JVGfrgLYoJkMd7o4aTlI8aRZ8F
lUxo6UJBWyHin9tHd6wGaj6HAI3+cxpj+yrPbVxPcLqFNeaihwv+xHoUkBuptL9WtuL/ZzOtsnRI
Vf/Z23IfBaOccUgfEDM+5Qqs8hkmp52EFOI3gRWslrFt9tbzkn5Wzp+0h5Pm4V7d7X+tontTnB+i
JVjwZX7JddhR/QedyREk7ZON1Fu8bRR1r93q9rc5Yh2EWKMPF9hdR3p8r3UOQ+tj/C0cir5n7WCV
kWuCRVZaYKsZOvYdluoeWD0SG3WDpR7S6Y1hvCNLdJq+JPMT0xcnLSo16hD1MkQKZ8wO/MKqcrp3
HC/xp7BvVPpxxcF+EmvW0ZDce6GWosuAjdsAgM8t/3vFEY/Ufce54WeKw5Ma9hxU83cphKNl6Z0u
Uv2EUBdP0WeGMt/EG0HNsrTt9Sje0hdijkALsXzvHNTib6ut7R8VO+YLZUNGmNrPNXvXELO2+iqj
JsAxs/S8v+eSFYa4GYwuUyn9oI/oP45Cj9KRsn3Vvo5R82kKdSwiEe/kKniCoEQEYTSOC9ApieP4
5MCUozdmCXNWEQnlM4l+vgZdh+EGYkPoJ0XIJRjbpYOyMXa9vwm3ZAHh0kST7UBwRusgxwKp4ou8
XfgIWexO0fZrMajtKNergi/ufuVYcgJNwIRw6VsVOv38trQeuvGMyQokpeai+Ps2Wsud3UFDJHU9
lXJawDueIQbz4XCmLjXN1+s1EnL250Ls7M3u0DH4StDCmIJ0fIGzCXmPNM6qOJZZMJB7x25rfoRG
OgXI73HyGfmX959JJtoM2PiDxC6tBb6+OHbnJRKL0aYGjLb6i0CYLMCRggPjjAmycbloz969oOBC
2FSMl+3gEmNP05zkG2JK65w96+6OqyyQ/bgKckDQKpi8FzjTQGCFrWi6DShc7q116K1hgQr2w0eC
w1XfnHSXXGf3iH226ln85No5RcoJqfEF9FA0ogKZZ/hjiZ1qdppaaWAyvPF7yvk9YwFqDIOCX3he
5cgX44IjKOg1ca04xFDDQQoUb1B/xW6fLCnbIEWMkygmuuvW+X6ZO+QbQFCduJVqT3mu3HykpGEj
TApyw/4jkzPYev2dYvgqg4c9l8H1C5cl9f66t20xzsH+y8D+4VNsFXGpuWZhN0ZPiv7d4NCmDOGJ
HiKGwT4btxp6Web1XJL6jigHeU97D7ST/cuazlGinX/t7YZKktG6MeZHR9+VI03ZYAlXH0ejmQ/Z
hBvayqQuIuS3SUhu5zKN1gKVcLkXAi0FL8mfU65bwcOF0VU3C1kKPQsd2lFiRlxyXG3Yiw4XCrSu
Fnt3XH4Cxaf3X8QhUpAP7PyxLh9wouO6IpF9fqDECQG/oww2zeSominN/YSp8iTrGIqBJhv7HF5+
PRH8tD2qtH4c6Z5zrN73rq8WaSaPElwFw9qffOjsmiTgNGegKwp3PSbcjLnhdAIkHsnpaOdBom03
lRa4PZF94uZItRGaZv6MxCiNREqVxvP86D3vmcf0+oVPLTNLYgXt5hTX8KLms/OAwh2YaIhlNr39
iTuMAnjbnVSR+9lETbYR69S3sA3v2zjxtophWJkOXuHK+EaxZaAdUJNWImGV4QuZzMLBaKCIfUjz
zSEB0TInKUH2xuERLVaxMKM7k8xS1sRVKY631S9O3zWJdsfR5VVWrfottPYmcc5vVAknbSmRZdyg
s0f1hcrBvkn09lJO919LiWdRuFJcjo/gKhH9lJ4uTvsK98UbQX/yVnMngH/cpKmXROMVsNH0FEWZ
DXWg4BQXE94uQ+WSnlUhOByCvBudw9v+pWsEHIq2g5DAml/guBB4sIiDAzOqt4+SKVl+VeAcoMQ0
gxEdXw5RtsywzqDAPG7yl5GyMJ4/wgurNH67CAigCKPugmXcUu0sPT/2b58qqOnuaIBbv/sxFbtp
Fy/LimfiZggQUCk4CcwqL8Gh4LV0nkWxZrmiJnGI0V+JPG/+APkMIjJFpzD4qKDTHQj1A72AjMBJ
z/LZlrRWjudaABi/62cCvc/+iSe3pSdzWCl4C6TNZvb5/Bv5Acmiq7UpWaxBrlNxqRWDAgK5BK8g
rnKwqjpanGD8yvsVQ2mHn66G5dhZ8eVMDsBtFlrQYecXFSO0ORpL0tbRVJZLfx0JcLSNb/dDHGgV
2JuUfP7G54GZk8JRNnCwiDBPRuBVMq/jZ9NDJ+tozYtAKtEhgPPzrVH4uRFuYrgEBt3fMl5m/OR9
MhlclZV4/zvvGBtHHnOkEDc/vAZz9qrsb6FC4Q5XENq3B0EjCzzJVIZOpm7XG0HDPte2SFh8eUoS
+CEREJ6JCbDRjTdkM1FRaS5vbzo7KJwInlIxht2v5aiKtJEZUlWbENogYS7U4F9mtZ20e+5UCvS7
MIt/PanN8Qyql76JvUr4tnf7A8OuOw4ROVdALsUrArV0kCLzjHgi3HtWLe2AJnUIzNupaTmLYM6I
U4+PZbBot+EAeOdadGPbR/iQVAoNJ3cTpuCULIHBzv6SFgOpc6tR0Hqq6iEgi9dX5l6f0P56SLTt
7y6PMK6m1TT/Lq2F0cEvsMCWAVQcl+9c4hU+C723XP0Kc7xGGlt/LviXIxjsqIJKSKoJXPLHIZ7l
8APS/yYAgVe8biqdZj+6bQoEHlf08ypKMty1ZkhOQ6f0IiAbZEyRyilGj1zTVsCCkdSlLB1lCBe1
yY+rFSHgsQo7V05HsfwxrLXMxWRkHxP6JwqLqDF2ZCbdjQiIhjkGf5DanXsOVfeTv7Hx3THJkhOS
EMg15HLSW+E4Rp+pleJXcPc9WmX/4bTFwvdAadlTeJTyw1lNjkrFzVTXgzBZtUAJXTFSFeEgYJeH
zDf94Ia9elTjhm6XC37hS3JYxZq1fUIida67yicCGFcMthc27AP4M/4EFzpx1Q1tcSA5di9tGw3D
ckTaj59JMDNMNsPCP/7+5VJmxMiod57T3+foLbGIwozSqJZKiuFDVhlhHIxRPwFR2d+urZRR5PGA
b7yr4O5CsoEuOHBN8PBh+ydDmCLGWvb7sRtsZNCm8S4aL1nuSKMswdeYPe5JfZohRtUP5fWZaKpx
jHLkvecWE4l9s4dRVmv0bekH0WL2TXFE03TEmTShUBroB62qv98ggCbyu/gaK+jagsHZbVMV5WK3
zDRpdSaRQKa7fao+34YcmbwM6/UgPi3mR8ZiCVjCRc+cAMMViJcc3mt0BuAr9tYZqClFI38yMC0p
bauvCJChIRB3W4DOoTgEvhn8HlYbfQE5xgmGiTzxvWdnP8T039xF3+881I2fLdlG6BowqxrepxYX
op+7cTz95h11Bwg2F4BFL8MSccrL5FKKpBNiZhRdWwWjy1mi3VZJ8bRIZjjsuffhMApbw8IlMDx+
J99xILMh7LBvEbEDgHW8GhSrGyEm0wz7ZL8hiRTCskqHyRP7DiQE6t+dg5Gysoh7y2UTvIIjZps1
GAutPp3Fg7ivaRSm4xa50+zEfKWkoZMO5xu8rpApoUxqMgP0nePTseSTmEogo8RRXM0MQ9xqXCkW
ffKNlMn956z8rbLr/qogu8fUQv9Wk9XjjONS94zwxUjQhAkCPxDJS3XOTns8Pr8i82VZKGG6IXNu
yGmcwpbUqBE39kNYQfVzOAliLZTJlOPbomzHZCwmDLe2ZsN0GgZWmQv85v2EiaUpiYFPPwl1BeFw
4ZdDBCCnpZf2IuU6UkERwVq/jiOsKmjybGbG1Zi1/4krzMimUL4FE6nci7RfkBTgNrdy54w+PZ5h
zLn0Wo+HUwPm2a3hSoX+BjcSz4Cvch8Eir11aBgoY/CiPkDOGERqKLxulTuFDtXw8aHuU+Svmvqi
IZnL9ea3l0Os7YF5LylgMvgaUVMA/R/DNk1lwhAiShaeoqgTOZlvjeqPrdTuuZzp/LGXvZsmcrdi
qOwHI3wooZAYf2hwIKsuIV1PAJUsPAxx7FzYgBMbvN29t65zzxozbV283pYh1bEQPsRoVdrZ4kOc
/xDpc3sDowuQPBfF7VCyyWN1advOySL8/lSXmuzgFm6fxf7Sl55rZpz0m/GkNl5SFHl6otJ7IziI
evjgXllirhAwr+V74gZfD7Cw2x0eAQLCIrEJFnS9qvbpDfX/B9jolOhX36ZdA3byCprh/tzXgqUe
ACqLSFX+nF0C9ZTO7BmnWtv+6zkZlsHP1/iznuLDtgLSSYfaXmq7t5x23Nomtn9wCOikxqdU0mQt
sRGnwBPbLaokoCIHHOO/QnmRJ2yIjqewgsPDhpZ8xi5DcV8rHjxsv888RR6vIAPV0yWDSQKsODUG
VmfzBb0g5562dENWlL40hV+6HF8OZIxoD5oVimm3U8kX8lrvdQkhN33u+mpUSCU2dbqVzH+pGY2K
V2QRU5XqcOqfdH6IemvbZ8ISobOBa1DtjTomhJo+c6cYgJcGsGylulBn8pUZIOwLLTlY4N0QYv4F
VgoDB95EPCMhBEIJoPNIAZiAfl6TbA0UajjdtBYXLpQ7aP4v83K3r6/1Ecw36j8WrYGj6H82LL3a
HnjfN06n3Y4sXTvQsIHHusc4oAfDdnJyo0796UD9KV8dpiJX6GESMmzOOxs1Nk8rZgkNbI1+5+Z2
F8mD33Nh2rOhRuBdWVk2famjpandHAMK+WiBMjiaphgUnVOeWr06xq/0Hv/Zy5gXSCzu+ow/lEGt
HXWT0v64FUcjbG/Am6RAvwpk0u/Se2qzhtkZNlIO3fuM1BuEefLu0w1dxXi1NVre9/GwylL80VR9
yEU4IRsppjNc9QXY/iOZY/dhqmfnGpfq3041fnpkEnuVK4rU6fckbRvYoHZ8FyVBDhtcxh9Rnnmi
q7thTGczWnMMtZxFtdEyffrCuN2cYxVcu9+Af2gFjwODsj6VBRDQzAr17L9Ga3yvIFJaWt3smuum
C7x28SwPsCDQ7NsklLafr+4DsdFdyXFPaECRfvGdNvaDe0GNGJfCG7U1lJi9gR0h90xwPr4Nt6G4
5s8sa2YD8BWM0p3zgMJyeiNc6zgKe174/CiYn+4ZK5PKZJTspsErTVB07sIiOqVxZD/NZaF0EJ4z
+w8w0MpAeZ11jyz+3aDG6VWVE3vx+WUYsjt246rBAXTncDisFFmQGpcJpPrMQmlfDod+RDalE9VB
p0uheX/qOwUfJ6eEiMOgefbcb7HbuS9zvBCCF5rjkVH9/SdEpqjIb+2vuqySHDNVpwyjF6QK2Ypu
d4RGXHtu9wME5SsvyNxr2b4ofoITaYij/zyBZtVj8JTH6OnKrvWmZ2pea/V5WzwtkoVdGqk7Ydz6
3C0hSPCuFoMDD0CC2pDloKc5qDNE5+BAhi9neYqTzizRngUPl2C0qpz3PoPe9NsPWPc3C0fCfXqy
csoiMgxuWBLu+xCR0U1Wxno3spH2wcXcFzjsGoHuy/TqViFte3vTejQvOHeCCZaEfjz77J8lIi86
JFqv5gqz9Qm+Vjg0X1NsFagR+0NGmWZAroOzFtoYG7HbHcIiTYuQKVu/46n5tZDzYkbNAcy0W80i
TiIvJJAIGLW/yQuLyANpaVHfNoxqmV+dqahZNNccyvDiEi97mqBqwYNa8x7KEOd5VWld40zxX8dG
CR+LiVXc9jdlJH5exCveu7rIJgZptp/Ew6f6lkia+0clgIr0L6CqAHs7GjpXMeW2BE2o8qqq7Ads
tCG7JKL2eSgGLgAM1H8RL4fsu5kFRJLwSSONfcPI5LU8h0sSnShK+xHp0x6LaQJ5xAsYUa4jAYkS
kYs9aUDD9RnnSMcBC13I9kIbopCgY/d7qVWUFMZEZbxgCAJPxGO4I1k5wu0VdIfzOKMPN4Fpsnma
lVG83DYQ2NL+O6cV3d4OOoFnP+RdBme8X/AMGkUHH+7qFV194mDR6WMPv5Guu6HqtBwj9DGAxE1a
1+6gIMaWOug9YAPU6RyuHutrn2G7z3nuTmE969R4CC29Z0jsnGhlaMNWXh+HG3mGCN+6VFD1iY+2
QgeGkMXBEVzVOWn+I3KIgz4+zsJ0g+ZMAnhbqTCwuVJ2oO8TzL2DZdAwt223XZ0012i8SJ29zp68
s7QK7ly5cMTT8h/BjI0Q2fL+slCSVTJenbD4+gqRP9xAV7J3b+mgYQg5/za138Nq8Cu+YDODo+XI
fSh95UnUXD3mSO4qI2xbITwKk1qQd4sfhGlc8ZX5ji8m8WoRMJ2my9fpQ5LbbjPHS8H56D4WAxld
pi7UV2JDE7JQ49j2ejsJ7v8XviaK7xdgsL7BAGvmMrH4zFROgYFLdN/jRySvwhyHoQyE6WGa2n8z
gdeT+Ev5VqupKqAZXO3yDyDMMRSP/zh2MZlW41xZtklU7svPD+z8TUXq7VL6+mYn8IQAZj11gcEt
nnmwlpzbJ6sq8AACACkb2D5A3QCSXEWYCjf4Zb3pOvALIZgkfnTgfalLp68Qg2yNxw4I38Aawnqm
8OEHwvt0bgTX96qs9/17ZzmOKPP1iwovyzIWXzMkPI4NGtNGO11dSluMYSs+bzXSm0LEegCMN5nE
0+79lFjySonQ57IvVLv9Vi2Mn4zG2YR0rwpgGRBEZZ+aM1+CK8f2vEGefBMMNHiSaEdZByKrQYAi
KrRTV5Jc0sB0gwnZI7WqGfhdq9h5KwQGXWauNdP5WuPOHT6Kb8wO7Bc3ZmeGRuFXcSPDiUYf/u9W
aX7b/p0Ej4qJPbV5xF1/lNcMSrmmErb8/GBKKVtE7atY9X9D720fkp4tKY/VSw8XHO+S74FNiVl3
z17/VOBp36XO5TAUQuRmf2peiNYHO4DDKBTpd6/8F2DlXMCgM0Mx3QW8G+V7Bcxoaj4KWi7zkux2
0MyrZghwvlcVL8iKrtvH1tMojRMA/rD//6SF9xO4yVpixXL8oJ6mQNjlXih3b2PsSTgpxXZziCj1
eotglIjpKCkTdB+/m+Gyph6i5DO2PP+DyoefqNkBfX7W4NYuil3MJk75xa0POK7t3f1D67D1jJ3C
IcBqIGWL11hs1hnL+MWeDuzSibDFA3q3E1at3TpJKopkjPK8XcRZaz/PAUVpJrqD1L9y2DX9VZtG
w/hvpfbal69ssc2ac4Y8bz4M9imOtijMAM1QeCYMv0rL3mBqpwM/hEfMehey/uZgSgN8n+Vm9XMg
3pKsL2wi1x7OGXM+t8TDlTphl9oTONgxDKenad4yuxA9+3nftic3tvB+m5wn2708t6eripNp2QdS
OoeYrb8+yqqC3EQNvJWv1yKYfj9gJT8sqgbQVh2nRUYNW2ojTcgiikXR3aZcr1AafnhnrrZhq0T1
MrQItCK3hcSxoOE5nwcbyidFiYjEZTX5/R02epnqgZ14b8rRM7Qwxp+E9DTKZSfY1TDmuf+zt4uB
3JkRzewLm4yP6o/2JrmToBSl07snmFn9YJbCT3WLNiogVn8rWaZmO1SHJFEjsjkZ1xbwZ025gAEh
b7slcKElILvvlbKlv2uC7tVuUR6iZGGGOoHVf8/2/U0QwQ/LymQ5xYGcCK8DzPjZJrEFeMd1bEd0
Y1BaD+q1Q8HkHKHh5Xi1mghTcmrYaERG8Gpzyk+8Tngb6cWBkNkb00q9J0u/QrBqvHMpo40gX503
k0T/fesihlYG7Ba8s7SeLuecDhynAyjsdCjnlO7P56eOubanvwhHzUzS501D3cAIKFeDmT/ameGw
pMytiMGiGKw9NgZ7qz0kUtX0T2u9fEqHz18uGjfq8YfXDjwNTfyWiUre9CQlaySx2LKWY39uVwb/
GB4p779EldkbOb6/T1n6rVLwfVt1Q9kMRjVJANER3mbajRCtbFyWxISadbl//g1hRWlBfjCDB9J5
ExuB3VRovk5XW1/Ls4j9akG6Iz0EAiIXdGd8XG3AJYp7WgmtE7PZgEpTxBgVDTHBA8yfeQKc2NNz
Vz5LJeWbWft/ECY1euigG1RiPPKKG5KJxbPQNgOwxztm1yT9UVQNkwI62stIo7eL0+EYToCcuRfy
WHF+l5bhz33BB+sL4m2tpPv2HFZzjfGxGD3QOuCDmldr+OjUpaH6fW0okEKaIOii6V3jRnfD+tzX
fe4OfBwcc+kTRhBrtcaZ0QjKXZv8RSCZehsIi4ZVcqjTCpuRwEkqCLIaucZ7NVa53aLAmGqlGPwx
a8oZiNLFRfjxF1mHcXnRrEjwwTZVRZyXrymJuwkN9HRQJnQYaUCOQxZR01kN3MiQ8Pz1DjtgNd97
aaVaz8Ce0X+a8XtPj+REAnAswQGa6afSIk9uP5tFchYKuO/YWHmlLScWdZSbwM+u8Huv1D7MvbLw
eSSNkObkiOgChr0If51iGIEGEEb0CcppRSkAoOjaz5PjKCQ9pfzAhE9jv388tq/xz1b5//D92/CN
TxK/LkBsSauYP4Ct3nChUZM7cXSUOVxX98xZJ3/p45OMl3NZXuq7wBnRjpyZIfoPL1WaKXDCSrNW
E76Uk57u2jsPRybOgbMFPQrHq7peEGIiKXZbp7ze9dy2CTQiqiAISETMzhAEmmBJRZzbvbSj6FMD
KzgILAK0kTxLn9YAwUU4AUo9b7JeXTc2xCpS8iCi3bddbFS8bR4qA9rSJ5TnXnsJmkQ/GcpQNjje
aKxiejVxcrPtlqygE31p9t2SFRb4Iwr4Sr5o2Pe7MFFHIaWvSATHRx5HPm/bdinspYrvMovfD4DG
m5B+BywOtLXd3ua9NmATh1WzazBB6Sg94ABGifkFJuYMNKwUTjZbn4VCkggyPajHQJV0rUR/Sfya
s2P8nLD/NxTCYta4QhFlp3M4cD2oC5MQ4M0fYhrPHMN8v0DHYQT8g0qfIhlENQPOET55sfEfCH5i
an96EFP9N20tTxXwVFboiApBeV4y4PIMlihHjSnJtDAp5J1TBYKOEgQBLtfeRFtFcfUhG3C9tcha
Isslg5iKCUqcWzjogQpKyQ8cdS8A7ID5ZCBGNr6cwXpLX3zY6+hYBgFIsUO5ytzdYkoNaRlZNdqI
f9qsCeQVKfEc71NYNkHf9ZIh6MahNQsgE21A8DulxcKYfDoQ/ze2KaFN18sWq4Bn2Lj4DKv7VQ97
t7IDw46LPL/aY0BUHHONr20oKhANyFdRmmiyIYnjiq4ODvpFnpvFvCJLKqLZmUOwfoB/6dhdFGiR
TycQDfrxORAYJGL90flwjLQr8Fl0j0l2SUQoI+iiOT+SFaxE6X7ZUj2xC5Xdnr8icPeE04Li7OIn
FMi0xFA9+nvZUFreUUUXiODLAQDnDPDV9ooXZf+pfkFPZ+cIoNSNckWw2cTVik+Zy/gdF1Vs0ZLC
DBZAq5aU7D6VoI+pNSm1tbQdWOh13uMYeZlIB4+Cjl2CAP7PIZ0demm5AtiC2lT//Cu4o8li8smW
rsKC9xlmUhVmH654JLzAKLiV7Ms44n32x6YDInQdQqbNou0V333tB9gxpqHJAHeFAj+E62Nml/7g
YlCwYckc+QqrCucqKU7e1T2e8hbmwmYWaJXIvIMzeyb2VUXjN3NPKg2G11Pmbrqqa/VUksdR+MRm
+m8HyXfoFpRowy6wZKd/kylHmByQRKpAyuQGmkxhrC9FB3HdyReR9P9mZ3ruf7SD3GhyBh0P9VpE
vEOZfLALPVvXusD2J1l/XYk+uCIZaa7IjXlMaAoiXjnZVjxa1jXKFH7Ww1DedtfioR6P35LpyWhs
L8LpeQHmEbVz8roK6zlRXWx29h755p+mkyKMkOMiTuHexFoBApG40NDlL5QIMpQcbn+Fa8RAzRTm
XZmtYtdDJ88Zf0FWQJ5+0SIWzSY66oEA+alGZzUl2vV/jhqVCaa4Q5u9HtIS9XF0mCNwNo7UQnRR
hFy4t3nKZ+Wbu/1v7dTN3tnnxUsFf4DdARgi80obOk5/2iQXw6cS84HQKxZ4CxTVS93MAZWJg87y
3yWmhEReI+EXp6Nm3AD5JiTpfUhy7I/s3NU6jNxYhcoMnYsTESKK8bhWOKC7KkQ7g6sumIAj30zM
dQLb/JucMC5Qzv8WKh0PR1LEJYk3XNFfheQbQfrlGkbYpVrRNRi37DHOe8soa7Dd7fYXYqNaZ2MU
7FltsnQlgatuChQXHlTew4eZUhbBSIPJ+5bg5eiq2Uarwu85LS+uMH0fwYkdxCJmuUYlKnxwMqXS
zbSOna2cH3DNYWTqGwkqPwlnmkTWGPcu+q07YKLcyOcvu4GoP7O6wIFUE3N5X0SYW8e20z5dA8m6
SWYQu0PHpAu/qoOwUrcS1rqWOKUWp2GMpJV5NX8htDgDD2pmQKaINlCVXzCZftuDzvr6vqlqrj6b
497F3i3cf3RS8x0tZE1HiorBdxHvfPyvF/K0aiB3rMxWQKdDOioMvTSGdJj1rIaIgQSB6scBKd2m
yN9OtBo2QK/+GXaVOlnS2AVCUdqDrlN5SWzm44Q2HRoc9TDbULERDcRmtmprEE+j7C6frelijALj
NiuZN+sBOq5mhGMNluER4d29vaVkcxDsh3APfi1XHMVLSlsbibJwVtEKit9YOI3doccYHFy4KSYl
fxkCYWKQZE2lsf1j+W9yJxeiJEYyIEkTE+IXJEW1447StKCcO03w0h61eHRJ/FnimPHcdGHxHewD
UJyM2PPc7bZ4CzNOmd2+1YPNBh2D9VaNDivJTFAtEHOP7Ue0GgVI94VEg2hwcZnut4+hemSmacr6
4cdGcufKwOPtOAiFvt4/pp4Qe0RA5PhU9SfUpkqpJBOuLqYLGMVgv62ZPrBOWiybg32QaU538Vrt
bWb3gkITK0FoU1+hybHCZ2pei1ApkdP7bbbcGd5jelHF1ZV5SoF4rdJ0d0ZB1ezXRF2Szqf7JB7D
vOVJXzwdGDIDhwZ9Ful1Z+JW0rqGIfeLnO5a1nrx3bwfjvCDXvXdotNNFHuH2o6Ik1afYTiP45Xz
yIUzo/2uAANHPgGOsWrSQDOvENCHtP0oz5MmoBgxIRuYSKeKIlF7NechOonF5WhZFdme9LLIjrk/
Ib1R1tVQKpw0i7HNtwjEsXK1F53oYUzyj+nrZmjbZLwtiy5daNF4u5QimuiPKmVE33HkscWgJ6OW
KxwjyRPwoDwcdKckfeJcfclgmcq0/AfMMg3LwyL094ecUwwX8AqbmPulqftaNyQ+OA6vM26jYM3U
wVDsIV79psa8j+5Z6FHvOeFaDYD+vz3vqKQkE9VPnejVA0BuMnQwHQfVaRm269qyca6uQ2sQPb3U
fOargQIBSbx4zG1DxOqN2fz2IgWsWtGKFWbyJAvTFDiLfYpwu/R3/08aX5+f6nn9ePV+aHThQOe1
lN2esGTc2Q02eX6FLbfUl1T6whRpuY09mVfjv5gjri4P4Ld/5QjpDx+IYs8lTJgxLQyyVY/GwXxx
WfCu4CfyD38Wl6qHbU9YIa+zXKisrRY44ZuG83FRu9QUs7V1wRZBSAwo+WRFw+eiVd2fW2Ty+YnN
a28ACzBO7PTjI0ionJTVzx5FpujH3CPjvBpneHx+bC1/2oJx+VgFPXQfADCkantII2RSPqrH6KZU
yNmJiF9PFfHbf/2tkYJf4IUPfZcGDV33byYNSaEWS3i+oiuQNB+fgVGuyoBGZBWAedRPTLc0yan5
81JmYE0CdXQsxaIR2dAKUGPSz3DBMbcvY70gxrKEMhTVY0aWm3d/eG89IeecfBWx5DfAHxkKF3r9
WOPkias/s9f7646qhHKnQO+gvMDICpDHEgy4LyEdy876XVvhGy9QqvrX+ZJ6NK4kKYWGAoJOuQSU
zD8BxGKg1BnIWd+l+/BZmLX9GpqutoVQlm66kPzFtHOpGCaqoLdQQAd2ibfZmxUjO+66ovSj8RzR
bLtv9dILP+5g7GG8FLYbdciVf6Rv4awKAbivef+RGAKhfx+bz0t8IdNXm3qA9eJt0Q/GBuErGqQx
XrsI4+mMuFj8JPVjHJkZt6z8Qqs4mYgSEmdF4PFLQcIU4ySwWfgxpXIbPuWLxezLQZ4aTvxE7juI
eLs/i/MqIe8O15NE3v6L5XC61aR/WqrGxrPrt8iAZUv9dhKf8F2xF9ZQyvIHseXu9c8aK/g3xSen
opGGD7/YuH5aN7McNJKOms/MJJvQzi9fw/d3jYXv2fwKZOo0FoapI97Hg7OuZtLLOyw36JhkYJJF
pDBURpcJICz4vRBUsntXo84KdsS3q8+/6lMrWS8RnS3UKJSQKwX+EDSnRbwDtN8dfgL6ZSUQxFES
29QXBbI74NplVql1vdU7ykhzeZa2bLrfcbn3/DgON5bqAmfZc1vLZ2qMZGpB6M3MEBQwXjSYREpB
/NXWNR7hEopH4C8k0nHnqBSbDxJM4hgsYF6VZCmpa3k+JXPZ+6fsOnqHUIrEAIERNuUSylaNCnMU
3+1XZLd2XpN3SIJ/YLI42l6wQ6An1b6jn19r6bnggfTC5UkycMD7OVhJ35+4H9cmiErNeLOTeeHD
WmoF/zlLqf4w22Mgo1/K8bsD2LOuCQoXmoKSbfZAtHdX+MhJLXusFksXYg+wI6gkY4lymi7e7pxE
zjrfU8GHBtshumBTQXAxs6KLdMqc9DFFnptYyKOqOhM8h1+jKthlUxiC/LvqsJYqFFOZmxOeil0K
zmW5JB7hZ7XdRAU2suyfHJhf3j5A5AiBEX5Orjf/nb4M4AVGofc/KGd/APn6JlTWWBGMF8C29S8S
WFmgRUaZLnjkasREriQd3y8jd6zvybgla6CW4Ylkrl0UH2Kb+TqCUvY3jb0lywVIHFA1TDJahokh
gV/4ISatpmEnnS01EWZp2aJUVe3eDaTclr/DuBJMacjaN9dxS0yhHOlDuUZ+SbL5tIs25i7DdJk9
/cfN+bGISnw6Uv8yibSBGxbmaRn1mB2yOID8dxdkYNFvxCaWNVuupEeFkaWxP7rVjETFdHAWu14f
jaEHt2VcUj587+27xfW7FIDeZVoqh1cDnImM+UJp7P/2VQRWTUX8snJO+BxKoXHyc/AUqfRM/fkP
cJuUWqMlX7bCGp03aw7slfce50P1aaZZZlppTQffmOaN8aTFJKq98fp7ONvgIYWMB910OcfmbzBm
geVKA1Ffw8MStwLmTamxgMj/AEdfWL2FlPaGQYM0CeY9hk2M825WyoNVPHKzA7SvswAfHQJdpcXF
lnjzaCzt1cPvhGzTvNSpFAZwB2cLt7O4n7dsl8jhWrylxudXKfCPYL27+3WctXZdKRh40oUBuKNC
sqUuyMpuDpPjJFzFMcullJCRRXAlq6i8KzP4RpMM0LFSZbfeJsN4k7lhfAF2AewQkLgfbGLx2k4W
rMgv+zkat43QHsaNpXDnKE9b0g+H806ljhyOTxrcNLfDb3/kppg5rwQhTDozgEx4B+NYfWRnkjBJ
gYrh/5xKyFNHWxeHsfmhR4Uve/lRHHIkylVqPaXyb1HFDcpVyvUx7PJllTjLMEETHJXJBoSroRat
sLdFrDPbCKI/UwDDr0NcK6HiLKPoWWtHbvDGX7BiXUuhk4MQt5muduXSlLKZZHAshszFf+IGKxpv
lGk+VZpY2bOWXeAnMH9fs70sSzKurZsSeKRAkg1EzpgH4ZKMHu7kbEqMYGHhA/vJ52XJXJ0Q+lZH
l//m8yd7WpxoKe7mxs3szPJcoVtGCxThkoBWaAxnzH9zGt2yYESbksHYx6fmTafUyqB8VVK8ecm6
PUdbttkyg5MtaPFPBc93tBV53deVbE93btMjYpGtVRUJGztUSZkaMqd/zovKCuJN1mtrzIPYyDDA
7D2Hah/S2MbsznW6dGsU16fZaySWEIIuYXSg2mkKgWwliRDQQjILLzoqHdlBOWiiCaWnMcgH38lV
YRtMaG9UJUhc4gOby+w277zbBfwd8npUifNQDGk5FpKy4EzdyXadsK5rXPsQUbB00AAt/J/7ByzG
TP9sOVASrS3Ojrqm6k7RGgQREW06NOiV99xMvobbEVURM+0fQjjimFU4w6JiwbV9QmUJ2DV22zK3
1iS/S0PZUzfy5aq/VrQ2FxIcvSei9mlxrKCOOck3YjKO7KmQrwupuAG77JIX32S41U64ctIvWGDz
ENhSSBSaweVhxHHLInuQdSQi0JTV3eA/kIMDZuypYjyJTiIWkkO7qB8HcsDm8T0wGGQsI+xBCi2Q
4OCNbvtzVSEG2oLTCLbanuX3fyJpgFCxQSo+4Pct/u/9aQe/N/llLDN4FFdZaV6q3asmNuoSQ18U
zVWDLzwWFX8Z+gnLayRKG8SuQ/W0lUcA+ry13feAShaqE8Iyvnaldyf/qALp4ZMu3ASXBawVdAiF
IZEC1BttO4SdwJO/0V9aSJYENChnbMbv4f7058P29ArWplohzlmLvnufwOrvzpW3bLInt+H8b+uX
dpH/Ug61XScvLapENQsAkuWEJlt8e26EC8dfMIz9Wq9qMH4txkgX4pOf4EGe9SoD7xqVpN1eml73
Etl5XpNZmoU0EPBVL+Leb5+/BVomV3DOog+EU+9e7VdXzVZ0+WJWB4p1dJ4cUlhfTHwIRDi/j97t
YIYu9szqVtQIAKkex6VMCJ4nr4U9WrUgbYtT80LKl84ZPHbKiTg+1Ib9zVOAr8XnsA+dXOFjwudh
7kdbqxleiThbCxTXtZo63WyCtPZMtM0dsWDoJ++6MOpmjsf/C0+upZhYtVKSh3mqIFosZjs9u1hV
VDLyK77k7vCm9bCGgMPTJhRowZSZfUVPVlYEsD0D5cH/yd5r00UeZF0TKTVroWbp74ZP9KcaJfPp
hSp45bvbMi1db61cL8yHRRg23ZVgpdFAvi2IdjB1mb54xngiLKb5v4eoMiU/tLISwW6lcJgemXJz
eX/dCHiC18XZDmYBaO1yqKWxR0hANcRD5byaMOIO3k3E5oVP7SGHdDckZe6GLwJ287b39IYOjNrU
rQKJsmJvJJD0aAMbt9/ElX/97v4vGOkVaaJvutZ/WkV1bHaQelTYpFCEjkom1plH4sjfg+ifztyN
KFPgE0nAXT7RRr3PjNyHXgNG3zmVFJV7qA7zMG0P6SyCFHtdusSoMlEk0Vb4KbwWkOzS2xkVx0CB
fMu06DA/f6/6s25JNvOT0TW62bhATkZARFU4V7gDXWxA2kT4GaPKGApkyZh1I7tO/7ghgUnTaR1j
u7XDqo5R5Fln+5lMrJWyJJeqsw79+tgLaPO5Pn1XxB8XAcAYw+uQ5Bb0MoigNAVhNkGBf12OrWBj
JSyxsA334Z5MkONNNnXJiLpFjKQnSYc6lyz2vi/xc71gmAu3kLsTxPBWTsVNgf2537WYzmuYFMox
mYbZcq1m7e8Vsz5Y+Ra4XqsuJ7RntpIww7WfvC3gmShbHIFPKjSF4IYPBMzIJgWPtDBVmoSHSzaO
IFv3An5XoeGu8twvHoJNzIpwJ4In7OOPbyJwByjy3z5IIdYq0BnDJ2ImPY+DCMP4J1BLjGqz8sWt
I4PRZu6OjRoj3m2Y02R3qa+QUwGMtwkMVQC0LYRX6T75qVdr+PNUTne+nr4Yu1HQpsfzE4jl5OKv
RHf8u4lD4nczrO5444r7cZn/8ZydTGcuNP5RLzwpPTcTcGduhJznQ52dzGXhG6CVXTR/Y8wUxdbI
bUgf1rYVL+xT/95wOvAOq6dtoYwxq3YraNPu0oGxaKEy4mL20QT/hWGP7yIayWoBKoPhfNpGc1rC
ZAV8nIcFfx/HgQI19YdtNH14KFcnm7/723XIQBShZG24bMiRggHRouNGtE8dZ02w9KIh9F7FixeR
NAD93eXKpUSYFNr+EAxGhZBhL9mm9MS+skVFgcJrjdkQ9jf0kUrW6/7AjlriBhivtHm8laqjxbds
l+AHnKfm0Fi874dFaEytbJJui4nVfejzqY2lbUv6meExhbqXbbIIgXZekGvvW214uHRxNer5c/SX
ItW20cnrjMJNY7xx3cF4dZ0ocH41pK54PZ5FaiSl+XpBk0LQBiW00HJena4W4B+5mXdyzbm18C7B
ta7LagdT7aBvJvQF6Eb1ye+a5F+uttX69hcYMPsf2g+ymfw/nV/GiwQmaHKvfgg66uSpM6a/Zw9X
kkmhqw9Ljyka/+RUSqbAdkmcCSWdY6yF4UCVQHV4BaK1h8T9+wsIIaBSNvQCrUyrz3GRS6FeSOEY
Pi+DC4KuSTl74obXbO9V/KYlL0bH3gfHDJjZ2wKIAonrnFWVfEnDUjmpxYzXr8TAA2Dxq2kqgBCP
9z1bVEO8D4ikpEXQqEilTvtRvQZE7VS6rfEAZ0bPcYpoU/yWZBZc7ytjus1Jr+zaa6OjFTJsRvL6
un07bnhL+Px0zPCE+l3y2povfL2diLTx8E1CJVhmCVkcHz1diB60YMzQlVlTScD4WU1uZWFy6pVh
CeR37zeDaimmaO29NMiydZWtpjSTK7teeC2ranWO8vFb+URosrKy118ZEsgczmFbuY9U9SEldWFo
owbRoH4EuYYW7FzpYQiABrAYQTDeV1b7YdDtWThtKoi21dPnVkLm8/5IVGersL2FtNi741QwBtXf
NLrwzv1RmC0AewiKTHof2wNH9t7C/7SmjuFiFLtKLA4f78PuN2JPCs4doYit/WgV3QdIdGmRVQ9W
ObE/vYT5ttlS1r2VWH2QJKGHd1N3c02N+IbEyTMOiLYLTsK1Afr09xswxG5UFvsFm6dJNi1oikUg
ibEVbzTwPWi8oKMfaU0JoopZLZrBavZXoQIhfXCOTZjTnfwcdEOMwGo3Qmon9/w0LygBpfQhirIv
w8hr5ZWc+jHC3D4YUED6E9W/q1OOiYJ2sIZozjrWLzXlFEsUjUQ5KvV2F3eZxcPfl0CIBCWH93Ob
J8Q8owBqwzNFlzzU7edVM0V6NJbp548U6u2Z3XFZpwIbOCoU/HOzUAVJ7dbbCSkjsaf3IUsYXFeg
t4R5i5v0cJkcSPSTGChZ2RLKBCrxie0l6oLhmj40eDu7LcoxyFXZH1u5CRuWRyh6vBOQ9+yIhBVa
dC5hWPMMSQRxuE/Pj3a+eoK3HujRe0F820hYhraKCGNUAZNY7mUC93mIlJWAaqbgBzg0e7r7v6Cn
HEHk+I9RGb7Ts7mnKQ7zCp6PCzYTmrx3tiK+e0CbY/LBQMWlhV60veCmlmUeAYQ9sg/9AMToVs2u
Gi2W56WOKoYLoeyN6G24x/PPyFJYzbyCf6WA+g0UIK8y7lvkLAdGoDaISOAbVVjNeNB9cIlyWJCI
61rfKFmXRNk4ALhVp4kC7NVefdAfrEBhjNsCxK1tzyKzUT9wcdBRNifulSr4kQrCxRStKut5AGS2
VnMtswOwOSnbkeKBWSr/svFQ4LJwCtm1bgwSGn9uIyEXIjW+Mt59GHpFkRhRCz9DjpX059kzz/TA
da+bjR3MsY8ahhRK076sFzsOAbjKLbTiVmWl2HvCl4a3gDY4NR+f2K8t3jY7RZe+GNibtUszirIV
5Iv8RFy/HkytHigdBpT7GXmhJPBkqum12K+K3rPUXqMWZ0TQPp+OlHaqdgx5N2JAE2yJVKW2uGsK
jw3Gow122nv9Mfpsbn3DRS+63gRv+c0o0lQuE2n/sI4PmLVosTYPMAXiB7er888qvGqpHWLD5z+S
tg/TSyBtdXcohzBp2emtj3qjTar6O1Kx3JuS51PFuNlnuybu9EfqAZdv7t/7V/5YXy/S+lKCsB8h
Z+2WEk403HiCjn1HJI7VzJxWBLpcS9iJU3xwMvxd27oGY03JcRqqzB5OpQfE85vZI9L2V/mLGCRN
Fje9BTbnxNU4eDRph2EGCwGSaubNXLtp9nXqONHg3/+IJpqBoq1g8OTa4bAgdjWstiPLKJJHA8hB
LHjxT0eP6CJi/Q6gbfmb0VqjRJhQ7cB6D/3sb5RNkUIH3ax9N78vCXYT3OpEITRZrZdUVxXk7wpH
XSJ6e5+OVy8lvq2uhJDJd1sf6Xa7XlBG+lFJEF89RdPYwlSUA/7CWZMYWLQhDV6Gr6sTqCFsu6ho
ml6GNE1P9v27R+HMty4OB07ua1ZgezmUCXrVi5tyF5zFqHVW6P35bDixc5y5INEwKBvnI9jzE1Z/
/j2Vi2jAz8hWfCFNyd8wVdYz/ukxu4TR2O+u23dwOCci97zhR+qqyCG0k/qYQFoTbSTJAUYRcKuT
Zdsg01qDhVnbCuEP3dANnnMhQ8Y2MetXfH2WetFPmrwYvFAO5pWSjKmYvzRo9mdc5xc6PIzMPcOB
h+T17fOQH5QCqalQsCy3Nx9VK7wUixRkBi9WwaAHhKp/2arN+vTq+xMiBEbuPror2OxkaHiwWxJ9
0Cl7aEM4/n3fmjDBnhBTN8AdNjqWRQP/K13t8UhKpcaoGWHgpPXUgoRgUIeJNRw/cLpmOqzqbVkB
YC2hv4mv2H7Tn1/c8AJQEdXPrpEpTkfDBopXKPVDFC0PDKdT72LcoKuNGsgUnH9AS+kF/3MHk/wh
yX09zNxtvNU3V4d8llAK9cCmmLo8QtkrxmE8HdDx+HplyQyAv0CZUfD4kNM90FPwTt1u9wFRG8iR
JA0MuqrCo7dJ85Sysz4zFXdqwa7t4yqsOeJd4aqpIMmSurU1Czjeu6EB8not1UHz3JvEUlIgdmX4
7M3kKm/McMLgN3SBwJ6Agu8Ly+k8jLUmHCZElzWjmoh9QwrLQ2VbYxIfz0gagbRXyOqgD+U1wYVO
q1pmGFs+YmB1ebmJ1egc2A7VaP9i3dSjvrqVeVPz00KZB+N2p81rkipWD8RzmzyVx30yaOVmeLrh
aCQVceoDxEfTziD723HkEOhMUhbD7qmWjvCj3XhH66s3pBC8lvk6mAM5Ey+e+S4ndHqQadofRreW
OiAxfZZHXsUaz94pDNPNPq96X+qcM1FGNFSlVoPTFbEKB3UOw1DsjlAnTq542E+1hJ75wzZbPFKk
tG7wi3ap6bTdb7cr24LJrL9+iUOj3xE2E/eT6KZ6PLrN9fcJROiYyk2gVFgEI3jzI3TzIfi4uSFM
mnQtKoGXpA255wbpKzkFeRxwkkHCFArBUpGN3KJIJ4a7LbzVde+s1519WfQBN6PSPEjl5QBzCPlr
sFMXONg/r8WSh4Gm8PWexgzXz9hlq71tJNF3EaBXIBEN27pWjoA3AegbhEMYAa42D12ZQ11vABIr
BZZ7ROR5GBpO2PwdoTZaABfkobk8f39GggwS94qAaQhm5koyGuCQNV48Chy2tggdxND4F62FwgEb
46m/4Xryb9nhrTzVR6ebKAjXMYjVXt6ADoSOrSPWt1qoZTuBUk+7e3kxxgOIrkBIfAO0NxtYw7F6
RkyAXoMh/0n8URJrj3GVe+Jx9/ZLJX/zZluF/MN47r8jhKegzyuK8+aoJX7Qd5h4gCXGnPMjw8o5
gPTHnH1pj8CTP60H4d5ghvkyzIYoI8nP+3qoJCzgxr4Oe7/2OhgR0CgmHkD/JbcHCGOqbclpUhae
vhni/7aCMp2PLsEh5N9ELG/7sMGKHSGU9Hr42mKm21RTQBJgXZ1GZYAJLUIMXRS2QxfKq4r9CqVq
A+q/B08TJfsWtsA+6DVK4X5wl29r2uZR2A4nI+oBa5spM21vJA9MoUoVjwyXB47/xJXMtIxEhsdF
DPx0qNfAxTTexDcLS3/gVFqZGFwljCreTtc9bOmOz74+5begy1/k8E0iOrjjY364i4wH5xAsRzay
D1M8aOJemNTswcgSbk16NAyOY076+V4x7/3CHv+CZhEZu5ODSxqejETMedYIQQSCmWEgbQvQZa5c
fNbVPDbULsv0N4ltU5BUP2apc5RdzqNSBHw6/A0r9+ZBbfmQF0gdcQM3vhfO9vh3QvXmmIzomL1v
G6IrbmixaJac1pqXqzxJcW2XbIFfjLQO9DhTTdiQYCX0tjPsF+i5e6WeIUmrwhl2kvSRYfNx9smf
DpV9L/AFSX5/RJsiUN0xHcSxUY3ifw2zd1Xt4yonT74aLrQMiQpijM7cCjkZ8myqALRNoyXNdGc5
ZGKVqMFB7lK7EvZZI3noK1Zq2NCQglI1wEmi4aHlBmKuDc56yJexqkBhGHjfqBqughk14cp1Gxp4
xpGTrmIwRoZzAoftBijCKJ9V1EwULZAx4mvmcz9Jvx79q/KwZ9LIaOXlhJtv6mVo4Bibb2UOqrRp
1qv/X2QA3lPR8qtQcmsNwkhHqoIKcD7Hftq3eKyn9DOB9JBtafccFBNHEn4+hi0o5cnuGOkE0RqB
qvadhHAqWBZbjd/+c8Ck8AfKrjlOJ5f3WcKMo3nnG81eV96JGN8cCyWGQlah5mcV3di1aBoVIaia
nRe8Q855cv5H+yoLSq8M4wg6fagxJJ3WTzo1IddeM4DsQeeMu3DOO4nU6DTl3kbvxZ2bMUpALLYy
bnBRNbDiZGPLv8MF22G3X1geDW8SjDsCriKEx3WilVYfT/NrU4o7x1z5qhSgGTz3hYwZvtJahGJW
gFKbGxpe+a9Xqdc84Mqhe2IClZWN8J9RCLAfZOAJPq0befkZ7lycc4guAt8gG2tdq1M2s1TY3Bxv
KaQF2QOZtZXz9+y5ls1iqbpBFEINeObsviKlg7LLC04IYx9Y6DdUbdGzrgHHzsk0oHiTiU51be+n
pe7BpKPQ3SpIHAcyzx00vXQpHQCWdcugnrt5PJf4n/Lzn/CngO9PXsHNP85KUzANFq4MUUHdFHlF
OHHH8r6OHg+5gZBp4+C4Prz/ITmB5sLai/s3moKmHcr7RFVOyhMsYsQTacn8psKZUzFHUcHDatQ2
+z61IWgKCC8yj5ikPLmDMOD2WLE7MmzWk8V21Iupr/jMoOcJ9WK9rf16vJhYEM2zzYXrCKkwy3oQ
ID/iGS+TKCIYRwSyRurhi/XSyfLB3LY10TPzjARPlydLl64uXVAJuWk//cI9vNT8uDVwTNdPgC7J
MLVz/O8T9BzSFoInJ56/q7hIayK1bXwtzXhL9NPHQQTzdvAHnamW9yGjR6GH8ww5GlGJQ5kPfhHR
tIR3EP8weCxxSTKP+pifXZYTw7dWd/jdS+MRG/V1nbB0zjFR1fyLPahGDC04TY2p/0i2WANyQ1Bn
qs80jN98is9xLhBAeFy+qWE61QUhz7zlr53IkzZ9tq5IsvkkbJzuXZ+msWdfSkpEh0kKqaZEs2Ex
8eSUu1oftM94Gl2yzlCAd05dnM7ADWaAsmiKyHRJNfmijj6s1MBIQxCHbfpdpmvMx1O/2tKi0Mib
+LVS/Wkn3p7DOlWWDi5x1e1OVU7iiqzkx+/9Zs3zK200RmujRCJ1GkL38zCeZ+Q3BaziFmghWwGI
tW9ZzsavLsfuixeaC7rtRtG/e93/v1u4+ViOa3OTKK8UvsEnsfBmpveBMbS5vFvPg18+tLcJPIqy
yeqCpPdllgHx2xam6byWHurFHZzgve4Ub3jHDfYcMgbWj3MW0fWaVJaY37Mfpcb02LlTPUDQ5hXL
tGFI9FU/FHleTQ/0oTWxceMLNK/t0sIO8LelACBvEbHsizj6ej27/Kw/YJWhtURV/yy8HkpiHdsN
5SDJH/WdZ7fcQrHW0m14pryyNqoKnfoZgYb3oh7LIuFn3xVySLu/wCPC3cRcbZ5SE46drtG19ifP
c0VApMIrA1a0bXLcLHo4mP9hILMuote7mqPf1nTvh7M3YB2gC+ZJeO+tks6ax14cEmw0Kfd3JYPu
srV0cBhGGl+H08ZMxyZvzBRbVnmMtkVZae8b1AYZZFMzsiHPg7T+/k5rFhbSCVrwC9wEPYUhIQnR
QGnYZzYUpuvUYrc1uwwzD76JQaq0ws4rh9vfXVx2W9QROodjMupmEpDFjJv98z2r29ZA3z7QxACp
VftdOAFluOpHaok2WJ7DWUl2Gx2QyNkkMrELxqpxPQXpgNSPUDHMv2ntz9i9fdFRzLEnqgkK0n1B
7MiDVAKZARh6UGvXapplQ87Zoi2lOaptED1BS4eayAxAvRJtdWXr+DtCiFVNRpz1rD2ZBdT5M1Ri
XypKpn6OONn4q1MV6KXC9c3LhbdhukX4oiwlqjpG6cdU19ViJmFSDAZnCro6G5hNOPeghRIBfcNO
ujBk6mmpKhFEtLnup3qwbb6EuKtIALymAIw9cRejWYP8f04ykiCOrgP2SzhGCYtQ+M+fwG27680K
J3F6s04tVfvxOkR36OHTLMF8JOnLgW25UQ96aN1fP6KBSwp1Xu9Cj0GDDft9B2CfSP5bUBfkxQZe
3C3dm7Ioi7NuuSQodpTMEcsCjxmb9kT5+UMV3S13mKSCVW8OC15qNcrFmDn41zNq2exDnNNzl34g
QCCArW7WN4JnQnxlKYhxC4eg/RiBVs7CVMnVnDVvkFUogizf2jwNi1vHenJmY6GyRSFCY128Xd/r
nwYbFWEOqOXlW4MZgWha4h8eQxEhJNs3t+ll0QgceIURozH0pOJMrxTIpHOV6PDGTBrvrqPVTIf+
aRC/re82fYFmnXGjLgn1cgo6KVuUO4MmeCef1HeezWnbii2rRXj8srrZgieKE8OuMdt6ebaQSkJ4
3mnUQmUuHIcsIDDUkI+mBpwMjXEoIXepDL3dgHB6Q7b80P9veoJdxU4Mrxv9TY9V2DLhn0KytyoO
ofSK5P0xmD1KSn0jftPDbVFMtTrf9JTBGmMZUluQFVx5LjvL0xDkd5b1EL18njWD2wfBYVN5ZhFB
zrmX9xPla3nN7Z4/yO8NB/TBehFQa3ygK94YY5PXxaRp9TWxHvX7WTUUd+0fJ/Yd23LWyApxO9NA
b8iMjwItqjayoKxSsWKWcjt5+adTryAVVewXKSNIKsIOTnhYCV8pYeDNDs+gE9dau7t+RUfqhgAN
CZKInhr4qvfu1PHG7NdaKhXrW8G++4XfSC0afPG9idBO/s/9apvBxhF5PjJlEObHXTHUfegZhfNv
Qiw/6FDasfdR8KnvfotWwkLeJLdmWpu+4JuP0q1osdWJnVMRbMKNS7DN5NMFGWp0xqVp2oSfMIh2
blklo74mD4KERoQsmzSzKBqkCbyC4GtY1H/l00S7PajLYrK2iOitTdmprJ0iAQv+4qvNY3j6s4hL
Y9P0XFnbErG4wsiMHrX1yFQnvMXN6pIwx+He764dRqWR/pMtM6yzJvUBiZ2u5H/HaqBYVJZIOn5L
OTQdMOIS27JtoHFuYYNZ0KRkfxcvZfzw8J2ULfUe3pI3MgIN2r/zgTiUX4orc1pMz4JN57qEi1sM
3j5NuVjUje4wjedbdi5KtA+L6LhWajFcKk6XOPgKJqWL20Il8iM4n8ARx4+grnaY5c9JWympjfgF
dk/rJE/pDslT4YDvrh8oYtEJm2xu3H6OCRImWc4x2vwIg+JViUVBRs8cnDkBe56+g//iU48UmHE2
MDcc5o5yRP4ezArvOlYXauOw9n8+b1Ucv53ThJUIZgva//Xl8tfswqi6j1+ZOTeujhGVN5HiII7E
sjsqHroh2P4wwmMdxarYXFCk2FLNSWS0SLzUJw3hmY/xXfl5oPntc6oJ/XmfYfMw9EwmO+MPlKP4
nUl0PjSFCateuIe32VTbazrCQC+4NQt+lMp9YLIoCSgb/7BuQWN+kGJII6NGZyoUT7jM1jPPRb3o
qMyonyOkzzBIqk8P9ALh4+CVnhsEHpKPpcwIF4dSPCfw5FERshy8MMpb8nEiYhoCMTDb5oFM/+i5
hoCAfGWE7MYdaRA/pGd7zrrasMl0t6OILbHBiewxhFA/MC77S9v+7v/RRzZ7mRB6g9G5cdaJb7N/
JIBt869ixkf8loXlfLxzYfMPqlsTfmc0ITRpscpBzqMXZOk7aufCofW6ScH+SHzWrZVG9ODxuH35
Gr/giFTxEhjoaBQD8bIj0shUw2CWYolZ4woP3TZJ4c9xosVKGMlRJYbLGLhlKWHQYv04QV4QUYnk
RNZ7IF8eZtN9GDcAYoZIBWiZZYDxpYf+n9zgIQq1ulju5Ho6FU1P6tfQUDhF17IbKwf7k4jMSX92
eeITimvKW6hhq6pQLQtPK0+N/70NN2s/7ttXPrrh8q3JH7HqbdZiYjJZ0QyJSoI5laKjOVaAmOnD
BYeblPzzvyLrZKEisEbzvH0h2Xx/csNaB+kn58KxrR+VPurjGnm4znWIbn/yZMZXVpF6eqcNkY7E
SF+0G93vUJfQkKh3idvoAjCXOAz51CqyX41nPMYWDL7/nLq9Up/XF5kIosfM8r6S4QIonFcKjTaq
gmPlxC6MX+8M45ilx1JqnUV6/R2FdoKAMgx54zmQWCy+1JMqwrDIhK20LkvyNBv08izWpgoMghrX
K3kO0yXMDiOP33npXg2xcIBX05r+Ay35xFSsIomVgbkvzCLnAwo5UXpL1C6L3+Tj7/r8mxXvQSkt
WJshpYSwDL1iw+w/dLHakMNIOMmtbydVmBpzscS2lE36QYkSfKY/HJ9cTfgexCseWP0i94mFBxLl
uOb+N4JbrKdIpe4ZyHASPyVjt1eE/AG2Getam7O7Rm4wWuaA4AGTtoCMRUTW4HZ8emtebUJpjhkg
WZ1RajFlNnWtt6gtz3J4tWnUJPdf4KyD9KKf5St93MOOa3keETOjYn9+CPGiuWf4vWkgiDI/yOBj
oFpESVnzcO50Ax3MPzORdEMweRqWIPucf6qXn0WbjI190N2iHO3Tx64T4Mle4I5NNSdh4shaiP2W
gDuMQQK3cDpGK2ixrtghMrnkaRO/ImE9Rnm0yMsKDvS4ZisbQAJGR4zcgf3AKzcIRjx9hWQCTucv
JhoJiUL9d/NTSwgBKGPVO2XUmZvSogMFqI5fseZKtt/0+kh/Fy7V3aYTUqpWqkJ9uzbvTxUMgRIA
g7ThlrGwNJdmI+R6sdK8+bLasQ3oL7mt3+4jAGAHrYCfh8QRJVnPAKw2uuP1qIwmN/gk7L1Hmj8E
ZPPsuaGZSBlUqkAMpqKoISPTPlHU+rIi19HfZs2AVBhh2olFj2xiSe8gx9qR9rx2y7SKHb4uV7Xn
UnWuQORQ43PGdBVcpwHbd/CuwnmH34eYf7Btqgal3jS5y00qdNREjQpW4UDGHCKCRdi/yOgnDphp
ksqf1dQnkGirnJ74Tq+s0xLWbposgbdS8VgOAkZ4JWLtG9eCfmC2a7NZKNq6+RDbTfxfCnpoY/CK
DYkzv9xfYAEsIrsm27kF2qJtOV9PxNnn2cNsEDoiCQqpJzP0i3A1XX2lFVG3MfVpROwH1F5HjTkb
4MKUzHrnI2aBVMADE6pbC6mFvE6ZGeNimqexwUoEq4H54/h1Oq/+z1QYRz+uOlPhxgpuOZz/bxgS
nK7hVZvRElY0HJCp/g3F3qH4wB3q8auvec/EhRjCwLDUuy8BJerkPhG7aOJFXQjYp8SrZMcMbykB
Pu4Nt6oB+i9CF40VJrSS0cBqSfHAsYy6rXCEU0LOC/P8FYYuru90LJRVgqmuwBAqXs/eTWqomWUv
89tP2Nz/4y+19AhDtsRcKHAtXmksoPAAXq5Y7YSZLRoJnuGA5MzCetJoXAZj4JevZ77aGf5AT/GF
KdpzW2KAflliAZqOIFK0g7ggQHCjlkedPo/jbkCUzYNFpiffyvujSzdefsZvKoGz9mEo3OefBSza
vXAH+b8boAYpE0E3PU8606atBY5DnqAvGdrSW1WyFN2ftPlnHiAUT71x0Gvr9ESznLy14axamugm
HLFGZ6wJ3cy2VAZmdhmfQ9a1zlLPez4lFj1w1rJ4cGkSY5kCpzCDLV07O/aB/qXfFT2PyX8qr/cQ
dFi9/mMH+XUo/NO/QYlpO+joeF3bVLlcIGIeYW+QVoex8ia/lk+Ac9GNxAR1ZCkY62Nu+ExGBm3i
DwlYGfzS08Bm/BAtJNoXKGyQxXMaE+ncJhvZGWNSt3254NelNxVuVnKTc9GEBLNRECAAQ/Apb7I8
0/9L+1ug1iZ9+P9SEmIoBko0PpA7GYns+sPtBnXWdh1Og/d8IwRIO/B7PaFoDLIEKLoZgqtyDMf5
fIVmu5s8B3AB9ddr7xc4beB3xJNa4ldHd3C50l+cXnVvoQv9S7knrXRUciWoSZLiJTZyYf+h3JWL
Yt8prAjWUOJuDUNefmbrPfFKokK4JA+pzeNZBp8BaKXV5O8JQfdjrbec5Om3r3i6RVDOqVlhsZXc
JCXnm8qgFscp1kn00DPTeSA6NSDriYniF0F4jRqtUZUI2nTdusKZNXkHB/rPx5hmIIUc4g11+VIU
+vlREbzJ8h1NO0o54Qv9YEX7K3lvv7Rhv0bGAQDV40PTlaQrIqGkZ/AlX1bbVYY9JRiXLzcdKF1n
zKSM786altJomu0lXT00sz53QnUm1Gxx7iS994OuPs+41a1LGKB0oZGcPwfhsam77JrHt0XiL0RA
y76B6jE18TG1K/eLLqvHkKEMINtfNu9XQpCtAOD6NUXgB6iG0W4JegajBoCoDxJxzn/oBU5Mk08x
uQkAddRh0qlm0PA5QTGKra1pPfNaH0uEVYWMflobEWjh5JrjrI8KWQL8d2j5I83R58Mod/r+M486
KfxWmjZSzbsfgnCsARz6cISpQ1smJQqpTsNKEuQEX/kpni/11RungnvZ7ApvVH9YKeucilmiahv4
yNRjohK/FvfoIUgyh/p0ydKXyy1fDlPgMwsidV/MygyC+cbuzpuqludVMjwNJyF1zWE7molhSRTZ
HqX/0X0kSZWHn/fevcrbjAwmeY2aGZpfH8bbtJpIMIgFnrB1ecuhZwixsUokxGZE6x5hsM747UhT
bhF5e4ebrB9b6pBZOj3eLez1bSDU27n0i/cgM73eGKA7hEnFsMPQtdT5N3rd4DGA8Ej0LJ8rDCOx
RLGjDzJblWVDT8RkvK7Z6L/blDzUdQhNhwbjDqvfjzLb0UsJeWV0nPc1zjST3rLmEqECQRu2rPhX
adkXd80UoF+TY6rTu1QYXGcd0dM1ZM8FQSUYY3bUwQgljvVQW7Fkh5u+EF4dB98SEJVcqQ/DWAol
HSaji8o8snMR6OfURNB9nVG/r0X5lnG/AcK7UImQi7whAX9hJVP+/+XcRCtPZbFpVr0G3WM7tx9r
PFOFLamw11NIjTPZIzie059uhNgHvv1xwW+EvTug6QOlPlT1HrDPKqN9io9w9giTNGWxtPpE2K0c
wKYOplTFdn+U2A/mhNB4v25hl9Dpfn4VkdJpsuS0yD0QyDIQyieegNsP+8IEYHK6XYu0uoAI2Dej
C2BjyTG72LNDoA+nn/bBf5BKlQHs2rLru48Xpz0CvuYxAhE2F3isMtmr6FfQoEMJotZp8cyp/w3p
RbUQ3OTKKHR4rwhdQP17MyRqfnpIyE9q+AYRbg2diafA8Sc+gmm2YHnAFXKOHjt+vUIUZrnYXQvQ
XqVpiI+2iati4FM4NVdTbV3dnD+LeL48n5PXAY87VsFIIIHkQ9ecoeJEmw1RwHY1cPRnyj2YulBm
HZLPrOHFO3DUBjrTTFGP768cTNGLljzHiNWkF9ZJ296nGjMGlFVLPb0O/7rnRKQNn+/CQvuDbvH7
vW2llT9Hx2iA3TjsRlCJDaUu0QTixhGGq4fFEC8U91L22iCEj2XRDZHr47SBFfdzC7dWycr5Ro9C
qRBF3liLe6o0yfPd6UFDBijBOuUh4LHiwHqwas+BfeB1O0yHpGDSoFrJvYXQOb+wbslG7loya7xJ
eYn7Wq28rUH2EBzgIR6CCTGLrDMjbJKe7zJIq8UiAZX31TVAmZjttGG6zB10ViVvXkizJOfr9fap
3577sMbgbYIOfiUGcR1XBbpIzltP8e8ms/u5qzBzwcaKgqBBznZo7E4os5NS+DIMRyzRLaeit8Bi
t7CEqw3obgt8h4Z+0XvVMQhvgXhE6w+byDbJTiOMbENyHe+Mow53zE0y9zEwNVAy1biI6SddkhzP
iFh9XSoG4MXNb/n5/2HD2i29ziHRB8EILpjm/FDAnp/5UlldJRVo5VbTNfGlBQuXe+RKrNrlK31k
AZXMkeV8wRBQ0GeqHz84QaSoPklNONxA+cYMwG7ZnAAM/2eTxgh/rnQnq2MUoWpke1GTglhfxLkz
Er6gigZcPW36EN3ffbDknQNsccAS5JlZWR+fj5qaR5hEhOYHQtTjhMVgw7RyNwcpVonFVJ5PkdH7
mTd3sGHwDcaqRfDx+RBLOO8/T6HLIObYXzajRvooIiWUQof7UIuZjbTjG8lznOj5kZVTWNsX+ar6
reFk6flCDxTsfaabvIHguCPxd5Baya4DVQqEQScLt842IYlsmcXoPSTmBHPOoRw/WUQfbenn4UHF
gWJSTF3j+aVfatRgJkmGkfbAAhUEvXAown8G2o0fZVrgSckz5Gx1P6f6lNDhOQCkNJKuu1Z12AMm
ESqSQXDXJX33NC2YBQBKKPlGOrvWjK+FtlTOrgoeqBVGb/l5pV53v7vxsMBiHx9eUhwue3O3BCF7
xmIBFzJzb9MXdXkZVoh+iWkYsmp7veIQrQd2RPojcEkHTOrojLnyQx6KMgAs8veER/yDRsvT0atK
J5o8M0800qY9QTzkRVNOykxBTHzavcEqEWf++kKJinx8JFEhtUnIuniskBBZ1xRIBERcoiQWb6Q2
zmbhrYN8tDbWU1LI1uVAjBRzcgB9WCiY6lYfj5BVCQNXRfbZ9OJ9CJx72bb2xySZegCQ2Q6JE0lu
S55AlIHgkYPmTsactiwtiB53t1TSHpVNnFP8SyuB+aTGydk5GcVm/fdaO0gEORC4tzeZSj3ist1k
bsThfILt/bYM5ZqCTXgwtGsr2lNNTu9vqybUJGzwSix7UO6WXGgYX3Rm8F+Pdr4p+ka1schx2qX/
2jBeDEKwo6PJXPNu6gidH9+7Sgi0jq3jWNVCaAJX+EkWpMp0v+gtQOKiZ6B6+8o2CRmyLVAaFGoZ
if3NvxHJqYArIc9ZeRJfIB86pQxbt0rNIHdNDUyf49u4oTogjuUTSr/sfi0BqQOyRk6vLO0buu+B
uwVIEAFu1edb1aSU6qxawJS4YFJhfKsEIfvrcCYcOCYAFU5BYXyorCo2UTqlvfW9pLr8hx+54/5Z
RJ//+nOJ8FZTgvnxm1vw/EuA7mEJ2VIxFtLISdP1m+O2i8JpB8V7EAApjGQpLBBSvJk3yFrc2LqP
LC1w7BheDmxT0ViKejFx+M4BYPZz9U63MwaTP1J+E7GirC5nzPowUoTeZP7Dev79e7pJQY/lz92G
hJF07JwEKkxoK9URsFuthiT5B90UVG4Vnn1qPcmOJSFF4Y6Zys6RCzx4/4X62Hk8xf9E/Bpm4gPO
Im6ZxfL1TBzINp4t+ZD2ZO6dN/cCXwJLCbBskP+oiqT9TC3H1jNwDn5nrMD9IXgBcNNim/Rids0t
rRJ44HpdRjELX3AU0vW4v86EmJMqsbR3O/7aKOS/IsFnUUNTuFQ1amgN5eY3R/tjk+Q8FJrb1BPJ
iL8rk5Vw8vFhkMX4+PiNr9frE1HA79fEoD69Cf1XvpZW3IKuXecl9HfnPhXyj6S/ODzDA8u18ynq
JDtTipmwJ6yRdgAUIupGwLSz1TPQphz/thjg8bASKJmZE7sBKMTsqM69WVuHqsohGpm4lHOmA9zN
teEz0LaBTJERVhp9icYO/xoyEylHgymFxsmpn5yPIIpqxkZZuj7SD8pe9VzI9A9SWwpqSOJeS4bW
2rayacfVqFbiCZUKqHCoEX8lx3hoPcrwqyO3d3KNzXyxjeUm/GVgVANdnoKOV32CZURUZcfYkTrW
+t97tPGpuIpFlZ03B7d3yJOoXUsHLzPP8p91L5L+2wz9dwsG+M34aQjsEUHce60DaF9yl8G7aP5c
P6PpUjTuJHeX8E8yobnYHWJM1WQ4od0swO3i0Cl1gVvZtgBCp7WDf9KNZn8OKGkVrjs+7uaSPgb2
tjjV4baR/X+1jJS2xcFPfYqs4Z/16xHga2yp18jBukgWh/zo26CVYFbwa/9zlTUg2TarDcxTfjJx
frQ9E2EKvxwlqZ7QiKfNnX2v8IM+hm0uCn4ZmKbW0AjER/XlG61sWwB2snNdg80iuwlYYBESD/Ld
WJphYA0sH2bBzh7TQ/pFavvJC/A/+f9ZSsQS9AMIlGehhhpBNAAsLa8loLWKSpOm9h2Gn2SwRV2g
KSpuCFGZZLPEmfe6Z+IAUcGTNGDmMhHryjVSqcqm8Vf4FyMlrukJE7dx/wtux0iZck02qSnmdq71
NqddqxjA9416v5KDlYjiIbzXwewB3sg+gVmfaUZQjoS0Dke41SWDGhO0fDr/A1tmRXjrotWnHdSc
BXS6VjH/LFbnR49RFc/zTsHdlVf5F0v+QTDNfIqTVldh9Dk+Kw/lmCx2qaTxRB0GCvGsHIi1UIOj
Ph3BoihDAzV+Ec2Ef3Im31S62S/UIQtAkI8hoCjF8cMNY6yLsFgO0/QFoNkvYXfGIivJ1sioMg1t
lLWNNUpwJGzaNuUUoMqcbA0MAT4lZQGo1zXJcLOzjCyG9zGyPBoLzotGORgSjwcnXQvWmkUB1twY
vj84O+UfqbzeCc3NYIjN4MlkTOyEuIBk2GQg8v1Zs2Izn2OXEOwOYtdzMxpj+/PSUokbilykV2Im
ih/GYULKQHol2shbIUlqoI3pQ+KjC2nia2/UOrJGdawc87Mp3gynOsQfiW7pX9QvrroJx8Ya7Gq8
EK3o3rrhwNjzJDNkspHVTSWPauqex2IbtNAkTcm2g8aoPsWJwtA6EO83PJ52uzyhIdiaUC9ay87V
YKW3wKhR6mweR6rbHrPZk6U8wDBKQq6o+tSz3RfXw3wF7rJYKNk2b7GkeRK8+WjXteNbnHd4bSGP
F1jiqQJcg+VYO7gm5GCBO5VdCeSDlPAoFOi0a4xfVcyKNbhCmNISwBIi1B3WfgZ8i3rGuqUoWX1R
xlzTCNaC2H2EuQraD46c/+Efl1OTpED62YWLDwZzenkE+vSYAEFSl2RC6UuecRwCUCRsId2GJeiY
OwecpOhabmCgWBmLYRe3NdYJacmfA6WuOxF7U1TUHSStc8zYPsC9XohxNmtSmN8LFvSP9Aw23eoC
jjHM82ff2N0Y1AWfiRG+FrlMq5uDsb+pfBvUgigJvU8RuLVL9WLEo7JbJwUnW+lxkU1mEwMq+/ux
Qgc5QWnbY3Ivte0QJINpx0YrdC3AwQ/1YOYXzKCVb8XF5pUlIU4b1GMDD4b4XYmtgJW7tlkoHd51
5ZWykkGvHszRCzOlGWPW3D6QBhlQopzgxW7KHKh4E5r2jL/qn+M4upOQMifuRIvdDjILjM8yqqP3
qRahfVNP66iP6VzdPqK1i2RgXZxBTo4njq2eqWUQEFlMe2icVXvG5DY+hw38ehomJhZVSiwiFv14
wciGcUZZIFv5q0QiOldfiv1VN1g/QXSruYg/dFLL3kmrn6/iBY07LKRZB3f2E+JZoxX7QUjWCufe
hiXlnUW0rT3salHHpfdl2RrGlN2cQDnTV3e+RZwbAgYUb2GRfH02T0pV9lrdCwTBUH3uG2AAKd8r
HkqDb/tylY22aoPdUe83SCjuWkI3bLJTjoMICEMSrsYrAOpEQNWBg+3201D1p6hON54l1e6rjA0H
qwJvsHkRl753v54ydys2Zqjc+7SSYAJJExZzYKRWhBv3dO7JV1bQRY2qOzh8DzxUuVixPQBvciqv
Cv9mhzuf2JCzfbxNrPStWm4GjPzKz7jYgfXuO94Os6usbvdM7uLAFdsAwClysPnOjhwA8kWZUIxp
TVSn2a5IG2F5dofUcJOUgMA8I/yYHuCOj7vjBw0KNPXzmza9iaT0mrE+JiTsfiLjNsnTPnPwKFDN
VBHAPVbFwTgt5UZ1uH+Cgy6mRrBnBwzlYk6AQyaDS4Xy649gEKkKvYV/tpguT3UDOX+a1lCUH6XO
Eh/A6M71jlC76JuotHj0GEwFmpoceZsa/l0ISMHtoh0Vz1sKjZmPjeJ80uX8tRx5GSkVDlcmG7Dp
J0SO1CT7GycqspxP4+/4Q1Zp6ivWAtATST/sIOU31PAvWjXEkK8xvuJNONiboqsOhN9yBkSX+QwO
achDbxDtpi2RPbVSK+F6BwD+AXpciC8jJNSen1wtzCMpHEx46sqRkmCSn16KBXRV6bdwaqP8V57C
efwqZ981VrRE0zRXK6P+IZQeim9oxSVWhyT2pjmKCv5Yp0sMWGxaLd0H/YoPvlx494GWNa6nAqa0
u9jIk0kyKNkmspC6uSb+/Jpe5Fmczete8X+1rg02yUB28hIZER8Iv+b1TKFAkWmwvn1al+BnDtPh
nTU+jTLGu55M4IG1HUpX5PzjRr5/iBE6tTCi5DR0dGnkWsFzfvOuH3sikxq9wpFnp/XRIo6ZSCCe
O+1OzRI2vNBFjtBO0wNZe4XZMtItpZq6Z4dLnqwkMlLA3cZVdStncl0LQbrPGb06/nw+/6AKxk7h
BMBfrhdJEiJ3D5Rp2iMRgkLzp6PlmE4X0TKX23fpNi7whBsSVZ3h9rk6h2Vvanp8dHUYyTdbqiuj
64/Oc+6f56kfCWZAs9KEIbzlbIUTFdAPn+5JA4Ebntkt+TZHsGGP66PUa4TolQ+Hrj7u01Xx1FOl
1ehV6VLL478El9gfefzwbVYkt58c88nhfqpWktlvlUQ5WQoGNQwc7QjdVxwd21/vAC6rQ2/RMoCc
r7Ng0b34uaI/jt4VawWjzNJmLQI1gVkDF/iSvGt8vjl+zm4OidB6+IfLkDu6liBM/c0UKT7/S07w
DKhj2mGrlbFlEfYC+ZDSoykDEKM8KzMHd6Dyr+36G5psEwdfrAMYD0yuc56dSZozuUJPp/EPpoh7
5qfWTSK+R6KRPQNUkVtsOfls+Jv6aN/I1rownAeUAqBiOfEwlM5qLuOl4DBM1wxvHJnJV/UcRCMk
AwH3iIKQqhQHr3ZSDO/65FD2hJ8D4pKCwcg6L5MxwvRfbGSreMkciHrkCrE6Bt7P06BWqXGlj+Bt
B96/qBaYYxye93OfuGDfd6GpVwdf1rcXOV2EoYdvQ7O5pW3z6POiKan4yB2EXKXC6BbBs6icbbpB
Nqr82lRxkY+V2gshzr81QofwF6h1YBbOpWKbsZVrgVuJ6OTqLgg+YmxWaJcYr4bVNAqX/c+4lRGV
zRIjTGhH6kKcasfi6NFsiudNqGb5Ot+PYChRPueu0qpouRvI/2wDFKqL5alxT9d2iIzDtdbD8X3t
Je7as/bNCFYiWMV0FGAStt+UzI+t5F7Y2qnc/LaKiF0/CzMO+KVcsXek68EeHpd6cTCvqGLOxBoI
Gg2kjJGzVBqVBapc3o6+0BQmuttYdTFL8sJgrRUPSLd/6MFpP2LhW516a+PzFlshm1f9fBAdXdcT
2VYNusanJUXogqOHayCp36z6o8Uod8TdI5P3dVy5z4nDkdi3AIY9oGM0BDwJauLqj7crM+l1VV2F
vUMtktzcx8ds0pyS11U6rgW/ZEOSMbu5jUb4jXG6IdJKf98OqfRWQ6GrnmZ5j0MlZ9CvINVVTjCB
KWS2u8W6joQs3pMDflaFX3Osp9cpBc4seu62OOw5w4CJwKmtAvhL/Y02skgN+i/Nps75AsLPItx8
8zBAg7hJRGv6Ymcp1b3hHWDZwna5ruv/I9yc8fCww6M0kILgN0TQ8Jfh6kiDb+EkodtxtvFn3dAg
BjzF8c3Z3MrbWF7NmDBYh4rvmabf+yE0YuwJj/T6e1VUuYy4GkmPWklsdZyXl3OYF4pengdNq1du
9Kx4ZZdumCLC1h9sjqoMqUdfbSSq+8LISAU7B2VL1pdVyiWsPqahcldg3pADhb7r0y0ZTJrq6RZR
ZMyNYx2Ru4Kt8E6vr8gsVMH3o/ucn7l4FPsVQeiM7AipkNgNPAckmieXoYSkQEd84/eogkjwYH7B
cA2tCyNejXAXp+uGQxX9HqkfCu18gF5CJYETd9aHpLk7GLc0igo3rvR2vN0oxrVuK2/tOGI6R1Mu
AsIFbfD3soy1v8jSlrC9ubWwzXcLVhwHag73DiOr9Nn4PShiZHOjGAkSwP/FomyL0TXOnEgw190H
SCmS3JxTrKrsN13fHVwPmI+X6q6ggweggI1Ylqkj/UPhV8Kuf++hqOEBjNz8LKbfc2tkDH02xVUa
L5MVs+3rR1gRqJDG+ajPNcYYilxOwzw1xyH+7s3d24fV8MTnH/x5RbuV0KvJfcFuKCFu0jQkQAMG
ru5qLnA0nJrYQT9QNO+VTr555Wvs3XrZICWeFgETyo6oVPSZws10w9OC/zrzHoYdI2NSV2t2inLa
jA7SzOK5kQqNpXgAj9tUTrwCk+mOLuzw6lClzN7yxsyFQdm2ww1q+a3NrAdh8EWcqXSOs8u6D+Ee
LF7erPI9FoXCH+I1vQ8Bn1uBxmGsMSSR1Nw0tcGv/ZE66prHYIdwxVM8Mhf4+ExAbjUsLRos7ocR
A9lBbfgHq8MRczYJ9MN82FWovKOLbhZV40dC6d6JTkw5J4NqKq/cS4vxKxs4Hzrob25t7mlBFmch
+47o086SaTwemxdoeIjuRsXNYoJJZsQC8knLbFHll274TMDJ5LKsaS/vpPVpmtxmwqnx49jq92cQ
HEM6p0mS288I1t1wQtaQfmLuktMI0vi75CUfhI6Y6s1cQ3Ny0EVABF5wKTGMEuhz3XX1LtUCs+PX
HucmXkqdzelmSsYoH10jp1zDsbfNMFy+uSaj7Yjt5YIfbyQEmcnUX72xyylLimIQX0eqac25tPri
ggmtjhHpXyUmlk4DbJf6yDcbsERLpH+PoIr5LvtzlPxb2Q/HuEQwGCfLxznR3GnwE8VTOs1YzdgQ
xh20/hgRiuoh3x3/OWtCk8pkSTl+fu9ud12WAn9cyZZt74FhipdEQqflNQHMUJ0JieiIk3yuOXLB
YzilGiyMMdv6nIAlBMWSa4+igJ5LZ8I7J3b4vyqCVJIRfXd7tpm3ho6uTvQMXzIbZwKaWYhcnLrH
GWJ65xSQrijPbjQJNsR8D1QhQruvRC7EIUYubAZS031r4zDJI9JbFC77x2D9jEsGTp7UPE0djy7w
5inS1dsXOhP9jdK8MKJNxYj4XQ55LuaxWnjdJEq6ym0BuL6O/US9hNVNee+fw7DQ6hBlhr8e6BSe
DDeQ4B+azPXk+7ogtMwgd1kLzL1iu7dpaJJLzY9ukqPGII8Bcj2SXt5xHS//wSotp/djsvk11ryW
lj8rRKpc4xmGzD1MlcJGqBNC/gII/TKmFrYItJit6Oc7OaaS9qtcxsjPFUxtTVaC8GE+nUARB7qw
0oNzGpTxkm3vjvzG8m6+DWXj76bcWa+9qatA6H7yqJoNgQ+8540FdahLLzGtvo+bZos5bQfRS+nL
Md9DbJNH8LJMS4HCks6AKHD2cadRKyr/DStXogxzCBlYGoWn9WZGzec6a6SUCc1bN7lVAvAULJbd
LhE7jn527w31Mc/mrDJGwuj9+kkBEIqdfPg3pO+VC4OAZ8nWPSNIUODVLP/j99XmIxPjOjjahHj3
cuGXNFS2gI/pLWMaVNG3lPoKhs8/YKFx9YiVxW4/HT0WJ3GbdBWalxZJgKXwFgwSpo/mHzl9ABkL
D1sJqEm/1HrpBAmNBC72dWxHVLCHt1G2k6j7HqqQbYYmjiJ+wHEwIUxq9yqpExNF+jrcK+zOyxyl
69FLlO/wx7YlwCqBTKXS/hUbbX+IErFC+vBNNmuY2WiU9xpXF2Myo+W/puzO77wW3/5HUPFbi6vz
CYjjlrLJTT22YUKjFZfpn7GsSir5vXPJCCpKxsuVsJbInjvlKBtRqdl3h6ajg8lTePRpsGIsEJeb
42bpPX9IKNAk9qa/YHJslqdWWFxIdKkaqUDKfvwIf8YD43sq+UC0P6T4dkdnK/BIbHXhrZ8SiTJw
SIfZswV/u/VhuA8xZBqWNqU2bzAGj/Bt9VFUB67xO3CD0uuDKFlmr/Af24IRdVoqrWf+fB/RRWo+
9lC48XeYnb3QCJdKIV7np0fi5gNASYbE40GNWEpi1cAge0M0srQUchIUnJBx6RPI/nkaJHLMLe83
4AU/GSQ+t2CX8Kw8m2fpIiB1kn6hyWgN+TO11GmZpJPRYhKtFVdeCQE/9KqW2AXiS9j/AVepmiSx
9RIqGpFQhZnOfwu2obIRHrbNxG18966qUyoCwFZnZXVwoLWSV1f9vSt31bLTFR2H4UvRj0iZHsX6
kL6VIlPSizLceA3HcFE4KRdX1ffuUGFhuZEGcwGJNmFuns8cHsIbh4Ywz8OOYjvh0/yBmSmZnyhB
P++VcFG+72m+8bJvaXsg0uijjyud7aoVb5Ku1G8BB/AlrQ+UXT2vFa8i012gNk38fvX0V6xB6HVT
fuFm/WVZGsEChmCl4KZU+34+mogTNPZ0nGBIeArtWfhxwM6s/Yzg2X2/Zvr7nF959+wSzRskItzm
W4UiHmQfT1HmTnX67mlPGe59bh/hRjTcoTkueACigKJJyB5Ge8Gv8wTGVtQz7HSCnLn7oLIM3eOn
PZwjUC4qrDZpUk1+UdXYIH0Y9c+hf6X0cfmx1VYnOISzQ1mFcXjZuL0X/wtj3uAvfC5D5HNHjZqy
5vy5G5AQswz2CYSDPgDaU8OQFqh4piPs4gifc+pK2lRgxgDKLftCYo5ufvC1wqUr7Xt7Glv4xL4X
u59SiAgJllhX/6Un3wayGgySSpss38z8bSj/6mke6gHj5IAy1eeSX4FQt2IJsD0jjIDCNfOb3R2U
AtTvrGpTywpCtgS0CfVhYz090Ygc9fYd2hRMHXFmd2KUmH2xyX4ejO6AkJZ401ypMnl0MMWZuNsQ
Igg9lgR7PZgNrFGC3CIvj/9+Gapwb2jPSbliDT+OjQ8l5bjHRIe/e2A8OhEQsprWSRIRaUQfavEd
G6PqCv6T35IoyIR4yMMrigIg1Bu5HRXfkGAIzqt0J8AE0ZvLtodzEhvi/wS1ZkCGbnG3KAYcPEG3
3PFpUJWsULDMOi8TeIAssUSJ1taAiaTZx38o1bBscpW70qQKkW8cDQHdVBtEmHnwgNgO2Yuh/xMX
cDFp8oJIYHxdQMWrzgoWbYtmkgFCK338aO8IEgqxqB6KY4BIaX6jeJzhdvePfHLVNlwYiBdsUqZq
MZdkDRAMyqoxOUwHkM7UvD6XFdvhuW08Bmd8fasz0HLdAw2McU1snKLPjN97FO/EfvYHYvRNTq1C
s83V9dLd7ZD7HkbpwwcMVjYMNDzku8uDPTfXNynYTqwGfb8FFv8WRgU0REMuSuAWpvfkRJ7EpTn2
u6tv+vTjFbBej2ncmV8nLrxjy0M6F10JQhj77BunlTQq8f6VxD4Vzl50OmwH/UyM7b56vYkiiveE
jL9WbEL3BkFtl+Yv4qcMZp6ZAA+AFBsgNthN0cHhsZLYtGGe3jtjky+qdiYPItbNi1X2rfEnOwve
KsGu5D0R2+tI02DeH2AbQm20PJ56duO2eJKOEDputM9MSdP0pQ2JNMNJvOup885UJayX1TPi3o+6
hWVdmFhPy7OAo6nDLHrYZqJvj1s4sSDLaOEN44ykWcuq0E0zy1yHlhZKpfZ7C8CQh5wlH65PHAya
Qp0IQJrrQCJXz2d+ua4PHjscwxwXolbyIAsQ/Ir+K28qIm6i5bh3/NeUFej2N8tusrN94eAtqoTc
mP3UcOxda/Roczv6FAfUlboxXklLrLvKSwueIfpS2EzXXEfpTrju7/xr5pMfhfdCNBUXWBRgyVER
/x436hJrhJWQrtTdWAiAcLnhIjrO/wtKJGEJSDz896K0Ha/4uqB77Z6KoIe7BV2QEPVWjHDVzINn
VycLZy9RH1jClOqxesU//4C8MXpN142xcjlOb9Ssilc4Ww6NvXM0ITOPJYW2JFN7+nUaLKIfgkXy
TSOfjuIUUyI0jsfr38o/05Iyy1t6OJAgnmpIfwJtO/1uF8XQ71qHWxiTlkHE9KOf15yhXfmnKYpG
FL9/K6VA2UoOqKJ7Jxc2T3CFDzLp1+GQwQlOFJU6PQJInDdb5+9vJ8Pi/+FsTMwnWa6rFBafuGvp
Bca1bhRCvTfsB1aDZoqF5s8adweJPWFIF7MmXjeQ+OU6JQY7GH5L2tBXTnQRNcAoGq4nDZSeQ2MO
i3xUSIDVItW2shlDmC4H8q98dkDl5YPtwzMnRxkdEakUe25uSSxeY2uVqjwcLBOYhw9LsdBt4Bwx
W24Wcb9c8TMpCvKKxWjMhqHv2oFEulXN1zJNoOmVOE14VtStQYhwUpRVpHpVnIsQilVQ4jkRoIag
aFHig7QbAiP40+qa4pBP5c59TnhrXt0KJhHxoWSqULqhx/SHvb1Jj9XJD3GZyRMPtAtrQNIRffLn
LENPj5IbbxQRCXL6inTHA7Zis0NWBpFQimOX7UFKhPF/CTLi3ZLe65jS+cCNweqsPjEL8WF3H+Fa
UD/UOW6qn9Z65T3ZYUEvZO684y+Y4NvQIHafp15VTs2nYxtgN5tRHToaSLqY11GiajUzsutq+cmC
zBN3WKtXWj+Pof80MWjOhhd5tQIKF5jVf3eeYyg4yZLTN6Wmr9FcWVRninGNI0EJFAVZtHco6B0I
WAP9BxrguaHIy4XZm6KBW5ctMChi0bmQANnahGZKOaTnjy0KY/6V6HNcs0zlwIlRn1QTrleCCUXM
LjIp4v9Jtb6af79LuNaok+YFKQZGG3HthXQTkUbt6eTWIjTfyqZnqaq3yEdwydg+MK2JGAm1tivo
XBfb0iT/AZoqr+nHqDN8VjTf/HbFI2loLos75ytRhn3wpEvY2nOUOAksNTRdXNzt++K2SxfjYnXn
HIIh7gSuWQRXACTbeWcpQO3u302XALRL3gFMSXXLMP7xkP4lxBdlK31vrW37bMHjDXU4uIWHF62i
aTVIsMFSBX73ydZfjvtI4VrNbmh42ZDAxlqRmLeyFzA9xLTWw8eyLLfd06OBZrZ/nVRycB1anStS
URAHCd9Uu8PfNa9mmQkOtpcDM/ul/sTeC2QSt7pP2+0IUlNrXavm9jVT1F6j+ZBNnvtBaWSW63QY
ISAvL8OrQWxSjtbFlCw8jSS9gGdz+nbsVaYj3J8R3YP8B0NFtMgZLl7x98NZ/t+r63EHBA2H/rdS
WIwzsbSTd0RLRlFGooVTfo8ePpl9WJpV+yEBXiRj3xBmMzkA2zaKCh2FBW+EwnDGuhK6I+AydokH
mJOEzKQzFqQH39VsN0rXhAeAAUqSRm3tQVdnqF0NJra9ruPJezj21DCcf8RGoqI602dIss2Pv33O
URmMIVj2vDUra3Tmy7wcFXELeTzKxBcNUp8TO0hCQaJolAJnzVzTpjI5TQ6Q1VSiV4rqIjQg+Xab
cmrdftnOM3zBNnxhgPhSnXwUOBdfDEJ6sEpO2vQwBxnJaMTKu5/Qyf819+9pHOwkf3fvrFgGnERu
bs7i9fn5N65z8j1+pq7qYshorKd1p6U126pY+JGfmhwNK8H1c3IfWLfizxSOzB/jMnX5S1bHymJ6
8eKrJQRnatcUM9J/yV5LgieNnahdsrUVYBRVACSOn1wdx2pvuZNWrfnyTgTH2NX8h92tgW2wuzA1
9HCoXTTONvfjIDt+3zJXl/Y/K5kxKl/Ll0aktVSL3hIrWQRo3vqSk7g0W+T/D6TIJ/TcmxPOzzCN
co9T2mBCM+nLNV/fSN7IAy/RdunMoBCElFNec7wZAw0FJH1zW9H5zwaK6KOd/XJ8izqyKvzHTrEd
XuhEhBSqXiGZfNMdDIu1JUg86XdFTt5Epu8/W6xmI1i7kunllbBhZ59huzCEM4PjHEMkKU0vbSS6
BV4B2HVoZNSpvWFGuuTUPHSMhvBZOxW5Rd5nRoUwnenQJ4ePmRpIZOJCBP4rqAxi7wShDNumZgWu
UQeXZPrP4CDa4Ncq1tdFYcipzeyWArJEsbD/z6+smxh7KlLSiQXV3rJ4AlI/t+JR/IF9AsqENO2C
2F8IOCmxYjHQazikTW9cvPK/jgj9rdKLdtlYU01vl1AX85jlX9CccYkWj7++zxVzU9MN0EIZs6me
m9MBhVOKaUJ/FocK2XNB+pr6X+EAYZcJ3ffJRAi+krtdYLjzMrDaOrwx+hzOLtFMy3hX19hr/Q5C
l+LzMxD+bLnl+l9qlmPUlXqFGF+WVUTbLTgFK0KzzmneNbv9mjSMIalMhOzRBG133ZCdPiO7iFcm
+sbs3JVN0DQJ0cx4G5nn2z/r4ee5IliAGpMuNP/RUL82t/1JhgbvhCMGZvSHG59Vlxjyi/pdvTR5
M4eeQSAmQNNlJERhvrCc4s9WwJvLKfQNAbfYlaC/IJIZZrEQHRzW8MZdvM7jeRnwGyuPhYUoA8KW
fEr9nAhGu3SlmkzImJz9eofkt1grVeaTYErBvLN16jSVPA4N9CqyL6VW++KgyNgIUv7WyVZREsTR
Fggj8wZKPhyaNdjyXDX8/wJv77LljQX/9qX86gqIrmeY8QX325N0bJmbqEM2z1C7XRZkxw3EImmT
Fx7dS4FnzTTS5nZNOgbT2Ty2Z6Ih4V7IZvDJ5+iWM7hsis6gHm+PI8c8mQFxaIYh5Z0XtQbh4c5U
wgS6+732wt+XKpw8VCt5wKOoRixbWjKK5ilt24nuVY034jMkkn6xUFFdTOfSQpqRqe5fyYuJJ1QP
sSbEDIBtqu61ZzE/yTNPtlQhur1wTZjRTYhvOgVWjWIwYZcFn9ca3z+DlEyjmNXgA9JE28+xI4H/
fb4HPVZ/l3D5g14ndDC0rFyKrimBK46Q3u1UKpYa4OQrv18q5UxQe3z278GkbV0evFdKiBYV64ix
Fh2ytmL+cIT4g2BYVaFwANMKhvKTsHQsaF9OuZimxzQ68YUEQYAEsvL3wV1sGzapwPSWV5tGOUs9
A8t0NGrIhVgXaw4hAGndgjDv69ZaPP57nS4/K1imAaNuobS904EhFIc0PTNEc4o7lJsxOqW2EIG/
biBQad6X4PJsqXx+PAd4oX0nZroJCtTrnQm+Mw2oOiX8J/KyQhjXfJEvv6wuRpwoV8NUQN19Rtw6
dfKrVmjW/kxonm4nG2vrxPxMgh2gRsy9b7znQmkVIcwp8go2cGZJLUx/YZyKRoXuxG98u1rHNgSc
7TZmqdF29UNWbZX+Z6opwXpyawGHzAsJGQbnudQR1/+lvggbJvfS3XMhI1KkLG7w5A+BqL3C/6Ve
r2XH1TlJOJ+/Vfl+zgpgD+9veCabmTDisAVmh7ysuSH3KVzaDfZJErm64Qs/TMiY9iePEom9NO5x
h80c/PpChfx4iewTrGSCYAQnV7ISnOX9KpjndSoy7YrXiA8N8mgPNR0tVCD0joLlmIj1sa082oNR
/5nuyjFBGyJA74z6jPb0WiwPcNzVmmKjMyrWfeqqv9oEpa/uDraaCIbypve2Lod09inwiVV6cGZj
+AOTmvnvPw1ybuLhKz6+cbBzHZ+mYmb2ESWBWXAWXOinGoOn5pisbx9K70+w4YwlVf6KHqWuookc
9doCtzi8zxwkzcGDshuktnbP5NYTSocsVMqLYMmCZCP8DVWq0zUQY7ViO80clR/9YkZE6jtL81Bm
SvgZVOc7ueeKSBpGF/zAYIvxhF4PfLNco4Pub+pU40P9jYvOWQQ/oZSFWR3D7jvN9JcNyQnrhojo
fUEGRiFra5kyonNfi9ryT60gzN3bDU5UEoJqXnqhRTBeYGb50qRMx0i+bvCboumlaF0IcOL4EwOX
eFh8IWRCK8dyaTeOuPX0+a5lkgGj2+f8sSk0XVilDIyVowUF5uU1lAg87nD+wlnLq5wT2qdYzVM2
glgqiO41QWmPM9/LjgECIe6nCfYj+SvRug81DwVG7mV74i9jhQbAPW4fyxVP12aQOy74Fid1VtR5
XaLP9iP/6y923LJ3DIgEUIHG4415SHoIIdnyAFcezYIyax1KBJwl35IhzapG+c5ATXxI3p6jal16
rEeNJYosuneCKXTFkYKoYk8nFn7F5xIToe9zbtPaJ3pkQiAJU7YpLZqF/AY6rM6b+IPFRDVziuVb
LPq3ipRVnuxofB8q5tGPnEbsuYRkyA++czfbWYNks6aYXBB3b/dfExIt0Q151sLAeKWEiwEJ0B5x
F3tTLxozWdnYHwhIeiYACmFxw9+RUu+FpJAO9gAY/dSl7R3Tp0+tyWCdY8+Ikn0mCVGXLiu8sPSC
FzYXquGq3FJXfO65CFdYQS3uld7ghlQovK6JoblKQFidodK3OUmMteP8PpWrSTPlPIRcm6jljOhX
oUfcsZesvxzlVkQLMHK9w3tmAaH7DW9gYwCr7VrFzn0UVdoHex5wdR3ryGs4CROKbUEL2ebyAFMQ
iHSF7kCOP477gDhXRo0OekyKMqGxvwy0QKZSBcnDrMMnBgmypwhUU62TUblEKO7fLyOcfCPycBBD
owEdWwKkSHlfHE521pbu+WxN/n7ie9R89eZ1C0PImsjHlxCA1N/GDjNnQN61Q3P0DjxcsVSFZxmD
gdSI4NXZBDZp+oC6Hb85wOGHPVnR9EyqrJTC5b6PdftRfZ51f+oaB0ZP8wU76lm10PKolPMmSGfT
MWbNCdkKnqQlNymbeFnWqQl8XY9mBro+3brt0jFVpvfoj5sf6ugP8gnZHRiW311PYG0KQ+fgNUlr
x/9uTcBHJtSe0n4hEVjIn6LUfPg55BaiB5r4gAYx0nWglLA6bZmXsz4YqjKHO4I+Ehcxv8cTS177
JtSXYfmy0YjXNTsffjRVbi8J6VaJddWhz4/nxMO8qnwApRJ+dm/q629qajqLyA8X8pkoMupMD7yi
wzXEpN8IN75JmG60WXxIn6HipLlb7VovFukhc34EJ2zJgZ+cpFV54Ot+0DOrPmx5SR4FbMZPr9Yb
vV7sTJorLiY+PvP6SOIWHEs+zkkXswHg8GQt7ZuzHoX6+5QV//G7KwdLj1obr/DPtkrOB4iBl1zu
R++2V8E8RfEbL9DnKy/cYNC2Pg4RzMl3SvIXZlK/G9S1JI5SefjChoWIf6dq7IaB9ZrMAnbABwAh
sHC0uGz0qf6c9YBwhsFHUJRUC9x8itdFK14JpNfv4iord7T4RvhO71gscTCqM2VLGZCiuI0uvdd9
DrVpGTFFKjla9zI2tUFJRPKjwPlfLKEl8dPquQkQIDk8219ZU+AiRIDD/sIvA73LcgoXzkCYc4x4
eiYaIB+7SWcq2IAN7vxdZUkHZ52n5DXeKSDdD08/EBl2++AVGEAttuQ78+6zSaVGZj8YaZf+L31o
O9uHOwTBI+ri/p/5h2Aih/jlZ/iy0o94byKtL4EIZ2QioKMzVYB6gyCCTadN32crBB3SFg3Z9Y7R
O1lEQPDaBBGRLmYqHo6SEnoeuAx8Qjd4gRrmkMDeGHciSV0fc/xuXkYiAUC4yLs8d7Wt3/zEw5IR
Y4R7UI48xCqm2Hy3TcI2+I050PsFuJd4yyqtk2CUKxy00Gw6HT443bM2Azmm/opE3oKBpYf79m9W
HnujdBVypiTdWN0QJ6LRGg/T24xUvcYNVp/5iD/Yr2WW38kpvLnVPX8AUHl3J4S8a4md9MFDyOvK
CJD5pSapf/EgzUGuzVrT6RX6erioEf4Ldh6mHfrS0TcXvrFU2RQEn6WIF9mr+dFrp/rmOWRXXwmz
j5EB+YeZjMF7dMBEnWjw5q9Ocfq8E3w+G+it9VtTHUgo7src3qbbwg6Crx3fMsojKBggymZktPS1
QvG4d17yOtKLoSo4BG4gWM90vp5hV8HqlypqsYw4BWSDy8Mbs2xzIkABRb/UGVg3jadl+nV0siFC
Uknz9eJ97Pn1tbtcjA9mo5W6TNT7y/4kq7ztkccWnEaVz/tUuv6jjf695XE7RxnQZkwvm7sOczII
E3DVt7qG5Ec7KBDgbrIOod55C/62W2O5VQG4KHbfbUIOT9faxEC5IhswFzz578zZVWk6Zb66sjXW
1oh8ce2eMYsA6LSO3snKYkjsDFAJdZvKqF9jIQz06oMkJeLmsuBWo5KGUccI/SG0m6KT0+9gE0dq
libCZ2DABG0Dv0dmRK8XuVygXrb4qDylZ/fBuyaFZZDkwmD+Gw11BR2eLH0EK4wPDkJaMEMQN3Yv
1PnYkgwzKdZ0vDJ5RfHRbQ8AibuA3CC0TYgRFDmGi1wzGoqo8OU1gf3va9/PXOuDPLHaU7E9UwZN
zG1m3frvXKG+8wdjOm3kFWxMyXwmaCsgWOSOUfMyJcaDKTbny/UF0uV1ciSLnfK+WP9sCbYhqjZw
ufbCtFAOaKFX/r58wGSHF8NIduypV1PXj3FwLLcFYSGz5IUKh85Qrzv9KyVvVl3lfENbZwLKSMVn
cb8n6VrADIT0i5/g4K5GEUTUX42geGsWvH1tKhtAXJkEq5ZKaxLTLZKYak83HeJ9FADZ6f67eM6v
JGAA9MPCYmtkgDcVAr9Z6/YiFqF+8AeWq6NHjWt9y97AxOvgXsDgZG5BmUkU5sPAC2uVCjx/+h1O
TGugeEwoR650HV/PYzTffY9TwlJerpb5RJWwhlViIAk4e+wlC04cpHOLRByo+0HWRgOp10udhp80
6wCDJnwLfwP8SEevlU9QwVzt3/CgFjeSqMMH+x1IUJf9aDDTFFOdN6QISfxewd+1ZjanpN/i+Npb
R8f4kAjyayF17L47nOEzToaUhfvOGgGGSH39JOQqp0oizkT89FAPpqVRL0XoXFgyOwjdYRkLE11U
JEY8dMcsL3dAKk/++iCFFbZk3NmYZ8Swhu2aaJcGSwLJdaWq+INtY3VY/6dighOlO0eXdIPLzVfO
HsGpoHTrHyi0rb2whKx5F0ZhlUxiuLGomznXNeb6witfPsG8p4owD5hP7/tiytsXGFpfMm133roE
+OL1qScC/unQwFRmxXXO990OBdHVJ5p33+688/5Q8BSm2+t7uebn4CBpc6P2Qb1UDrUNqMKtz8nk
MdqAU8ZsAeQSUogUZuQIl06y9dksfKWedMd8mnlPo6s483GWXllBMGMgZLKyJJ88pdUpTMklCQiH
puOVR7vOxGaoA3fCAkSCA56VQ/KAYvq4/aMCtnw86N7TYRtUL9Ca9xrsysWTEEhlqi1hQojzFluZ
A4xi71Gev/bYMdiZN+REPWh08UqbMZV49vWpbmCOPqz/VEQQcR0K2c2sD6f2F8xfXvpOmj1eod89
YeQlkpUP1YLGA90RHYg7I9+nnBefM5A635f1tZ4MvTfgJ1R6DLcVGborXvJYdUQbUx1tRbDCgZrs
wMs71Cz8+4DBxeQM53BMNLReNMj4P7vWj06787SZYoZPEfPO1biUDPjz24EaxNsEqyCkZyh6s9DM
nXXqyV6JH8Pyh9HKGRgH1Wx8C1lvuD+82dLfyMvmaFavo5NytLYFDYH5CILr6pIZzWq9U4iyrC6J
1rwj9QAwHEbmOXvrUHsqPcPZQioOjiCdiFeJzpPYvXEDWUsIDOrIYoE7uQ/p4avS7EdSzI+GAiu1
jfOcqfGwuvP2NKfY5jekFPr3ib4uxKvOhOknzkbN16gbfmI/1E9Y9CEQgBJkV4EibifDHGPZ75Iq
qbqHIT1+SJXx5W3044mBnf7mzxht10/r1rRE2avZcciUgiaUIflfMTmtIZj7Cz2vk/LgFdOXXDhS
PysIjoIZmGso0d5xNhBvp1KTLbFYq4q/J50oKgBxi4Tiv0p/zCGW4mQTbMDV2SZ8phYhCWXON2ra
8EUTfEarkKCIIb7kg8vFN4o380gZPg6cZ5MiYTBF5w0D62s/agUAuFEWD8dKnuftOUQmMCMy+BnK
qCGCOO8eE33m/Q74nhfECQ5R3+c+cIk8y6bo00v6AJ4c49yzDe4HsUHvVr7prmLLZ+8zWm7cAYNn
iY5y3IzIXoYf4TuCfIio5Rxl7ibUtPXA1Vfjr99EEUNYcJGg4/YcyeJFCpEPRMa8/edUEKykW0qm
lNau7yxJaCYdch7SecU4XbB5cktRgn93qXW1M8I5ZgBS//jdczQNClvsDQXYdHTNUymYp+zO7+cJ
qY8PsB1W+sdZsk6yGgVsxRVnXe23c0SnGFLolZTZh21o4EPIHnRTF9IiRx7qK9c+veOIcapOU1FH
EGK7sbfzbTXeRp5+HrY2uNUnlBYACFu7CX/3r9w4PN0dn99adIoMZDli0R13TDAtRUNAEhVR8l5N
5YBRPDnAzIu3bGro3n/5gIL5+4DgDhOvKrOFp4N4RDhjgLZ/YSax75s5FBD3NTOpQk20ub8fB/H3
uVOdHIw0i3QBRRwO9oPWreyeUAxt1JzCC+Wkuo+o4xBfOo3Ialt5mIaEyq49iV9uRlcJA7sG98Bd
2QcE8D3pbpgvaN9LusU7zB2UClABDyr1fDNBXL80dbC2xjxLERmClg3FoBNNw6lxkRkFlYXabgVt
SkBkTvyZ2g0nyfgZCQtFys2IAEWuUmkOFtbxHysbVMA9PVApPiYdi8qdALGSF1bHJxchl9ftu32e
aAl7VNfZ6d4GrV/FEs+dD6o6jWLkxYd/wJnL71Md/nEX3RqkLssctCV67T/k2X3p26ZfFJFYF4L4
TacMasqzJH6v+dhN/I0slBH77MeBlq3cn74jHsjcILV8lqp4lLcRhsZJ/WjpTPAjpWOVZAgyxMFS
rvPB7xJnrX1DTrtR7CYXlwecpuElvqIVOGVsLgVQlHqfnmP5Wwt9T2j8vX3g+vccOFTmwUgLWdrg
bwV7P2vb5L8dWnF5GUGil+HzrDj1WZIYHxtfdae8mWCfsAee1l4bnsTXEIP/5r/tzon0si+h3WCl
wtM31v9/VE+23gc55pB8WwJhdnqpUUkNdxs47empWhBacDVWGCYTJDXbgQFl5/TyLIUHWrYu/eL9
FiKs0s8YZU0pmGA3kcG49sstPxqOBGzBbWCSFZbpimwKZXSHq/A8TwPSdvB5fdRGgH6DAwnLTON3
IDwdWb3SMY0sEgfD/9T0TDIZkDQLKRnDlaoLuJxEIQBZ3V4Q0aGopKTOkuRuwIQCroO9YQ96L/M9
vor5s41uejILB/wvW/pPme2pnwglh37+O9L9TitgoTMa4OGh7+DiDJyJp2A23H1CxodLc2d+B2aK
IZQERM3vsWf99MYsB7uux61zrJXrvatGOgagU6uWnBAIuGNg86uhu55qS6MZLaojBygCt5Xik/sj
2ejKD4l+dDdyxWexgxozsYIfNATAfVtu4OrUemHEJKeqjpz8qBvl1dzvvOLB7UUEd6Q/NoxYDHMH
4JMztw21xBHz6rzyvT3uDtrHNqyaxmzEmvVhIKI5rsNTvBw1SVHT2Bz4Xtn4g9fZBsq9FussOPoL
EpQgYmOhL03CbBC7vNuXJ7SNgFQ8Iv+NElIimFr5ubwzSqiJ/VSH6bs2uZAJuCS6UxJVY8NEtzqg
WAQOExMRCj+4bbCksynLDX6D2cwaqXLk4AW/I3l14Bu/r4GScXQyhHWQgIFReok4LPFLcFKO8AEj
VecTOG8UgYLMGYrNkhGxncQWtTOd/k+Lz89NcpyQGuvetaHLTxFxu6oRy884VSzaVZnCn3tTQcsU
7AIkQkEsMQwCiRjdqQxSCyAtkdlUbBTwW9DV+lbbXzDbrgOYSWllVqSF9vabtAOQmu7ecSXBL2pf
hEz/kc2SG9z9s/n1AC9cRiXHjoQ48/6DLOy6N08Js8CONwbBfRd7tOdPO6wmc/yBVqKpisKRmUvf
oV/4YCi/3gqJUpyW1p5je/oaOJeQOx/KY+fNoSdqoZ2CbDnn52iZAhUKzbK93hmp1KsPAgLvfdb6
5qVlBP/o/3bYheIJy9aIs+GK0JQplEn1BU1ezPzmzDiKIDH8ofUFhCG4W7qiERXmI+qelVNl7mgR
b5XaStIPPhdOlyfElm0k3O2PIiNC7KBx32jdyUvSLEBb05FVOrOAOnR7/MZYHl1E75jWYGIL/QGI
TeyEB5XV/tys6+aLGIYGgkMSJ/VGazFMaHyVfwlBuupCzL/4NaM73tNc0nbYzLDyuJ2L8XtqZyX3
uXPYucfvWJVOEIKyUrI34UKUZSr6KZaH65vq6xet5gcZFU2jVDjx4+/0EhV/iM1/tvG900OYHk7J
vPP/4GuuGjD9pdifKnokA+0L6+8ta88mvusNgDzeo9/q7BomrneUS80YeuJUKMsLCR3krwUIcBbM
63hf2PwMkRhe4cXo2RuF7nQT9GD/QUfbiVJSJqg/41JT6atNCHdzoNWEkDMY66OH+GeAljpWVTxA
rPkvEDtWjWhGFPZ2SgNUlCmrDYN2iu9oL5NxynrRlpwUm0GYcWu2ardshGjXVdp8yG471dxkqMaP
gTOZpxo1bMtF6bCXrOxxK8qnt4GivJ4AVqzPQlDWqz4w6VlE1kbFGsyBOIaD1bkh+1LIZ2TKnECZ
jcPtLlXBJo6/drI+QyGCs3pdDlgkxI4VCunF8tKbdjHZ8cC1kgU8R8J61CMluvI7Ol2CEiZZwrGO
tm2VZVG4wvYA9MSe+z8otmJr5rKB5vMYYy8Z9TC7HhBpJvdaLisyGo0AJ/plREjbnlb9yRAcoJWp
7DlxULuhZ9ftAIDmZPPvvnSFOpBisRWaPI9B3SBaVY1N6yXgkGaP18PZGY+jL2k2xRVXRGumKO2J
pCYem/lgk3mnLa43ui/C6zL3hP6AxCP/LYP26qN7+1l/fV2QfuEn9ZBEbINv1e4KbnvExdNFwxcN
1w8kZE9IaHvipZ7aUpD8pd8OViRw6+WEAJLY2RKNeQ4RHawh0W2t4ldtVHZQ7FuYkdyWQ2Vp9Vyd
ffrlJjuXQ0WY1QhvpnMf49FjO+k+2/Z7F6V3om6hd++sIGmOCb6hEul3e7q1k7HZtJ0h2juuNHsj
Ve6bgKiQRyFg5HMJVXnXyB70Fsekz6LTAyJRvxBatBg/BWOHo2VbnFrZ+WHlCt2AchfnmQCub0fi
BYYBCJiztobfF9sepMQWLvXDGgFnmquWFBCMS1qkTJTqIuwtAArjCWpMor39XJ094NE1spQ5SaOV
D5pDRIlUgbS5FXA1BVdw5BUFds+3089oJRVuHANfpY2c1+36vRE0j5DoPVn9nzmd2gksEwDBFYNB
5N6lPoXVXCBhGBNAcT+r8qhIhu5u64dEsyP+Pk0ccZ292q2idBE4ttaPG51/xT+5SqXmB2wJobed
G9JWnlJp7FiJ293ODFiUWpk1EQIDkHjiXnDVq2l5RtBj4mZ/xHKbgNXPOYU+eRhpeZ4jp+Jogj41
y+bfIltpFcHK31X8ru/UJDRiPgLnIGYI8mlbfMMY73NXBtKTYW0YD9oYmeIMfxUMmHC17S971ooU
Ai1AJfhugOYa6V1wBFMR35aQsiu8OqDeeDKTKTnm11AbSdtrCXMhdQ0m7aviZvROuAqizabRgUY1
XCeqStCeXqv0lxfv1mv6Nl9C2/1t02GXA4V8qYOyECKPg7Jy2lmL/l6L9YZCiBQME84b+dtuDRnD
YwK/3BvzoMweW1ABkR0fU4ZgroR8Mej2ZZKXkKtki08dkvqmr7xxLNbOVFZrnM5ygj0eGcC2ImPH
1FWrpDRX28C69NHA7rhmirwUNsVWpp4+OgdIkJbYJd1LsWvaOEqYICunE8sLYUnrbTHYFJ3fOSHQ
N0OWOmD32SH/U4frmMGwSsyHNv4w2vzBAiG7hJjxFSAntd1Sl7JOXMIndlz5eeRm/C9LfugetTq6
BMLgmBPx8GOpjUwIRXP1u453dSbX1IXJyYGTRX8m3VDQpSV5nONPK4D4VA0UptAhgMX3UjD7TODq
3HWzU+wkK5QOofVmhGModIPlUwELYeiYUdtnXqHeK728hqFhTdI5/9Jm+EfmNTABLOvlx3xr67kr
BQwT3JOxLjYIfUZkyc6BCReDi+0GSF4fXRs0OCR7oR9HLjtKAZ2qpADNwLRvmNqSN/+ipx2NOkO2
K2896SmC6j6wXBnCNO2zCGIHWv6oms9+NYcRekBhUBimPB0JQl78CofAhauImYBHcXmNMpXD8N8B
6TnTq/GjCjiQ4EsCzG6nnMMuxJuLVdYNCbCgM1r+fvAuUqr8aCEZgU7JN0v3SYJ+nc+TK/1JoAcZ
uC74QtDStYrhh3FZMdc5GW62DoWdx9mTqmOEwcWe3uKKXvLMvVRzh5pHf8wokiSZJOAT4imQgex0
Ysjwx3IE9fLoMg35L9KD56KK6J3clMcAIYQmMGnpXASKFeGmuFtlDkliffFWH/j7edfl1Ymi0bPo
6hFqXhaugeXwAr3QRfDgivcrrHtpTsy8mcpolTUKiO3q9vlFy+2K26rt9Su27XLliYqp0lAvQxFu
+A4h7zW31u4YcPJccg5Iuyd5kSyGqsjEk86gWvpk5e4uWOCDy7OJtCCkhIA6c5Fun9/6ubeS4JSX
MuUsk4gpNHwFlA/RwbRzXgcugcQMGB7M7CdUQyGlhIdcva7dzPU9oJarffg2F3DwEvRqy5wfl7dT
OjWsP5qVh3SPGnbtqoAxb9DOBwkt20uBONHU79TaZzGviisLW0OUVE9k3cc3CYcXBCgiWjor0tCe
m/382wUcR4N+/F/e4PRQ2cmsVctQAefIdKkaLxxdVMEP817TBkTc5X2B3h7wPcVpYrQNgbfBh+Lq
ZF2CKO7GZ0d2iitRh3D7KhEtp3ht8K/Gj+Ch8gVekKZG47f8shXKZjRBSTT4TWI3ZwlxZ8+2VuBQ
NTAfHh5XMSBXgDi9RjUJGR+5FV4rYkzbsTusUZRB9pam1//WNyYKYZn+Xjv0ioAO3l/w10L6WBf9
L2HxGNARSe9kIjDj5f4OCtVv/Asp4sUtuNelQslYj5MxtthCTmKTsh9f71ShKgC4Y/xdNc/QGItY
rnJSyaE6p1V9vM2OogMBIMkNlxUFaSG5z9+FFw7bEGJvfEy59n8Zym58D1AvEFqNZLsKW+N9onBu
L/OJ46tjz3Yx/z4K7gpxg/nE+JyxlTy51r4xZZ0jROR6cCm9VJPpPX/8cYWAKDOHtMCFFqO96203
lHJ2fMqax6Wr+dscUVRF7ywmcSUMr+FD+BSwRdvmOn6HLHUklLWWQw3+cq8KZtEtsopLcIpLZxue
6Esu5n1ff4ZPG8QaEH6wbvmBTx9dMcSkwzTgtvLW1NSgcRNU9WoJqMGD3pdEZagzua3qznKxf611
g+V1hVTElifkEbKwNYwzC+oWY2QcGlddSzOszXpKVpP9M4lUrDH+lxDzYrbNFIThiGNf4HjpIYwN
iA0VXt7+xknE/19+SrX+QTyzNS8SU6iCZpDfv57kOfS8cma7LBjo5RKexn9npN1GtIHlgTwN6ft9
ZgupLEQpUpt9UmVHuaJZ6w1w3nEaeKEBJ1Q3ukpX+RY10+BzmQ6JvfinQ/I1g85pOFQeULaXo+/O
EuZRkfnPjbS2C3MUZVzv7Iymbj2aL718J85wonZPzyL2uCU+thkgOojeGMZ0aUVdWk1Zs/bIn+0J
k3cVg7SekHjPgJnU1aO7JJOVXPm48if5xzXlE8XQbJbrTxOEQmYhZNQRrpQrJfNFo2amsp9sVT9o
mObIw9JiWY9tXaLtlPC3twe7ENmcP4zCx8NREXybwNVoMa8aY4500MAAQ72SZ9vyxdKiY3DvhORu
99Xijl0ifUbfHMCbo+Hx1EVVyFjGr5AyhCA4DWF3+vi0z0igZjKVlKh6xLftHbrpIHGZGyNH3Llu
rcyIiSUZ//OohZrDiwaL9ObV+CYgqTRpsy6hLW7yz/RiHcS5hmL1vVfqlhUfRMR/H6N2ag8typ05
hOrOp2YrBxr6Hw2DiK8b75hqJQN0xjHveLFOVWn2fizPXkhlwTYU8s8Oxl2gJ0YoWdorD84q2xIF
ATPDlwEivt6ytxOl0gGZLNjRm9A6D+Kz78QRKpY/rb2VJWzGvGbqlAO4CA/FN/Hwlr16HKDsZ0oR
k43c6MztAUyb9Um+zh6kXU5sSR94alSFEJe5a3ESQzJqj8CLXHak0Wo1843iK16kbJtuRAc4cD+T
gJWzVgeS0uvNFE7dQwOIqJ89JNivY93XOziF2TfSUnQ3zfxZ2fIEjAVE9cDDhX+HU5ylK+oVFdgM
UXq34gf7aAa60us6nNmgq69tD7hXIXwbIBQ/B034936+8IeIMMWC8H4sfZq8ygxPkbh/D2c9LB1T
L2M6KWCv5966lb9djx+sp/tFpANsOL5UVEkX32I0CdfVSUphK/WPX5SZXwod7A28ESZJzh0O5cxs
+2AYwLxG47yWCSTJgJXO5+UVREhN9B3SqcDQ6UPeAxpl39HuJxH3PtfnJK90BWot8GdQExBP5pMt
7IGCH2Rz4ZadSJkxq3yGLwhgTgnN+IbI0QVZ/P73EYpi9X6cdFqZVSMwsy03fIjzSLQ4A+MEiJy/
IH+8d+IXxkTCnYCNGloXEGR1U5IEYfN4wvYkRQO0n2JyMFORXRc+nQ1iOJnoc3dQGVQcZ/6pBBKs
3RJQusXoTqdcltvqxPyyE9cAEAJjgziN14tXiiv+l21G0OwO6c14nkOYLB3ptTSlZobdPQXibuwl
NSgcBGldQHNXOhKT9wUy/YwOSQpT/Src6MATLA6nSskQQKj1OrtJiO1gpMkltTxIfIyXeYeKeKhT
cqGHY2U0LYnwuVfI2SdIYvmO+Ysqd703/b4b5SPehAf51bgb2v5h3lcRJA4yGXdLGMyWlWfar397
WZ1xfZfpEuZtqICEIdP3myEL21ttFwQEmkz2gakExrZDXOaGEFfhvriTvqsptv4ucZZdFITC7Z97
7CIeyfbaMyYd2ztRHkmSz+mKI6CgBcXUhPMJWr9pbOFs1eRQpmpsWerThGKoAsJOu+Kv9VEnmvd7
EnTqBBqD35vvhGmxkVeFToxVqTHfNO7rnnidbQv0hZKS4VMQjK5pZ8v5GThWX/EGgpastBxZacXL
wDULQ6wSwt7VdFKIVYXxb1CA3UC0swVOEoKszf6acE5tc55UDkSUBzSACxQ7MHwf/KPsJ2qkp53i
dhMR+4sQrFCY/jcWVGmn0sbVHt3SAQPCl7DVkGeliHrsArANUv68mm1BNWh3Qq5H9Lvvm6L0GLEg
WP4p43LjmtR+UuJCoZtaEDH2OvllIlbCEpz6/uQVmoHHEVRF+Kdt14YAe2zTfIql7kegDmmVMuq5
xAgCA8PaqonVD7Ly+vQjjvrvg4hFNL8DRIE+Ruc941XC5VbOTiYQFzVeJi/2lp/M27v/ZQslTYca
T4wCeXoTWNPoSIyaWEv8wSD+dZAXJJfUam2TcRl5G0fuhdJkahJrnOAgmXm55lsctEH/w91sKrg9
MDh1FBdtPZIaYQvhdRfvRaPtVPvUaFqvUd4/ie5df6uOTYMNe4foQhhqWw2RhVZfkYNsjnOox4lI
NwNCdEoTX8Focp5Q8hczrhNbjz1XkBf1uURQKeF+AFgdGKbhlxugf1/Hg1Ru5EBv4Vd1VLrQWEc1
9PGuxIcZNAR0Ms9UWcrbRpSq8AZ42ctfpb+01HOvH8vuSMRT8HGUA3zPxxOTUjO4xVEPBNM9qpj6
V1yYecicWM42P/jgGI5XwacKtnyoyavoxeqtUWghv4H7tuA32RDaKF0cL+Tty+N7paom7mZKkUv/
l0lpGcDhzkVJ5Qw55aN4ZbQ9TLJhSahX+OJQekvAFo4M9PgKOwqMBehn1qXkHGUBLerZ1z+oXVrM
EBtfSoaZlvCsAtRkyyEF/alqAI8sTgC2CLdCOY78WLwe9ZwzoAIv66zJBWVL0KUHlJ5oR4KrMhyj
DCdDT9C2Hm4jS58YREQR0bYl3eizf79DHvYMG9VTRyQsYrkVgGZs8jvsMbT4DNGSUXEOcliJc5Si
oLLD/e2ef4uTfBeoJqFMqp5bKS7l6SYP/qdiieFxjWx9HI7QC42G9pf6pQ9mCJLaKCp8opVZv7Ca
B8P1F2NAmS3B1QRUHdQnV0Bv/s5FI8u5cFgkeMb/rJNff1V+YHi0nAdNj2tTn3lwv9Ru9kK5JQmD
UNpaMiyVcaeR5JJ6jg6KPLJn8fmCvKu4LpSSdbZYqSpS3VabAf6NpR6ahYwddZwahXLDcE3I54Y3
CHxBbJxbj3+15w+d6sp+QmoVElJSLmP8juO0CV6ycbT0IpfsKZyvLDwjP/d72FNKCsRgfyCsCmxp
BCDmojgWfbSWQL9mTXP2QVHztWRLhlCcLRieDGVyAD3SeKfE1hqkIOHM/d/PZIO7/Oyjt8jJgyj6
QPzuIVknB+DVk8PZg3sG3yV1EevTFx3iBaKA0AASh8ABXpLVZmBj6gELGMr83H9/aiXJ2cKrHmuQ
C3iWANBkfchShPVmBKnb5tTh8L1hHE1M6pWH0xy7kTd79VgFdvPiVonQPj3mrXfoxiJsyyvHcS9Q
C0GlgWM6x1W1dP8bD3d6RarkRC4JJBhPTkNlHEI9fRce6goYHjS3XWxuSp+sFd3gsJWyAyN62g6N
u7dbOSCDiD11vdPoKZDsJF081sg3oE6BQAQvBquEe9WfHk1w9a/x5xg6hI1Tky4jq1amP4ZhSrxx
J/v3+7nd4BXBVm3obRnDuaI2Iqtjbzc3PDny2Ud8UrrwlcfHbw1SZIMh3yGYS6516eLBhe82RIdl
txEL50YbV0qinIbxy5kLJ13GFjVX7fCBAIlfD29VYQi5CUiWbVOY0GNlh2eH4VPsoMQpjAmWg0ni
uejsidJinAOw1wxjPSViKWOyibha7ny76niNeDVLzLovSqPAziWP9Xx8laAjppy4meeB0VTB3BnW
hGcydKQzdRoP4bokhDSkcURnNY3hrIhCGNoTLPospScMz8kkCPJdkTS+lJX3dEgRS65nIPkK5PkS
eqDI+F2kJw843UP817Fv5mN/y/vvuvx370i/V2HZ+EJ8iV20RTQCk222F2JgJhUni9bKZZO7PJ6C
+N+3Nfzh1yaqfR5XM58ZT4vfEng/WVXgkD38wtPECyEXihbfdwOLvJlHTYRjF+YuFmDiaUOeDNFu
n4GuID3SS5bppOXRiSqa3qek+ALgGYtqSWIJmnS9kGpFX67ywhyfvsX00vlM9ka2wr+tTvZHtCHt
3RhiPYTkHTxPXZR1u2XVFgqezQEQZzqZEnBKZN8fbz0WZCwtI3W8S9TThE7V83YxHPYs+AxtxKk8
mSFjJgfJqBNoGcYu1qvOOGKJ404lSxVWU/Giqjseg9Bex9NX8znwhZvoZiGYvmWRypK7DXDYRKVC
oVB2rN83aKP86TXTH/ZsKMpsprfQz0HAXBP2cNwgxbToP5T6t09slla6VfLFHMgtsGpqIcpolbap
nqUL/Mi6bJ5zzdfeEMH1tQdBK+317qCGwt1fgefjU16S1IOMXN6NB2V8qNbAmNk6rGBqesbSUOCC
YYv6LxGefVwsl8MYPcl4aO+lcbw8XssJE8qnRMuTF7YaJvbkHMCn3yjT+zUpXUG4ZuPMQu5Bh6UF
nVcUD8g3FddC4TxJ6ST/Wu7iMEB73wBLaphvgz7ZVKWE8L/bwhb4e1nMVOycVQsX+fwEE+k2ZXRS
5joh5/xDuxFYMweQCeIKzt1AOOEHy/bfUcsFIAIWwouq5U7Uh3LCh6+11HfLqH/HJ4I/r/oWuJq4
KtKr5gLHxMfmjz/OjV8zcC6jGB4i7uOr63gq+DIrMIdRpDA0KnrhKmmgzR+lAmE8BsE+wRObnMLY
pIMThCCLStoJJXe2cdE8fEkIUEJjDKHMIo+bq4U7SIS6pVa9Rcw2X/OELygRKhaa96TP5id9vz+h
rQdQvwKT/d12zakZgivvjBoDu+3qGqOIt4ghd3Yrrt8h3K/QFzgfDdYwoFENwSUUqfZFSn6Gxsj4
4okOH0zXREWq05S8mXkJoXACndfrLU+52HCPKZe367/Qt4FrWEUTXRWuqsrmkqamYzv1Xu/qGp4W
s76de+CwX36czg3v9kIypewn6DZLrP+hdf1K/wGJPDKqGGKaNB+Wl0ryffFS4vKhUbLpNR9khfn/
UJgWXzJvimN82ToXOqKKG6K6kE65UVCu9NxE/dUNxMWf8GmG+OlMtJHlIZ/dLocMhJgWiCRTdsTw
gu/EwrZWqMufc0mpNkGSq43eTCH/NWYrJiiD0UUegT82Z3uSSB2IytxQ5G2uHvCVTCvdtIWzy+1w
B+FUqgl1dw6RzLjZ6jYQUYgAvcMC2v1L+IljIJXkUbXf2AhqPlaPfQz7eJRXb2PnrTTkC1NzcNQ5
8M9JLmoMfjWE91wMkl0sjnt+NRd1l81CMu+vNqHrZw98/805HGXzHQHCaz55bGXba7paQ6C+03qt
c90B/+sN1MOLOBg62oIOc8rbNSiolAucwTg4qxKn6GlY6rgcv8T+jkm1GDFdWhpQOQw9lUTUdx2T
ZU5pv91e2SHRXFG8ymXqX7J5JqBWocFuMDVqy8wC/CBFDNuSVcfs7uPWdh92kwdih9xCAJEKWgr7
+eaU95lv4E5wxi0F436418JgbI28sIV9Pfm01Wvp6eGNWDR3ZExq2aqXyGVH65vP7nbuqrBLaorG
lpQnoABfvvrCz9BCrEMy64kPx50W4Mi0lGyog+X2pEH3TS92ffFHxuYaoBnPedB9tCOHrn905iY1
SPfCKGIXgkkLuTaF6wHVVoMxH7nEjTHo/XhIweQEU/pStQj+ZiKDTFIXHdFaAJ2akR0QnWQ+If20
hGwWZ7NI7ptrqAirV13PQRhBrOOEky0xcybIcqca+xCvbFL4GjSzJsMp07NfWVKnwKr9zWfU6gz+
Gz48nZEwDAsFhuEGqmiiICzx2tBZfbdlHL8Mjcv2Ln8T4hXZqnHQb3Qg+PPiLXyst5tKUO4jEUUX
OmTENuHi/bfQuWoYyXlZDQQ7oX/DK5OmuB9NRGYH6+nrJYBPXio1W7R1c8mVAH80qFJCMgXjKFL9
Xp3yCu/l02x2DdWQirmzPohiJoKAA72QY45dib8MMqPjKlzI7dv71D5AmEmSwwrm0yBSS0KCKy0L
YyZM6G6YtGwabUGOGyH0mEpHnnbNS4zrpgx2/y2EvZfZOkoTPogI/oDS3jUJ+2CGQ4um8ngSkIjl
mAytaj80VeMnSXzKQwd1R27fK87H6Zg5N3mzW9c93NCZViiUzaqHlrMQQOob4YrRLSwZTj2HH48P
e0Z0XbT5bmw90rT4pok1AV2QV0BGQihZRkl+hHoiO8NEJkpHsA/Ova29v3jXmnnVHHnPD3QabEC4
TlQNylDp3Hhx6zQYsZENhlUMLwsyidLX3N7pXJaMfcpP1lNoFbxrfNITSNOl4p74S2gtZYRh6Rcn
61DlmrX0iof19kkQ9lFiKPC5FxHVRLIK3o7ZRmzJsuvJtm3BtI6owz05jRjZ10w7d00nW2nKYcEX
EcdJO9sIh5Eveyb/slPmjSZ/vUwqc9zrGrR9nfW+Je+GjW0ZSi7CxwJIdSflrvHh6xoyuz3T1qnk
73KQbgDYSeq8JhypVjJsitOsK6/fL5khvBVGqriFLDbExhMCamcq9AIjMbnvmucv3Fauj0fLtQvq
O9NLybeAEWQiHAyCd83/tMigFr4weJBzbLhXPF9CXsuw+XLE7QcAcYL9qN6A3Ti+9AL0lFyhH0uR
KMpoQpF5TNYnchZbjCZ/AHokDvEzp0NZ+i8aL8G4r4XJ5WoBXseHQ9NQDnooKZwXsGX82rNQZgIM
3TJGlBGKlNUggB6MV7RbQG0Qzm9y+q5MI2ikojOnJjlntCWns6kDNaJc94Zxc7VTlxianLLSFhwN
O/sp39IGSBsBXNtHb6tLiVXDACQ1wzchzRMDfZWi7OlDnfeFaeg+3499w4faFpFQArRH51OXadln
i3CtNuBanCtfBm80C1y5JcbbyNiK76PNNAZecZuAwcQmdLHyNwun31chUCdE6QNGxESMZcb3U34X
7U16DZf1N4JEDfPFnlNfseTnYdnz4y1FF4OaqXECxUtSSwxg3nd0bPut8dd4pTsG2U40wbSVLmDd
/EKHTnEGOEZ6RPpLp9aRCggVgR5Xe1IgOEfG9rTOztil9CaTGEgEeyyGnre4Io27XftdeDWSw8wE
ormVMzcZRvRjOfFYBpDveTnucPeA/FLPu9+uGmJYUC0U4YmlVRw8IklZEf812YMnBzuM62frVD1g
h/A75HqWC3mndFMuwSzpsVwDrOQgkqPkqX5yEx8g5jzg64TbfaioNWoGbAKevbEhtDMph5ad23sP
EI8LUPaLj8hpuj1lL+0DMZsMyeB1c+wroljvu56ER34xFm4w7vsr+gi3UyZf6dC7Vel+MW/IcXzZ
xhIRuugqFCqQov2U5lU8uRGMYIF3O5WcSQaQjkMKFviy0YrgU8ZJeh8iqAZzgeoq8rQpZPhYICWN
IqAiI2LhqUMBEej30ckWCCEg+oahv3f+7cxxPAstwTLsvlj9YKKOEgeC5i9n0pbVQiSSUh7Rosqi
cSdfZSPiLJC4J3QxSysABOdokZ1Q/3sE7QqGbP8V+rpLiBjIEFfji+myrf+gcDDHWASpPNH5ckam
slKY+OckYQsbVgInTbw8mGmS/ciQhndnt4qnICrtNjIfARBx52ksxhH+nwTo04zEyEtw3Pw0iVbf
mRwp6p2PETUn9vQ+3Ezf+2KAQRwmcbkxtQHKeCDbIr7beqyoD8VYGrfEmgMHexkAji2IADX9HxWi
HyZ8l659ZQZF9sI1CYr4t8VpAgkdExrhe71KLQf0jsGoxSoiYkwP8C4CK6RZDiK1FkGs1ys8mi1l
/sGaKkZ4OzOAJc0lcqal6Hz8cPGHlWDRCmqKymm+lre6IydGrPbRwkYyCPWTEvcsUZYfNXmbB381
kAIaBe8n1LatRKwwh+6XCK2P9HfIsPfLETQObVoN8ATtyYAWqIPNhOCAYIcdm+SlFxwiUWUvsvDg
b+RmsgbXw27x4PEtn1RCU97eJV2rvES8dINdO/n14Qp8uwrvQCaM8gT6FHByPlYRNnm4tVCcdln5
woAts3weaCmC4w4HwUBa/Wf39qB9ekcXxC/CB6hgNDdIFbqrOz2awHonAvxUW7qVcqciRkGuEeV/
3sBjhx+i/hKRLx76TeB1dKkcZ6yZoBc2O0NVkQn7EqL5S4sdVcnEc8Ahpg2lGZAZ5j/UKaU8HVPH
zWc6wS/Y6wyRVHbnYpAzSDPVmI3VoekItufRYQc5mP3GyJi2jmZCFn9UR442YrTFz/Ua1q1bx7IV
G7zO8E8oMCtWayh9FM2NKiA1OXLmeweESytqBl58nIpXh+CHYhMbWn+60jBvceKvk0lE9pfwT1aB
paGw34G/uF3ZcPAUxVnoRewPaNve95nfOV0Y1givu0r3poDr0Zalu5W/sA65f7O6ZuU78DRbpfMm
2GMmTZQdDEVM3cZpyJGl0SlmgwvANol512fOtYGLiok1VLWu1mtfWdEs05r71Ml8MsmPlH8IVzwZ
69/FN83NPnDdbzNU0YxdUpSTxc73glCiXQafthRBAlz4rvBZfgHnT6MeKm0q/YvU9/WaY0rve53j
e7Wv2Zw8CAYMIYAgmxCDFF73VGoD8hebXlCwNHVK+xrBeW1JEcQRlGpKEAn+fhP+ytNpiuIas83+
M4NeCVcDNp0K5bdnJ64SwCsUoGW3pLTLxsd9AeTKCpEtXGmmpU6NXqIuiAbsIsFgzhQxeTs/qyEN
9ahXzE4LpGy/jqfQwG2IixRnYHTEecLbN5VCwc58XaLxn/fxdSD2mYH7WgR23UfIBI3UGAEya/8J
6pGUsCKU7n7H4PfOGez7GmIlS8pscH8ZunePbOdsbDHKJnEQ+nRLhMuscTczY+bOS0q3fYUtaFoV
5D8qFtgeVqkEtp9wu95gH1xdN6DtaYNQZCkYwsaAShQXe8//ODLh934dWDlKgsJo6sKqDomK1Y3S
BM01DC+QIKfoi0vVWvBjAllNPoDb4D2ft64e3ywo2yXgPu4oAxExJGFbcayLzgYczu7toO5/b8GZ
JVBBha/G1oEXf/wXzjlrizg4C7zxEYR6KjU0XTMWGFqprZVGOTnSPEaQr+P//tOmy6+S3HAmAj2j
tb3JQi8vSvCz+83WqNi8YfGqGbP/Y5MgC5MLhTkd3U0khsSSACtg7KXGHGoLhgSL//nOjP6Tn5pp
3owCFMBMZuNRZgwU6p91XVuCYt3lUWAmUxPUpanWgyn2sJIEn1qcFu6qPTgZuY/RXTTVvVbMM+DX
7JlbUrWcicwKKgTKlm73QIfhTA+OJbw9LOXH1Dwc1QtjBpXhXsrqXh9YqC2sNFaZwNxak5PbYZGI
QKQbhoSduz25S77aKv1zEJXbNXcEsbmeeAHJaGcXXEHyznwpApvdtQAeZqfoGAy5vxFhuYhxs4RB
9g2Wu0prdusY8XKn9nDJjCtav6odmU+MoP50pVMHNOrTcx4ccpblQmhjrz3D3EyFByQi1XC7X3dY
zp1BYANaUaEoec73nONBGA2A52rcU/rPwS1Y9j0zBb9qG/3reRwbNmPvUmo4a2lUGdCv+9WeuKvr
AN0V9ZjXnqiIspvmsPx3EEjg4v2Dxew81aLqN+NZnhoYJyB9yJah1yuobo3S2NBt0q0fKuMSQf5k
rX2Fj+grxcdiVmuXXBFkxTDDkxClwxGkBnuxiiC2FZmLhC5qXNY12ukjgwH+8Yhgbu9NXfnJP/e5
uPfOJF3vUMt/oHtBWAA6+JhCoTIJS7TX5KSq6RtCovjBNbb7jfqUUmUUaMfgfyHls+vgYe9RqPB0
oKIOYZxFPfkRCuia7QhMJ+3UEXlpji0Qv9QliFbjA28vM8hVQVcOJ0beYqpjz0kr+oaCaviam0Jh
9xublhiaOfORMEFOR2PtkSWDgND1fWjgEY/gx2loeQmufrbOrTDofWjU69+Oq2Z0fKziKhsWuSXf
WJ7ECZHrl9pR109kuS8qRizZgAMVUSRMs7hzwVca2ToIctfkHjanpPDvR0G9alyFwx22RADnaS+9
iJg7UYcMCVpcbZqSnK+abPEhtjSpCLGgOSmOUNzYqLgbWpYhOqKjT9UiApfxdZko8gczblpvOn0g
Y8MGr2VJGdd9vsRfLz7wTSNUNfyCqX9vUVZpSHQQN8MfvLxDbTH7BZJouPyXyDfHp4MXjRTepNkw
qAvUXB5BUFZPcQpxBQ4dZmf/VnjLfjdt2LSgZEIZgD2kX+Rbl6F59sg+FXdzCOWCMP+BilVBCw9S
hpYdi697EclTOecVZuLhYnvacZnY95e5r/EZBf/1m6IWb8a+O7LKbkgtD01n/EOXcUbayy8w2dsp
yWHt+CrnpRdWh94t5FJriwb8SL5Yaj3gOmaNMrxBQDCjTOkL6Py+CJh+sKwYCsoqBiQQGnGVGVQq
JvskPCN40q+73v7gfO+6OTsx0lbqPdqtGaxlbFvHe0jZfoFrMNi5UEWqhzx8WtzdaGGFi5F7XPBg
4NVMb6Vgs8bg2lFLr0ws3Bx0kob5Tod97Mm5FahTEVx1bpSnAJLJsoxFaPbDfB5/r4hSuGFIvzQT
patrYEeI9jkEW4DWP2kHru1b+GI9AoCMczny0SxrMJSmWE6BsuI44C6UUlKGgCE2HLugYZ5hBWaN
+QFu6R7wDUQ8YLSMF99zyS9cR9BYOPN7gMAZTmnKebWORMx1cFasdWn7Dt+3Prkv0dJUCTX1J4OC
jRxgTAaPhDqWPm0B/3noVftAXAk8irAqwTRIIgn5goDE9Me9LOf+FHC/3UATayIw3twPnvElk+OX
jZAtRsKpVW0f+kjFTOhu9Vr3I18hpQir586f8ssTN9zQRat5Hc6S5lq6Laq8qc/rGpxzvMLk6nKq
8jBtuvjoeAbEKJSgRVSMomA4zv4TrU/ELDKX1/cfN/SMWoUD+KJVDXAEGORD1t3LAOV/e5rjbVkO
mg0P+qft+7u1d7ktEkjFeLOI+qYK+a0j38vhvkuMDsggzbqtic/5irNcE+q1Vro8qL5TF753B4I8
wN5h/KU8SG1ZaWs1oH6LhsQfv9qxbvPFFy9S0SHICwHESJOS6l+GaR2Ugf9n0hRLnTRBDPY9DM2H
IM2OV2xuZ3TRjsgetAaiVQYa9I781k5/mRSigQ6W8xS4hf6wtdUWOplV1jbB/Uj14b8K8xm18rAx
gHVF4pxnY1f+OvVjqEcjapWyP2NxW1uXB6xAMPc8U6vAcumUJ3sV07QKdJBJx9oZjSw7dEYsEkOp
IOWTJmIqGEhXDlWZFiGLQVGTl9lCkOi0lkldWCLuUr1x1relAq0q143U76BTOyD8shmdSAj1voyx
x6XjGB5qH4lGGttkl07Jp3ggyhVMiD3V0EykZWzHp7X7VhTdjSGyLytFznJSsCZ56OmD4LDvFBG6
Ro2CFBcWF9b/M8D76bKiEI/YFNKKagSNZjnQCqE6BRPvJfxJ8IlddvuY7bwCiusKrU9ViHVoJhuI
7Q/3PAeuSYiO0Zs3cXNyKF7X2jT9He8v55ZAdPC11OTDm2PWVMVApPPy/76Kn924/NX0IpQs22lX
QBqW5U/UjhMheGWlQoH/VlgDQD9Z/eitJ/a1sJO5xuLg9CuI/UcEPY0HfbbF5DNlZzpkECLmERjZ
pFxA4CCgTrBmJWlsXfQckRVidfUBRtKjNIT+OSHfgx11cQbyS22VRJ/W404INw+dBlShm/PV9PeC
l+Wh9ZknsJyDfUiZx6fXp5u9K3G3CdxtugiA30DaNn4NNFv0g6ukbyAexgfxQaoAaGQwi3L6zniB
T2jsQUi4U+poRXSmEPBE/KSmh8ebFtT/K9wOqabpjaRWhUi1KDfDKtD3K6ayo/r+qjxoehVBaxfw
D4LTeU7NKi3HXFpXS6iDpUWgzTGvp+/CilERQKI0/5cN3CQNZXAZWFtP/lfVv+GdhUWRtFq+2YYU
djku4e7bTEGaAcyFpIm6vfKu3/++/kXAlOVXoD/dJwgdND0X5SFedDQfTs51lborKHI/v+98z+Eu
tDytPgiI73tWW+kKUNQXl9/48Z1tvURMvHLSwEAhc6SmwWMTgd0YEeNb7+ZGopaokYkefkd4AqY6
2n5sRRtH/Cl/r28kUzaMKn+vp8wRTDdajqGQbqPuggcBjt5nRcH/DdP6gYVaiZpd5yTKYHLFiqip
cObPc+uGSPSmQiUAo6BX9FORqdprelvOnU1TaeDbmmHiNOQtxQ+QhXk2F72LurFk+QBQBzofXIrq
6HnN7uqnunq9C8XMO/tlZWqYaltJpHUKBdlhWoSlijrUxIxKuW6GNYUw4DrlXgNyFp/0eb8iE2Gk
6FFlh18FVo1hbKshyRNV1UmqM94HMm7kJydGwXQp2MFrRLMeUfNywQb9YG28ZZRA/d/v+NQ3Vdby
bSr3yRJByk3kDGMDwTdzr06BdCFEgii43cnP5MtERhoDqTjN8wxYSAzZiw3qY3Kp5EWzytztv1lE
KA5jD6DcbImGB896R+MUjG8fHUOX8sL5AdJ8TJUc7MmKGOS8j2vSrZf2Eqw7L7H21BU+6vBrE+do
OcNNOz6gyONdFeaui0R70XC/l2Pi00TxTrAmmHA/mn7M8QHEEcFoAQiP6xwfk86JiHVTa1NC7EG9
6Ta6r6rBhrlwsLx3wYl3952Mbx4V8yWyCBZx4rlnVDpwV+WKtb614SS8H0clJCVozO5VZ4ryTsny
G7Z/MxKKQoOM9oOicsZa9OjyAP6V9hH4QisVFZp9DXYlRUHjt8ENkHrkT0/QWGsaTy460LAoYHNb
/inPiM86T+ftRLdrTuBrik4Y2ehJ37isgLhjxclAuJRjFkChgJCEHwaQxJ8vulietegVJGBFsbxW
osG1yzmzxHluKocWWCQ6X7sUNSJAdf5HCd40iL+sSf8GTvjyAIC1dR1lWveLb+0ILwmQXNTC8TKM
Ih4SRiQuACT54Jahi1fsOqlNIV0AxTjBuH8wXnoojWrDtKyMwfCy3vd063YKYPD9lWoREIMadOi+
rGGleXzLg3VwS+Vw5rg8T/ceqqt0D/+MHNp5YngCcheMxOqCmHyXDKNHGSoU0jvonIzenaLVND1X
zp5hveLA3Y3a/lZuUnJRdMKskC3TaBB3HY1NF3qX2FXuGtDskOpCPl+Euv7U6+0AKpAGFm37YRvt
BdSx9pqvG3L1DtZ11jktyJv2/PkIxq0FysFjGDP/X/gcg3SChm99UAOdCDkjbH8lVBXSEtsg7Vq/
bu+wypBt2y6DO1syUbdBgUa913sFVyfUdaSRIkD+q/txAShOAVrp9mSP/pjyQcVvG0gUUemKp5wY
WI8kNa+66kTv/E1DkbcyXb9sChG9mY+UBJTABl1BSOJ0tNa+IaiBmuoAK9xPJenvkcJ3NZZB3x6W
+I7BMTTjzW6BoEv97bjR4RHc5KZkINxUXANuDZhDndNhvnTFCQ8nXtM1a16hu6S/9K4x8Wv1m4Rw
uzWCZsZDu9ZYRSe8kYpzPfRIzPkNAsBeaN0eCrsLMLrBQFWWSk3Hac2RorOT+InDBEUXVsZmAstU
UD+pC/8KGm4CpN3qd/g/ucZk3/U63Tt3m9biwLdwBdo8/SzUO95dIxmrekaZoqOGRWkdoj5/EMzu
7aETm8WiJL4wlmCauZGBy7ne6alxOWGf3UdOQ+WXnU6EdlC8CWRJXi9j3wxDsiYEoyB/clZa6BmI
nmKTliRv9PSX8S7QFCpM2PlgJntX2sv9MrnTDX/jLwCJ+0WfUh7A5wLcAqNyLXbAB2IGn0w2+mgT
SVuvsOH9q7zD5K9G1Zn46I0ujLpi2zvunjmUxrgy13pYTUh90TQFKy8bzQFzPlTv2o5tNyLYBIqv
ZFsHnCHYkkSEgxYWtJNBW9SiW80/IDAbZ03m2zslku1s9X7kc5z4ReFnV5KEoe0UAoDYN6xGA99I
CbhbwbbBQjgwPL5SSmzHtDkkOwYKfFn63f9hL6nzWYSNUKUw0TgjsWB385Cosy4XJJ1OhpczvfaG
alFjfA2cXUWHoX9Niq2tAjKf6PNtzFDhWgaClLsuWWwoHubAlmxEyThVUwHfdzJBx46sxlX8XZri
bmUthHY+DpyAfiVOKPxBMn+TUf/WARYRG1lg1aIt5A9U7m54MV3tRWf58y+1BLUJLk40e/X5OgFM
9OsRWtzdIA+ZhwKnJCEQy5pT4j0ivgZaHShxue80mnvrPyKNBk2RdKnu5FVqjpKAoghoHGEvQz2L
OeIEcSb2oUehI68+//ZxIFuXlZu96jjI38l2fembr2bAhgpHBecCsas/R8Ic0Mxy8BHsShFMA16v
mfwuy3LZqoOq2wBrMsNangiD2XAv8UMyTc1elDlx1M27L3DxcVnO/+oiTtk7pjt9DRJnl8cpey6o
vy6HBF9ZXf9vaD1/6fbsxVJI8Ojtf1+wPMLAG3YwdMLOlDbNSWaYxwAHKxg+Ja9djKCrPOOG5amQ
eVzN8WhgVTgZJiTnZk1EmR7hYZ1VrpKqWcd0ZintSIJNUZt3BsayMbGrOqslw6AfO/q5pgmzJSnc
Lz8Ll58Sm6FxWgGVaWvMFxmcFrx/yvzUdVFJKJVI0svmJ1/5a6lmWnG/+eRALQgTpsm6/DYYbnWD
pv8xgMpYcPg9tE3nTYUomuXfHQ7CsWV4LBSn5ZzMiMThT7I/nC3XSsxkJoXUcjiDHW5CPoHLJaxv
0L9z1YJ19oGkyUkKl7kZ4gdt0+IuTSsYDRM1bnrVVXNByMMdImmwsZ2ECKsqSgKWXR2rt3arvFI6
tx8pSafZq7153RxhMrJ4TQ5mvolix7rQlaM1Gal1/vAcC9npxwT5A/86mZjEwNZFuY8tAD+TYGzz
I+p7nl7Y5+2Yt4z5n93Ys1CP97xYWFfT5xc3krfitia8bmtqUMBem4zotaOdBPbEr2P3Zw1jYEWp
FB3vrN40UvyYXpZoUhPFoCb9UgP9jeSi7whWFRwgVQz++L7NbX9BrYzo6SVdO07+Fghq9kazp1k9
kfreR+H1D885upxllY3vCu6ueyzT+En5PWHF8TyoeMwnUKpHsCXOaw5QlHLG+IxHC0oaOerj5viw
bSCKbF8uWczJaFH4cC71lQa9i5s7tQb35jccsZHz7rKBkj9wiL19fdzd83MCFYsQ4aeTa8w+/Weo
vx3TU/xi8YYbmcvSsMM+/KvrqyH70Qtzn79+ed6ZGCDokDrFyalD53U314yPQR9KUloazolNMoWy
EzvAQU3eoxL7Q5Sb2QUlsQReO1hMLvwdT7yFj+OZHJR5sveMqIDolVT3STQwAjJwgKhQtHRyJUUj
XcjMxvkH3394/x3touScrWJCtVucjuwjEU0TTugYg/0n5iZ31fBmIjFBtM0H4m76MPWhTyN8ag3G
ZW/bhtxTcv3pKuy+lMPWuCyjcKPfVLrV+PHf2mTN58u9/9lfjx7nKAQywvnEDZAMDKmpgM47f3ys
mqXCytrdDEbbKSUvziHW5N83lV61GBJJ5xVrrZslgqe3bltwTgOK/pzhEPE/RXRhXjdfpu5KAq5K
+RYFDz2p9C8B6oRQrniTjTF5DCK7ARAmbIQhGsWVIYf7Rjv//v3rhh92opEHbnhiZZ1Jsyjot7Hh
uzxZa/gmEpt5Bk1VT+H+yj5ChtKLxiJDxrxI7wWs9EcO4qscbt/ESV3EkUmiLOGzzUyq3OZMD4dQ
n8MO3qgZ4C+NDKydu70zjV4NmIIkiNaL2Qkf8AornrVSLMO+ZwxxBZi/VclyKmEzvK4nryV0Z7qw
vazaWnHV3ItsGgtox41nZqIFKkdpc2sIMGLytAwXnqbyU8Sv3u3uBepRg7Qt8T3JjlIV2dy54hje
693OY3LR/tdcnqKqgonTZXvx3Pl9kFFID3AFZApSJhjIdsHXRqtj9beCK/58kwUR1O7PdlkOhu+T
4ScqM0itICWShXOvDPQppLeGhc9nEgfWL2pnEG5FnuCJzE0Sd+ecNqIzVrdNRU9S6VNnT1iyhZd1
ktw/Qd0AU5d5uuGJh0X9Cz4mJvIb0YawdEesfMjMCAzLGpObo8SSnuH+5Wc0Y6UzexIsFXemlcaO
ZGRFH8qXQgWR9ohhmvf+k3xbzo/gka6pgfc63hRJRmjhCzWWYKfy1S+SUtxWhNT3c0BlXlP9b/Eg
iK25LRi7Wefz4YJ15s/EyOp+9B3PtKFQ/8rCUCLl028NBXiMcnVGXUI9sNguhFtJCZoP2HHta/CX
+1RF4qj4Qv+A98BTSi2SiLziR/lQAMjJPquZ9I3vPD3q50tUAMR54FcNy26GkjKVe+eqmxAJdsm/
WWhEhGJ1u8J0v2J4lXjYUIKjltMQQuvFlhSMdUf7d+UayI7KFMyO7O04LZxucOK8QntEurRNhpQM
0UApV67xfh5q45TYcPb6p7hQymJAUmEsQsiQQDH0J8dIABjgP8Y+3cMpvK/vNHQQlmHzAZlhWmJy
35C3USYtwmJ22i5HwvukMaRW2ssawWk4HpRsuph80rkgXZuJ7usEzvWr8Xaf5guFh6X13NbnAITN
sOllgkaqjAKImjd54dydy6cQBRZSPy+hXhQfFzMcWjo+D6L84B54woLDpM5EL3Sdbky4tL1s5b1+
P/10cZEWAIyvi8Yfh+XJ0kYvfyzKA6PD1CHhYoLc2I9zO2Gwd1D4t3YyTZ8JSJqsdfo9UoqtOatB
eXHeUPJHOvbynaBtvswexc3QXvJrHZZmCIwc4yeNfRDC4k5aTj1rbaUYZ6yBfY9tUHJrl0HPWx0s
GfNjdUYGERwMiXaFHrFDOrRyrqyrXXK0JzJZtfGlvAOafyfI2HIcdH6uZyqqkswj6zdwdpkY5TTg
8olJpMMwaWnjdIx2UvS6g6a1fnX6cVXbXOXMS69qV7UfiNz/lrdTBHgexeUhWunfLwopcMO1ylNh
U4Ff6KxBoL3t/Q9utUJKCCMjlAfInhWLOfXMu6gGGoJvFKLz9xzdLo00EDjcjck8tEtlo3kcj4sm
+oRMgLbCEF6keYrhLN/8tRWlNiryDrzRSNFvx+45B+4892JoC9tDGxc3eCIVqJSaYNd8Qdxipy/f
Krv0/5oEMZrfAhXLP78o8jmQikm6SNfnJBuWcQbRURQJcbn/9YnLVGLuMCbG83fIm8qW9cgXoYWs
bUxQh4M9Px7P5kL5NpqL8vSH9jvLj9fsfqhFK5/IWXcpt+IuEGeMHSD83UMIWzVlhb6Yoe3C9lJn
R5JGivH8NXwnDWKXTXFaFjNrDfrjpPceJ0C8NgmHqhg+O0A4yH+ow5w6TbsbPfWONLbgTBynDMJh
29hnGOy3uvrgmbJXEB+DueRCb3b8Tk6RFGWVosNoXJ1ULkAXGvgnuW+x4eICIzcksYjt+qJVt50A
nEpiDpUt/usEmHv4TNvOLhCoEgIl0SzLLrDyFHB5eB1k0S5GhefpgUxebk10jwuYHbWeFuf1g2ak
0lzedvQqHKBll6PUGZ7P7hL1tb02TG/jMqkS+HyzmyJB6Q0pJ2WWp4jxyX9tG5D6psXvvHN9E2Qu
sGTSoOHU4DNK8gryj5tlb504oVCq2nhdmhmPyGFRzDiBDe134Ba67KAOBxRMDNuHWd3VG1ePKaEl
EatuCHq3iq3BopAJRlCGbDadRcLxd4brz2jYj4+QCrBfSHWsBdPWyo/NzHt5hQL6wILg2oNW3oqb
kfM+b9JdgM/gURCbUa40sh4QipVQalkKPREmp1p2EEasmoOFfw+5oCphxXsQZIKKz7+rx+8G7SJN
8Etrt92n/S8d1PD+Bxv3krhaUJiYKbj6z5e75ZpV28Di5fkfdBSrOqrsc5Endgk0yxbxXimuhBp/
P+nuMyeJVqbcue17lFDGv86i9G6+e9vyiUz9FkSXnESysvVvO6+stKRyFLN54No92W9gGgtzR4Rk
m28pmZ0orCMYy88JzelusNg2ejddQzx0drsidJOwT7J213fktdDc7QiPbd7ZC7NDfYflfBaVgtUR
wBH8jzSAplUuXCxjsFTw+6vrYhLQcjONfNl27Um+6BYVkA18vY2lh/09rUU9yP/JF5pkFXP3UfiW
RWglF/9D3t39y3thfqTyEQvmiOZp1DrZHfbzAfCjvHtw8b/xVleMbiqgqPvbhZ7taASj3fNLN4zD
qeFghj+lbf1crVufVt4ilNF2lbFvEWNj8V7HsbioSoATg+sZLB9XsGvvWnNvPkJdUnYcWks9Yfc6
zCa29TFCddl1Xwjp6B/xHxcE4X8zz6Wj5oCf5ma3/2aKAQpC+Mdho9H9qqj/8jCyxlHT+omADM1Z
oi1JF4zuvQiLGVDtFMNquUZWxpEOoEvLG56tkn5zd+9bqu/6kfDae2IaZ7nKrfVaeRIrcrhPc9tc
mi2nZwT6qt+mB/t9cgR77k7J0VMIx1kkOKfQMHxqF/s3mVOYHp9Wrw2E/lqO5q5OMhEUMoh7Erhl
8OtIRlcRos9+HOOrYGRd1NWgswqb2OFotnE+CY1bKGZ9MzgRe4OqoEExVX1JBPWa9uUJrOX84rO1
62j9gx+eorJAXj0zwZB2QeajwZFAfGxL4BewvFqlu2DG7n1JPmmVop7hFwG90ZHtg559NuTrBXO9
nfkzdmuVHvN7ao1+6WmBeGJLacRfvzgZBOEZC5qjivYwnMoqd9IwjoAS55n9ccZ2KGAqqHrB15xm
ucSSxbHEQ20S2V0fFr2i4PwMNJ/Otod8rjIGmnjZboP6I1YKy0CR5EGqCIQVJL7Y5HKiBDM+Pt8J
mEj6buCoK7L7ql/jqQwbO3T2C+ZGRUDuMA6y1P3Wv3YJHScbdCtuwYs4fb4mA0v6GKBaKECq/gJF
Li2v9dBtD7nMqFirDJ/zupYhs9V3mKDO+F8hEtNbAzBSRc5ZVqVj/GY8Jaz9VIDV2mOOpeM0stHt
QX1vZcQOF9rzG8SZe6paiKDQPJNHWT8qyw3w1O12T1Yt82Pp/H3pmGRMfqZWquMBrgcsXz7sSw/I
x/ZAwMgsMfRgduty9Z6fk+l942+FEqdgZoX82flQriEV9rMbxC3zdVNDGYCJ0NnzkSwR/deTQ9Hq
6ruB3NVPN+Sif/KKThK0vygcZtBWNFA8E97qxJTFcSLajq5NuwgUClAYr4o1a8cH1Gcu+ZPFMzwZ
JFT12m9aFtk8PuIEblawYTXW4G3qk31vrcqxOipv5ubRw3BHWjy7LuZhAFoi3Ttk7pzk2SDgjUK6
lGrfwzNxbsvBM3izm63okC5guFWxMCzjy7/9VxyFevrygY3++cC8w3rvPmrUEQvEc9MYBtXT0pnk
DxdrUvkTYcxUdGsLSDSvgGt9Wu7A/rxzgEns8+vLY6BeaZoAPNNmbZlJqKsgwvL0Rlc7fphg2/B7
qLSpjllJS9L6AdqGX93ixjs19xU8+i0/qqqKrQSVKC6gkLQ+4+ygyyLGIJFVJksXHtOqqBS5Jblv
7DoKRse2xFiLHmmXuAGYXHFzj2k/1GOYx2IB429DJDpcOHpC2NvnXI2Svs6U6JUbylODFvoIq/Z4
BtszowfDplDLAZr1FzOyYyLfqxIzz4+kidw7+izNs/Xmgr9dko8xBOD9Kgu3OXGzYlrfQyO5HvFS
XBkC4eQkAmuF+H0RmXAyVLRXzBHA7MdxRK+oU/AqZ2ZAIRhxHL8P9/oykYtwEznfMo9gFi1h/MGS
+WYlUr4z4msKKd0/b1h1g3MFJuoZ1HO1wq34v8QDxE3bZc5s2R1xHk/7kJANC/AjwG5jUZVjb+M4
0tr4Y4LBl9Ck1Or+PcUfzVWbWn1JqK2bHbu5J+V7lfxwKsJeMj/Z01622Z0bgrQ1QDBvkGM8Cxjy
1HymVoCFZGRwjUli2QCb4ER0nuy0CBOYAV9YyNo/VbF7aQTXyp+HqCTYP+1vmlWqW+5MVaQFzyzW
tVsY9x484IIXBkotQBkHniXrGRv3NWJKXQQnm2WYdbjclvTNzWx+0MCog1g24DL2KZmJ/vzOy6Gf
mSLWS7PV+vVt6WxiqPOieUz53JbgKi2BHEZkAV3oS6piwfU1LFi3UUbOVeqURkr4xvgS58WL2Jlt
upIcxv2/opK8QcUO7aVuOB/rZ7jTGGzwcTGFRlKSQswUqHncauYmG62J5xHC0BbEvniCA4mqinNA
xaTixQj+qoIqKAI8JTFrLibh99pf7lIxhzZ/ovjqcrysRxzyT/PYHDhJgQXJmq13AlIMgRM6KUhf
KCZu6cCHxGxMCPnHDpvX2dyNxcnaqw6p8x+OYtPjKVZolBTjYJah2BZLZB2Fj1gM4/o3Hygo0tpB
Lo5gcAvociTbhc22bEyeWwSYhUiXRQLttFey7S0I/40/nO74GhrB9+84QSWTh0UQ8PUWZII0y5fQ
BpMI9fsBScE/T6TmEgRy1EObPDV5jYozM2VSZy5vKB7EUBxGlhFDLZt/5M7C4u4zdB6rByg4YCGG
oC1Le7Qpnd5Qp3NBPQaVhA3UYjPSvS5VNqIDE/6IsdYW5l3fJxMuWccgBJQSd6Gx2DrhvFwrxiRE
4hTQ3wBwDfiGqh6KgJta0AOymlLbu/ksOUg6Qhs3f5oZYmyq/8+IxcxQ7PnTBssjq9N+X/hdjPf+
5eqAdIiXDmDZWb+PvxS/cGPhR5lvDzYMVzS40KcwW3SDxW46XE5Lt3OHkvyiST2v+ZEjRJiRkphk
2phwoXSQ/GeXAFgkUw6N4Eupddy7DLprj4Os8/E+bZEjgCfoEKqK+uX/zyLhtxpS3+XeACT090VH
U6RZkQnegs2Ncu5KZJDQl6dSaWPhbVBYBGTOLgg5O63Ko+gWI2KicvSytw6jYN5YQyTHdcjLDxYX
MpUVwV/RZ52PC8Ywt13rxlKx8pj6ork1UT9Tjj36aqPte90zYpTttErHPilnI9rhOvHojasnshIq
J+ZU09Hbup5ga/E60U7mVOl5rNyE7k4k1A4BGp5/+8r06GlR2GbmWQ6z3FYwRWsD/AMTKrwGsb2G
u662F1DfTNn5LQYZgpGjiQDyJ/mXqZDxzb06x/JxzNSFvkqdABd4Yv0I5gDMOO6F11bf7GlLFp7d
AmXq4KFfNQXyLpErSrdC9PIwDjEbBDVJ/wB0BfXEhRcjf31cdlSY6k3qdi225l92Gt1L78VIojri
frjVyX+XixB0HUMNxas1dUzPIeZmn5rKI/oYRFGzu/2vhzK8eAVKdDwQd6NvTjI/U7jak4yolyHo
yUN9YDgej7zEYInA0Pay0G0gC/2S0zt3Vy00vxhLNJg1k46b9Oh663EYucbeSIV6qereL+RQR7t+
EKyl/wxPOR6B3FAswOYLxKIsmOnEYkzenROxFr9L4JxUchocp+/T/sv+RHenyCpSet9HoMQ4mNwa
pc8A9hQoCzaeWEL4k+um7sh1jJ7Y4q6vjArRvy+NN0S4OZmUkYTL7JaWbwzVh2Kf2pr4ZiDRdlV0
f3ox48fnViAG8EBU0d5e5Yn0jOoJMbf+YaucFHkQVyasJc1queyPxDTTcpbzhpZ7O4KYARUjgJs1
4eSZOYhOB7z5TovtfYWiPedMkQAFIkE7ozLgEYPWyfO3pKn+6rx7RZ7aqtUYZyOEWVdqgTo94zCt
ro7xvbiP08B411Z4ne4aARd+xMVnbje0drITfglJk9eF+zjXgMDWZ31n9DWPf/Y8ABWOcjSe6uJR
DSiZmmmdifzuIfPDSENRL6I0abjNEEZm3XxI5GWBndPTonkSTBppbjtcsWQ5XZvmrrxdLdgWjVUX
XfQjB3O9mmxeEH3oW3le7mTfQLmmsywBnqAZRFKEjTnC0KrEw3PqdNv+no8PI2nRh/TvWcpLwBbH
gnGahNV932ipVkUOuF9PYgPrHZSS/+VixgDwKuV63oztbczTtjb77/lmzPIncaDf4uR8wgrdOKlc
YMPZd/cQb9Otpji5IyqSHVqaiHHecq3gvrGFZhRTijbU3ByEU363920BX8KuLteaFDzp+kIf7CQ+
OBH7mrYYfgAvK3YW2JXujRUzP3Z+C4Bk3P5KMEXJZxf4+ZgN3apgol0sJ8kFrpzP+0ozQfVTQK9Z
5aRoprA/tszVbx5/bTyARt0yc4HOPdAGrMqWwKAE5fvLaycpauXwcKt6b+lhk83+h1s9BBg9Zt2F
3OL6iz+F8HrUrCapxqLlqeDa8BfVT16dB9U2z0lvPliwwz9w0QcKpP8FAosc2J96h70SyH/H2Vc1
h8D2y8t/x7CAsz0qpO68RoJj97t7To5e3/VlNFBajlCTWwMssDF71fIJzjq4TZ6llwNIyTC5/NVd
8r0GBc6YFO3q4WcTjkRIDQBByHvRvw3/g9cO6kWogLA0IJgf8AkfbT8kh2QfptwFdTVVwTxnEoP2
421n9qlbfcqVWuhNFW9QMem4Or4OKk+pxpTsD1owuwruC5ASXe2ppxvqZnu2JdRFan46q3W8yUNZ
i7OzPX2u5io1uA0QyN6wioNNQpv8Uh4xT7Psmt1D7PqZOxjbmrs/kDsYRtVflpq+lebWn+l6RDQp
cu2lKaiW+rGkxpopDSHhmYz1PzSsd20fXfbqI3wpT6xw7stTRhysJWSWPX/DyuVdkm6Q8o6PyYlv
DiihDSPEtU/5H3ghWLj4huLqfFSlWjUZqxoFSuxfCDNjZRfXRaKgqxurRlq4JwDLzX2m7sJUKI8y
tm+kXGdaXojdgyr6skZB0roN+FdAhMzJ0ogGEkC7+ZCn25NWPrtoWndIGQBfINutMvgGuxzUhoWr
KDBk98zSUb9B3DqBtpCZOKpb/14CwzcvtZ/AjEpv0R62iNCplPkv4E3y9c4IkJFWHySQ21TUuE2X
Ei8bv9kINLteemorSXsbRjF8Yo89OfPcVDu9irZtBoygMBQU4z9X1jCaJimXwXOoUrMvOOY9SN4W
yQsiroueHA1xwf2Jmc7oYPAi0iWt/TOOoCGHB81ubNgSUglms49ztikMhgK7vEwkXyjVzrV3Kauu
VE+z0JpJrqlX0m4rBrP12bb0LO7fPG2thx14vGMKQCpB+ay6zkOrw31nC+UsfNs8uj0yFgL8uQF5
ihUa9hXmawH+foFwA+HVljI3OWFA9pAdith1NsAZWIBAlxAsCWGrinc+50rXSCQ67CUBxuGxZV+P
ihiEw9DHw64Svk8uhvIQCQrz8/wUkJw/BkcwYc7qTDbj6Ft7yL4I3XRTYr74YaEys2M8pC2MKen4
cngKkSRGT8s+rfxjiZfB2dJ8pDLvZa+bNsgiV7uBuyG1npwFgF+de3O+gWUKb+/4BtR5ROU1adp4
2zWN5HZhDbZ1YNtK4VHXMvYcvJkv1agTqv8oxw85nea1g8uMjE0eEK69SQeAVBiJKpBa/mJq5Cle
QJpZGpgvp5clsRlZkoAt+I5DcJVpHooQfpQoIAr5ya3YVrtNSC8ikQfOI3mj3gTvi7z4EvsQJrwT
mLYuRm0Klm0xty6n+WADwXHLj8dBGbyeWVm1Wmqn8rdddnrJZk1RqBOwQuz4gODlkw9b/IlE0qJP
gd9N///Nb5O9blRGf0Mav3y1sAjdOB+7fSnSicVyeQLKVojM/yToTaFjZToZQTp2Z28StgCprKs2
FLOQ9Zxz9s9IrM3ZJIXcvbcKLaEHJbmW3mB3rz5InTBHsS7nsJUyQovGl6tXs/PYntEjyFRe80cc
yKNq+XCYZAYiNPCrMRsrvNQMksgjXuCd9ICU07RAtaYr8bIkMzIZWk3QuyvLuwjA6RbshWsS8xV/
9t3pEJpNiK9wR8vDUEt02UzZAFuGildFDAE7c6YToSb/CsBU/0dngrV8WH6QmvoazE1cCVm0DfMr
Xn2IZjvSTNqRJGpA+Ihk12fy6SFBudCYOlnXGDfQzauTGHg+6iQkOYFoLLnYwgUUtuwd+W11DG0p
bpLcOuV9inujpNKJ3ur927cvj9eY9jZeT7Urd6B3ey6yb3/VucxKy2SRhZi3DC+iIkvwfOaOe+FW
mWw9/w4naIe5tA18iJwxehpxEeWs3fpEmlFN67qKMxsgGllPHtbeNHhZAKpPAaMDMthKPaDMghOI
DpHOz8grHzS5olLvsc4OfeK8I8r0uXxoSWG7Yf1hKTXihZ0CGSzWTVWgfRPSYWp34F+vhPoMEgzS
BS8Jt2TfSPvI+IBip7ucnASEtJSU9JzBi+w0YWMJk0XLv5GqbfsI8JtxovbxXTWXHNzjcin4yFsu
u4ar3IXXRjsoIqiWplH3R2CJkIMDcKkGX/6Hcl1WswB1TZtfpT/youU7JkoI24wbAJZHK9R3unR+
tIH3Uyr/IDdp6tiPHfFlkUtNuy3ZIIzRXxPt/NFWIVDwNARezyCg6H5JluEw7rwhejtvykZo0ytC
LEB1MS4g0Fqj9h+6dSBMJVSfFsTkKFCd9GMOH13vuNNzeHhw5cewE6OCt3UYamy4oaKp2b2bIelA
40P2Bc4W3PCGVNE5oPSuKnzGqSn+d5GLB+A6DfLVWOb6SAWaGrUvEIJi/vZB7lUgQ6rzOn7hlYCb
dz3KVrcjUpFKPQjpBONDG9CsFdy8Pc4qlsnPXQ9BvQAelBYiAqPFoo38FnAUush+YK1EuBk5iPo1
I5GUSncuoD4tjg2T/kmAinwbnXM89Ui4VVU7uNZeaUvGdW+7oq9Ys9U1Iy6M2kqmBoGQfvZ4eHOH
LStr8IHfvDiOWXDQUvbiyHZzGdaz5c9AiSqkeBGRepOIvQilm2DMztT4lTJG6IVGdw/ohiZ136NP
DS4Td2lW6rSMfBiAMJeN6ZEjzBxOjccgpdLXCmtR1WgO+69PEkC8gHfjZVLippxhWojK+VZRnoO6
HVsd9AjL8lm4xFkXUCM3eQvPOY+o1JnyM3/JuEzHhjhZ8UB2IjT1AtsLEoyHU3Q3n/XjGMWhhU4l
0R7yPm2VorfPZjr/kBM52gGMEdaJexkrZbFLo97kLS/1lx80lkm34YOg4k7qKMxlefxqbkvjTTAK
jjNHtiT8a96NEGFR38YQyEFmXeLgkZZEzxV6gvngmOVlRo+cUby2DNx4vSs3SPN+6P/8fehSwb+D
zTPZSPJ1xEf/EgM68VdXZ20MgNqTjee/3L4xrpFzTZv7gWbKZCuSn/7vQfiGJVjGoOicVjMoUiqM
J8M5EO6HvX2nOCpZPvX7OtAJybNpXrp2ZzUfRzdTMC91tar6t5NW/0UkWLW4eAVVRznqZVT7pm+V
B9spQTYuvRPbJD0AWTVbuCbz2eCf9nk71tyEks0YeN2ePAq9NOTEgwsTO7M+rtwgdM6pFTvtYZUu
cDq2s3lWQ4Hys04WxZYYd8OdhWW+UIrebf3twAQbxFXpfF5nkSpIJG4CKyryqgP5ffHTQDL0frzo
PO50tRYRfGBZV48qv6AZHH07wqxr9Y2675ILtxF9lQs5lrk3mlq2srZTaDUMojhZ77+5rUlJocFo
Gwe74fZJjYNN/5FyTDUjvlfGf60xOwsqO2+hy1H6KxNXaVZ2Kh0XixqoOEDkX0AMtQJqf0nkdg1W
lP1rLmkURf9fqwh2S+iRKRpsfKGBRhCwaFTV4/Ryb79Rdf9JoY5dQhWYEaBdNX705Kt+r9vFwWuq
ZYXZY5JT/+Kvteai6X3giDi7g68f3xL7pHxMawqU+tEpMHLpy4HjYjzd+3OOeEe7qBDyV/m8fGvc
62NJ6ND/yWeWeEqaR4FEO5i4SwSeXk+RQzfxjbq7gmEtEakofTLSvFUccEd43tAooWVBShVFeVV4
V9OmynKKLv8wevyXc+MAR/zmiXtjo2EpIl6fLEyQ7KJgVwS7NdHqdF5EjGQDQ2ILCPch469iTqkg
SHyahYZ4S0JDN7ApBT/wJzOU2M/xKs9bTPDZy+Ti1obahhfcoaTR5GUL0tHrJrgWuibdfOtvkF/Y
/6oOfledft0ZmZ2z4peNeDxpRNb0cjkPvHWoUCfgw6GjKW8jQuocPN/aHRd0341V7YCFLewyuCdq
6qArjYQGwLzukL0+A1a0sBoixazgMHfXs9P7vQ8nEbh7noZi8X4WaoYWrh0XLhzte6WAEFSPAUd8
HodkHS1cPsEUL3+wem1fcXy/kmiAip971XewivBHS223CPfzlu/iBFnj9DaREStKNmCUGTKP9Tny
g3PXnG0haaoLdenq9hB0g7LCqKN9bbd2byFLZ25vx2T4EV4QvMTGZOw6EpzyQ0rOSJNpWAhffiTd
lQ8k/MF8FTtW9JRlNM+zdv00aMfJjlwIh8bGlRVb312y7bdrUDyrf23/RFShqZtwRrg9735AY2mL
gf/VDvItdYLb/xnlSnPaHDeeCBygEVlpYeL5rAlkrsXcTHHdz0vfTByVt8fF+SK1i3tk4m09RRJl
3T+GPUaMQCbfWYczET9fo4fdwbLH+/ZGmgksuVqt5tOicwyQN/mBMxZ6X/67N2hvaOQIrBjaibtq
+gvgWmg6ftVURsPVp84SKgKQBEVxmGdSbVWn/Qin6Gp1bcmOLni081SPs2CsQ2IqFULcLCjJjDac
irq6CNkAl/JNQerCqHelHZWsVii9AFPk5rWAxhVXauPc+9h1hx/gbtLlvtLk5jG29qF+I0y6DNL+
4a3tBPg3+PovMtr/V9wPXDd3Zka7jZ81jdkFz3RKrQZsFPv+I0C0lLjzofBqN9nKzqfVJ7uVe/NX
N6xrCYkAqDtWsRC8SrNM2MpEeWuXrTjfVSoj7BLGd32XcCh5780NOzp/kA106mQF2ReUzQS2M5WK
UZP7hDmg8dU7Bb/6rtOpK29B5Obff5eY0bRguddtzG0HbL/vOBFegBUcv8OLnGfQf3wkgQD1Admo
XOemJD6p+5aFtH6Tx/IH7mYSVf0EGIffefJYcxVtB6jVS3Jpi8bhETXvSYHqAD3nVYAHTVMLPOUg
s1ZFavYgi1m5rFqqcSt0PsnV32Ao56SZ60FxwCxBspJgdxkWnc2Y0iqaGoKMixFWu3nOfdIjeh46
RcKYbz8KColbFpGZGGKYw8ZhKmNM3FDfgbXWjQh2ZI9Kgk8S7bXys9WfopdiMreCJCFpqNEAUdIZ
HZZOk9hVb9q4FCtmfHcZ14KGTC6JJjcI6rq6/N2WffWI+KO/KXTcTM8STb0o6JMoDc2v/lBJ7VHP
kNF09x0DwLtRQvQ+OufgHg0PP52txsYhYci8q0b9Du5cefuv98ekZMcpovOHmEI9LhsikaLw+6FB
GFLsGzXSVLGlHgomtY+29Uq21JynX66Uh40EypbPnOv4jWBcDrE+riJfx9yR1MthwgMSKDBVRq8L
PH16JWGGKaY+lL5cRXyGTxij/ihjulalq1HuGZHeNLM4uU7NQ2mgC3KpWKUoVMYIWCLUBa1iRyxU
R15sh9rr/yNBER94PoChafLE/r89eVMmadeiekBedazLHEzaXv83G9zf+9DAwfljOT7gaPLfM+4U
nsf8TIkTzBhhO7iI0pZvbZ0J1kdop5oelgkKTnMaE3tJz/hCoxHXvQIQ8YqyuYn52Ux6TvYNhTit
HlXtbN6KDBeXMoJT8cNfY2/t63+OEwIJC2KvnYryurQoQ6abJxsPV8VcgM+RxcZq7kaHxXsdM0RE
Pt4q/2gYlUphK7JlQKui4K1a0zzPmw2TNWCS3P0tyD9aUgqq6ASwk4Wz6eo/lIxy4F09X2IOZqri
ZTwhNpLPmlTTjOk+e4jTUOZnnmEGhbfZXSU/+9gK+TTH2kRDb0xJyoZx808WuyiTlK6Nrs3iW6aF
pz7m/ZhJUdpMMg4aSQN+c5Z70baBKgQ0mtj/zE3h5JOwgolczaNdOIRTooTgJF3i3OhLQRSQwCHv
hXClQIhKw/WI5KEDl2CaIdFC71eD2CxXxmdLNdxUH7V7r/f7Odx00BvgJP85mx+eWQsTLvxVc0F7
fx772ahCRem1NpHvKRD/hx49eALnl8Ys1W12aktZAvE0CBUdH776c7MCqPN1Uc3Z9ewV2c3WKokH
4X97yBR05e0jfeA84eb9eeQu4Ij2wWPj6+QO6YpJF4Mi7n6ATCaOf9My29fOPLCiWsWDB3s5F0uU
VMhQ9JAAsQy8ONIofJGORvu6ck7K7pffUOGTeiiWnfAdghAArKFBL7SMC+y4qwlnqMLU9iW3ySah
wY2qX2LFcRSt56PHOW9BtMxQGn/IYKlHnHRmm9ray0jk2/c3ggSkKrZ15ABxOts/LSeBHdZbNSG1
Y6dw1vOvjo59ksOq3qKG9AdUVsKALIxEMGi7S+e7xwW4VGl1ANTrW5UYrqIhgJ1QBFjITj/2z++W
rM4c5v9L43Izn7gHm76/NxTd6BQuJaR6+qnesQ1ABbwGX36ugnrV0vjM3/bb7uFBqLheoP3yi3OW
7DyBY/uCi4cNvMNXnXaggITgqG+mcLT3B7uvQIeB1L/wPkpA+STXIBrIAQoCP3UgAxhf5+MAJWVs
g4gdUw68J1w7gHFKm2IVdhBbZkHyY7jlKQ/XRBysmblZz2dorKjRPmEQaa3MLK9N/CaKEOaJdUGx
nPAr8e0bj9gi348sWhCTv+d27es4lUT9C7WwhE/fG77tx3KcDvbbR8eB7AezFc50dFtK96Vr2Bq9
uEaoXxA9QmrfAE92yuPljmh++dtPLiXeOAcqYKcvcZcZhgTlDQ9e/8/S0i6nGSix1ghNQly/BTup
MoKRL8eDv2e79oJpYklLKogZ3x722NI2uz18eeXkAm/TfDWF4oAMuoGcbMjKdxFyWHTumT+bTwdi
9tegNBI8Mulgr67yAja7ECumyqOi9TYUdLlYRUbTtERkBY4Z6WMGYkCvU0C0TVkU+7jx3b3m/h+w
noqAyojjpI+VHoOAOo3FRuKZwG7TDrxAB8Sn5HNHY60bbIUlPuU7VAv307qf5+Y1yt8AWB7zDh1R
zKCP+DZNBxBFkjo1P8xJ9GbYk/T1gaRIG16W9ht1YgV2v5cC2cfFkaTSk+IA0riCviurajcDHUPC
sDWwjdq/NhqnlxZej643DbuYhrMiFm5xZ92cpog+ld+82QHmmzLg5PP6LLKqqNoYHN9AOCTEaKm3
i1kexgEq6kUg0r790V8moLv525+CTJ1ukTVr+iMoe0YDxGbE1m1jUcwDoFfv8hY+t0av+r7HvTEK
FZNaLVMoostYPO/Hhpxynk50zhWFTMa7ck88WTFiStMMsCUGe7NmXgOSu7PvZrKISfUU+f+siMIh
oEinX/TPUI169++i8bSZsTYdvW9fSWnAx/dHsGX7Iq3TGU4dBshC/faL2CQUzqnt55rNKbUuGHS9
I70kGbk0UY6F074F0tu3hJZMW+a8nmhjaoX03zoDd/GU8h3NFI5EqxNePTkDJnmI4tQ+4F3I21mX
ue5NEM1yKELvOKxoDjr8WaX5bLjyZ5sH9UcuWBwuZt7AtEKVxwA+AxaU/nAtkiOl+W5i2IDkVuDr
sybZAHFUyRhzkNKx/g9qv4jCPvGSpOEMlhB6YBDVaSKZC1Cev3H4/eWOkqdmtZlqjlOjuH9H/hfL
0m4uumn+lPeaeExGSlfxfOXVKHgnI2Q74gZK6YiNlrVvnnzVlKWqY3C+T3NIqOlpzfZnLJeUulV7
rAc/Qrq0X7ktFIOlXX+1bwHeCsrrANPs/0T/W2yTs1tMdUkSOUilXkHGZs8FtAapNIBV6GqUtKdX
KoRMRu0SiGqMMrjTr2jSaMRuruBx7KERPjggRp2HZANEHekh2wLMpJWyN+gdSElITVoleHCT6LWG
8suD2DJGRKlUS8c3A6zPhMN8JVFAklU4iDWunWgGdBhxwTyhnGMTnytd4YtrJmJ6XaaSsxVq74OU
IwjyMG/XIgjusnztJ6RTUqyDl9vmOQxyE1tXpElvUMKAIXC3cipWEUbUAu4Tnx0w0hYTkNKtW49Y
2x86rwAkgxhxUABTk7x/WNaqtFytZJAP34/HeidU2wM03N2whR5KVxuzgJSp0a0gqQAOIbGQWxcH
X8JNUZ2WPQqXZQAa2DBAdw5Um7k48TWOg+b4Zow5wk7w64i0GZhtyRbnLnLggMx9sxrOyCzm6FL5
FGg1YSzcdK89gTbbNdF7e94Avmp6OatdRIb6JhsswwQuf0yB2wOWjsuJqGzvaFUl4uQyfhb2fdRb
U+za2s/IVpvVZH4PN6BNiMRdaauIb6i+vQHfy9SF/aJvaF3sm2XqNcZmuneaUEkypa1FZDxgAFEh
PRfI0YP5ffAcUMp2cLNXIAWjm3Jdr0SJznLCbTO/yNWx3WGb5hLB60IjnIZDensnv/PPbCIxwMnB
A0DtOj4cSD7a8dkbZ8rdIbjfkNSpf6Vd2mHkTV073NnOIqEB1M5TV25MpuZ3+55XF1GyXxNrO7wY
ZmRwWe1WK7K0NJSlzPCGg/fqm1bF5f0/lHqET/NV+0Hv0Spitbtorf7J0SOCz9oYuNU93upNqNPa
+zeBlZXN8VuSrPENa1iCgQJPNr59IdSD0WfQry9Ywjt0BFKMBscwZZPJb+gIkfwaLiyX4oHidYZl
vGZhA4cOpkyGuzA7kxkWKUxxUKemVbPGPRPZjB+UIBx/SrS5OOlTiZD1Hni4r1Z9owiDYSUMz1Ts
OteaZybdb7KW7yXYToFsUo8ThVuCPnlMIIZbsyNTOfy2UuLcWDHedvURiIC9KsxPQ1wW05UEVrPw
2dkWI1lpt1d6pj9iKHDBB3CwlLrIXM4NO2IZi2M0fvMzsxL7/e8GPmui8lse/trb1qGM794ZkEyE
0gm70+ihYiZPTSpm7m+QnLQzDSXN7hg7YW91vg+SVLjm48mgMVuRZBJvatyO7NTfqrTC0RiWrneC
vG1t7Lpz24hFj+V/VUELys6JLyoRgOf4ysm6eWPONRhJ9XQTuK10Bh+hKfP7OBLtFTtDRkQ2/6v3
jaLq7T6zUcWXwzZe1NXne6PzkVFNf/xpqnUZB4e4q2646al78TK+P0QXerzn7FcBfS+VQoNfxTpn
rMK9S+VaajNgTcZzSE3/3tGRmRT7b3qs4cdZcKC4yT48O/ynirWstIt+K6n+ICLUnXXfCzVjlt9E
9bSsU8pGEi44MdKtdDjATP/0EDZDR0E+RsMjUIfr9jLaKoqtj6qhxcUKNEYnE1TAcYFkK0ZZe5Gc
7HJ/GB/vs9N4HNZA6y51BSKUj3glYa2swqDRfp2D9JA0hQx7bxEVjOO/1TNnM1DoZyKcO8HCgMmx
AV8hoC+PEKCIo4lSS41cU6/Cr/44pzCMzuH+wkTAzM5fm1Zn/1qT1eQh01sK+NkyZ35VyXMXZ5ns
bPwV3WLGgR/wTbYh3OYVqccMm/9NAHo8hC5j2TlrEw3Qdg6ZfkBY7r4Em/1Qimsh4aRVebd6Xt7w
+Yee04LicIqvCjmUJwI0zdpCEyn2I9UjuvSCx+wWQ0tUs58UvhdLwmwR09uzRfM9RQo11t8BhDMD
6RRgaPqmg432XKpF/teQWd1lvi2zTasRDIpsvFQxJeO4I/q45dbCa6tbvFEvZKj4gaZIKgn8uYRk
0cEO4BSvFHDlNsoesJruA29HS1HCiqGXokivgMBJQ5VxBElsEb3Pw662hYYIrpiSwU6jenrSiLW4
HfmViDL09Y6UJq7F9phWoTfWML/MyC59fyTqEf88Dn18WpSfwpMbQLCab+vh4qMjjTePB6eAIfpp
GMHsp2hCMCAMtEvTpOJ1i7wOuMd/TsoRs7DNFCQFChGgFtmh+jTF8nTGT9jJG+Sry5DZ3UiOcXEc
i+dA8XSWMLnHeIKeCPiDusPWizAKrxGpjbhfUI/B9lvGG72cY7iuII0yYkmxLNQJRqY82V0tuy0y
pZdGBOzg6O3XgohXT5IZ0bN5EHQhkZQMC92RARy3fFHKEAc0vBNvfjDp2Agj+FhMefRswq3VlzaG
lTkiX0ELYrsv0Vt9GYFfDMWDiLZ1TzEl5qopZbI1yDBF2R7q79CRxifRoIM5J2SLzl8DRvIK4x/q
a+gFRBYyLfNjsQ6wFFTLnLkBJu4M9/rQxyIAiT9NRBnO/gHPEEjHjDElzxTPoQX8BnG9nB25sez7
RwNsDyiWjeHxxMh2vZbfIdpuNPwLXyhJYYQJA/c1pGB3oVS5Eqx7TqRK52S29D9fRcqs9cftiUHD
GIRn/qmsZi8xEP0FBJSY6iNDmsYVGiEUX2A9u9u3Ci5UtzFcXbspfMTQRc9XfKQ2wFKv7jAaKd5U
41vzQYPmiZcvdgPueRcn5P0BQ+ljwp9ypnTYz2XhVpOQ2vAHBJirTdLhbb6nZGxUrX7TZCi4VuMt
XknYdUuSkA+a6nLCNdVjo9ad/2GP2nSpPUIpynQ06sEEwWb2L0umiWeIcZcDeJGOv7PEZB4r39QL
2GHWJAjIGG/IIX7LUF8y+HoIfnMJ0KenbvHWmoqZ2Vg7+tKerzUkV1PIRSjhKSilrCDOq+jycWMx
ZhSJ3E8hhRhEV8Q8+J1k6uex41t/4mRGlH38vYsE694rLSTJd12In+2JL7odN1jr+VKBTwYmrt8F
/kcBX9tpWKpiImnJM1T1wftvZF95kobonKJS02W5rWlRMwJ6f6IhUTeqaPu/CGg0ZKtuKav1ulOC
m2bmCS1J7NmNiqyL87zMZ/ksqPMfEF+z/kTMJxpRxfd4CpR1bGr52Wp8339ITPyzyA6l0LWyT8NA
DJ8WatBLbCP8VW46u1WKUhA7ZHWaR+NAUgm4a9/Tw2Ex4IwOy2w6SR5qw3tW82x4yWpDr//UwQ8y
2S6Q5WV69wF/jjVLMHWyIHP9x51OMQgP8ioQ55qWR1CLYVdhAPzwZ1Z8z5sjxii4TYZp3/ibtyON
IQpZ1J6BtIvQrSY2wySLz7RHYM+pNqW7vGsQlMczQ8ZgL4xIL0RFiYFr+ccl6HJJvHIoswNeNSng
BNvlvogamExIYsh/OV9kD/YysC5jyl9QIwcuEtHSiV56sDtiOOJxriIPUBK+YSPaiiOEPV59QLeG
x8yD9XtEV5OcK4rIq2iceq9OtxCYCQ8XiBBAnviZD+P10ooAjCshuDqJzFdlIJSbgUq7stAUUYYv
1ZBVUNKulLCk2LtQzXFVaQbHVO3cKLG+UdG50xODHNrRj2t6pPHQBA1DDhy443p/AuD8/T0pay4W
vUV0iLvnO1HftZ6Stzw5IrDVfUYXfycqbOgpxqySbTjLOOuCmo/4VTIpuqQTnwK1uh0aPE5rka4Q
ZYG2hSCk4BeAlVpnabT8gWzVKwSg14nKJtk994nbLISj9yIzA+eXO/NK8dCEz7MjJWfhfTyVUNhl
2Rxa9yWq9VnXvu/t6NSQ8awy06Kx2ehOvH6Rfpd8kxNhD2bJZYKKo9z8+de16eJ5jFYKVM4A9tmw
zg/BAEoUWNBb+Y2KNXoxRZECk5nRqG5hYLocMLv7Iz9PL5Nss+Y1BK+FaPFPSM4GcVCcjnhV+g1f
RwumUBwrD4FxFy9t6uDXHLSqJytNbYmCFEbllaWX4aQzbQeTA2xdxO0TqI8HO3NGrlQMTXHD7LML
35WLtab38C73sOEbNlVAc5CIzozbjuocNgI5EChqu7YiD219v5kXacCGPoXVUomTwanq/vP+QKUg
QeQEKBTg0w7WeR0pVPfyCq4iqbOAOVA+gpNM7v19PlwQeX86K7yOtfxWlC2mBwN/7Uf7XNqx788Y
eHPBt/5/Nr+d4fez8jmuewffizzQ2arcjxInX+3e0uaagOGmiaTO4l/F53YvqTttxiOegy1h6h6/
S+yvLUu9uEF8/3qMvjmA5XGr5rEj2Z4VdC8zrnu7BkbkXGniuIsu2iJHiid1zMNlQxxoXa5MKLln
ZJEOl8VMNedpVflb1yEahAb3a7TFCTbtsgQNaKbZB6CRiK/lU83Eb9YJ9YHDZz4r6PkfqiWDRNlZ
iEI2eht4clniJ4ygM+ijHZQ5mBWpGIZZzzb2vBdjPhCzyXUyFlbCuHGkt6OHU9R2o/dCM3LW6ux+
EatWNDGt5tARqWMwG+N3cKXLjXUAB3SNJa9KkdWU2Tz2QMIYGrmNcrHpdabWVnQU/6+K+KfttBAM
GIZsRJuzMF9XmuGc+icB5kAWoE301xnXF2C8Fob57WOkUyoQp0txugPv64UVve8FyQ2sl3pUTwdA
Ox8cgYz6ro6WSxRmnP1sj8bdY6WgwILcHZ5jTz/wU93Wh1a9dGsBFfWX8NDWKZQaTMJKEay6B5y4
gXSEFKMxV1/w3ZmZpyVndN0QMmxjoq10QndMYyOvE8X57a2P3w7BKWBPtU35EFsqrUheXVy0xE2v
nOCu8rrU5vbqrfE//zHDNA0+40kxD48uQD8zk+PlkobR706w1m1A+ZBns/mPpbAR2M9HjDuQmVgZ
u3KmYtt8OFkG7TlhWgkqnOzy9lzCpslP8njAbXU0rnkIGUuWxgyO1+W7tvZZ9ttxS2xNzutgKSXQ
YFEdEz25GoYt3MImGfjzMhb7vob6bt6RljGgOkTaZamPA7lDJiw6VF6M7m41nl+ZEEe8bHGbjR4b
Qe+ZC0mv/PqaiVYlWDEOfJW4rWeVZII1937Evm1lti2jJ3z7M8IFP8On6KwDcDiTjroaxu29tXTg
tClMGT/7F+uV5OsGwtUKGjaCkdsV0lscPqss4bS3qtA/8jLv7rduSMECkowVbV+1vHBO6rrz14WJ
mE1XqsEaPcZERRTVa8LOLJFoWVTI3UFm0o7UGz4x0YXlTNryUweKKFWLjYAtizzMYmpZ8F6h4qMJ
SBEuU/1EYrpVW9LazijhPoAp52wTyJy0WWT7r4UQCrt0imVhXxDe6p+sKUZQAZQ4t4Pr38AeOBlZ
YkKhrO4Gbntq9BOkCv9LLROaUPwkEgfgMgPKcZdzm5ykTl0iO/xzC4HusMQdKHCdX1C3ERm1wyfz
6hWapFOwklUmwhhquBiqBAOEvz6L2MCIjmFtnLIyj9uVATRDJXsvUeDR3IaZF3rS6FReGCh5elTn
dL9o2gIoBAkCTmyxlPmOR7YN0IdE5KGUCygIEdwm4asB0cO8Af+RV1Jg+mMYeU+ihwYUknOH9WOm
WWjSlwBcqp8Qkz0mKdLghoY0y9PnwrRf82ntR93pebnZmib4XjmzLaF0dZuUNh71/R5O6FAggS9n
Rd5VIGNp+4Z9Tezh02ocAurTjgsEriRBxf1hBIty2SX06t58nbROC5tWhHQPWVe47C0sQiNS/sIC
dvRkLIBlVEAhn+IQLtYyr/UBYTa1m+Qf6G0htYuv/JYZgjQ+gaTT5gl0/a6EKQmusOGd++358k6Y
x/orrWi+A1r+2KIpFVs+0eCTDor5QBY9R1NUbYO22ipjhOCtzXOHxIVIhkKD5OTXg4Zicg2jbCf3
+t1yCzNmMvqrZx4C2QWymhJVjw+NxjsuAFGXld/natlqS/eFF629zSZa8n7bzRlX2/GCow2x9MSG
XVJN/ogwFOlR4TTeDZ2y9q7eEMjB0e/KdBWxLfd1ixn5qIRloM6CGsabXnychT6ry3O/t960gjI8
OWT9vvc3bRfbzJzVJxvD0IH5Gk3sm2Yd7LFJfyF32huqURifb2q55v62mXtvIgg48VGaD9hfuf3+
3jVSvRA90HX8QH5JNBz+ijbX1ap8R6O7B+IzRp7oqU4KVNNO3B8pdx5zEc5WASeqxUwOpqAtjqxn
ZCEyQ+Vox88n2tV4qJP5bv5EHCYCQ3wogeOF6dwTd3zH0f0qK3Ls+GwKRpfLQpBFjK4F36Rp4oN4
/zypRk8OkGGTa5F17YzsRFjwZLUQc3IYoovHmWlcKiuDOCJbCuaE3Rox//cUKxn6rYwbCra0Pcer
9r9I4fj8MJj8TaMHxF4kVyHGpxO4aEILNDRtNNfcqx0f34fyGBkugNfHiC8Em1gtmMhVatSro5Vx
pLmHdGGAN82tQtjRYq9Amyg0lIqiHgyTUgIBKyxWHBUuyp1EGt9lp/DU8fzMeZJ959toVMBr0kss
Xwz4KCF6UZxQidCK0Cb31TLcWfhtHcTRV5/tE3Byk2zTGCDQETN0ZEmoP+jiHVVW97WqyjAG8ctg
OLosv9YcXlgEGyTHTZ6IiBQgl7iyVvLcJlyDpdVJmMetSIUK38C8JQYzzH8I1vOHgHpEU56V6D5N
PPWvz1O51QzkGqHgMRqkpfVUShgpusJCDrSjxCZiKsLEQCmUgII1lnkU3UnhHsr0FRDzJh3NRWtF
tdFKTRsHQnus/FgpPZ4gtCLGVt4vif+40rErns+qlJT6v1A9V4vK+R2grPjuOtMY3tH6Ee7BHgWp
9At+BfI2QRCBv34atm4hQOxrMLo2kFYJHyJOALhkNc8sD4uWaHOUzqlCKhSuFL9kSziCruJpPNQf
jMn6bXm6ptQe9anvrwBpioDbD4txC/G6RazRnRwbH8tVSQlCd4Bnsy4ZRcEWb8n2FdtHKRV4XNUe
t0qzOlKRyWBEYkKG3oDQmMTpU+kUtNVddsN4YBRsBdxwSZELDBaDGuHZFcC2om4LAl/4284LeTZg
MAk1v5Ad4X7PBdvXOMruqrjJeX1VcWQ8tLnkzJlKr5Me28FLHxXDWSbRcb7rZ5E/bzojvhQc/2rg
M2/jPfjfIqYFliJWW95gVc4vXYagBdmHobxDJ++06qGUQtwmmMaAkL0xxWJ/nam6bL1NBOAc/XAq
97rw1u1sz60hBtqx2Hs9d4w39Xltm0aRT1QiP/sC0tyho8bHRYQTMAwwNly0clS+LKExDy7CoiV1
D49UCoOEYFKLTXrbj9bqem0BjSE/eZ8zBi3JEatIVfPwgs//fDPMLvWHjysTRZ6uZ9Mm/GT0Oy7O
Gr3fDQVB5KWkOmEyQSQK9iwZHcE2gHnD9oBCgaG1BXmJXF9vBSuyFxg6dcYxs9ijksG/uqH5W+x5
5yl3O7xiD5CrIEFKNGY75HO3wIt+SLr8VuyVFwaKz17IuvIp/6yNtREaiv1CHD1Psh1wG504gGfo
gHHPsIovihSmnddpsTHVIhLzl0G4ZNDci57WNzIpMocxXOvawIAtc4zNtbZhpc2h9c9sqnROtlHe
TR9fJRSJR30i1LZqDBXPbrFFPBZWutiHNSdQhagCSTTR8tWtI1f7elH7Fg12IM0YeH0en+Nrjhlw
yCYZn7Ab4JVgOL9wjo0Qb4zaaqB9QL4DFTkpSMx/kjylmN368JCi+bKyCU4H8ZMfLZe9C3oIPW4p
WJ7ik+09pxy2W9WEPjmiUx44OLXEb10NvonzpWIAbdwXX/ehB1r+g5dgiyq9QqhNxEuHNKZ5ZcKe
0khv0CrPGGcVI/fUBHZaTXLzqXuFZhN+Zajm8vb3tk4kl8ayY3z/d1XQWMNB5xPFp/eDUB90NwV5
sOExuNszZcjGyEylnylRvurrfQMIOfT55JmVn6T9IQU4InQyRIDE5ch4dKvxMzkw3tGqH/qkZNat
dFDwYMRrONmFKwLGE8txKTSoWnOyNek8SEWCiywMrV//uyDlXpuyC/RpVrPLDHfjL9xc2nEXTXX9
c+Vr2Wj7HFEsNuH0uLKkcJzxdkMIPOFQN2+BpmZuNLVfTyhJvbzhBRsVPE9drsQAozigAohZuPMo
7ZiFZ0Wrphy9FpGUgEaxLgRMEiAsTzSAjgWczsfsjTi2JLjS3lfZ5dKurfhN2VvMNTqlNy0BaXmf
zCQcOMSu65yBKktrIazYTsEWjKT2nq8gNVNptnHcPqGynspqQslGwqVEww5OohwhwfztpzflZhaY
7blGFq4wZA+xXjV63qYgsqxDexfI+i4h0IrklacmAAaMjLR7BGOEOSNJ+J6dX7MxfCmBHgrcLm4A
A7B6dutTHB+KFq/p26yxRHV9qcZ1jkd1SY8jxp8TjFhAO39VDgBZEkzauBnnmeGCPRkt4XhZ3nVo
8RiiexdeMRyXT/dpVoge7/7XRNFvjbh3O+LtIMANLckrH0dRdmaHBK8OHvFg2U1aXTSN3Ms6+rBA
YDqk9Lgj+dHFGXczptmj1FkZlY915C6pFAS8cu+dkL4yA8dPzBorEHbKeJMgi6WPbdeuwE4Je5mK
Mv84jtQ6EGY+q05lXGsCLFKStbgdnUj6RBmBj7YBAHVAKSfICDqS4aKjddyYWLWpQw7vFX4EPXsV
3ghiMdC73aRifMlkyZ4l54WyczrzVWPOftrHTd1xonm+rIfN5wMo+JSiCo3tSh4HLcjpStTvSc+i
t20b1BzCLOkLarUoI077uPK6ZwhiFbOwSjWkL5qn+9YGcThOsjUnUneqHN92125pCcMpl1QgThUS
nZYAIry/IDg3nfH11zqbYIBK3bZkMnT+ENO2RfgzE8/meYrFs1+9uPGTG5RsJsTaLWQkNlz+BvMT
IrC7qoUVCUjAR5ttFppUP5sJscpip7kMY5L4M6mEoGSiDp7Ih+Na640HafCXvKyhfmjHNT5ikHUg
mhHe7172b+6buE/msJH1rcMhPQiqOOpr2PHz0ba1ri4z0mjpGI1a/n92/TP2FaoC96Vmcs2XvfoL
PrucXwWSJY53UJ/rTh2DXmq46D+sZFzlsV9IiTQeBP/5OLp7P3JU1ZIlC1rXq8ZHeLHWexTFZIoM
6NcBCuuEC+jl1+8SqFQYaZle4XI5sK8xhLlKW802m/bvPE6ehb93/cffe3q5Ssq1qTiO1qTeN4jj
q8W5gEBHbOQ6TS9xzHDgsJ+1bNjocdMzCW5BkfPW2Qr8erSNlaaOGfNQ3AORpiQxQpEvPIPi84XA
I4fDnO4MMfzF697cqw/PxD0aqGpMsMAcQW6riH3oqugfmQN/64tQtHG5B+zmKipRDLe7v5BrGk4y
wWYXVdeOsN5KdzAtx12wAlAXaxFxyM5Z1H6h9LVqoPQuULsVFfgAb0ql5NANY2BiUg6VdD3ydUkd
ozmpvt2R5nzggXgIPRNcieRvbYR0/7c1M2pd9ZgwO9D11QPzFk+LNKJYalKcS9HR3S0gpfn4DQAj
JY9fCeJjYpMARbDUABK00NOPOpK9ELLSMtuU/cI7FVAS+uoH7Y8kfQcQ/Q6k0G/oAmT5u+Mamt/k
ebsXXWmcE9B6vhoBS8/1IDjFqETJ/MOIiELWBbGfCg4cPy1iQRSHJOCpBi19jMspycuuRdi857Fm
c9H6N/o6IXEB84FgTtwDEjQLC7mK74DK9QUTnuhmtcO+/MQg4v3r3NCnnEPBDvQQIKEZqf/49bd2
0JHuqO2ls7KB1zt99Nt+o0W6GRAnpreU2q6UHYWEzsUM7FTGKGGvBsq2lBgip0qzZKUgtnB0uiLn
rDt1LX5UcvdHoj5NOAGMHlCVzv9SG4tsJvNslnHdXJMdVoHUnUkkFQ24LSUaRbZKvrH2ZD4eRRaI
6Ax+Vf/m2eV3cUe8jag1fNPkvo1HiKaMbkj3MDEXKfej4p5hpnhUqyFpx27H1p9dHNRXAvemjklc
B5zgeNRJjSL6Mu5gTwnltQ/QEmuUonYYe8r0Tf5ZpJ7GkFl6m93DP0UEWpQNLjQjBa35NVPcQWDn
wPF6TaEsZaYOgUm0gqCWzmdZmw6CoguIX1xb4exctg6Md3gSez8m9mHBjnAFCuFDTJZoDLqvIA1b
+sf2Pg1wifx4hooC7Eii49GkJP/tTykycwSp+yS2+Fd1iyjDGGbpKyjpsJX0JIMRX8ZoYj3y17kZ
CDvq/LMKd4g+KaL6zKw4lihwvSi6fKOGqSksQY2R49JzNA4C9juiHqDai1wIa4KLguR2sJBrRfOl
x+ZNbPFr8TJtfjXqn35JV/W/rFO43UQyVkhiatcXhjo6TobmLKds+zJ2ZWDuYMIrK0NjP2FaBZs3
AEaI/uOOMjvK9cu7D+hEnEGdfWPPyKdpUuK8Vk85iVhZH29ujphmu7mtFQr/+L5rNH0Cg7+cQBIB
JjRsZpFd6s96HV/Ysvt8pXFwV5TgkjGz1zMifmUej1PJDoMd3ihPoPvKfLrUFHpDmrPOOK5RYMzY
EN8X62UU7we8KIill0/EawNDp4DEWsmHgWL7eDFybjUeFvgX35N25ZKbEfQLyeRzkjmn4+xuq9bX
h72/7XrXCAQl1l1O4VbDcEnw+ZACn6K5rmESijqtxRifL7r3P51iqHXzSnFQx03CBJvFM1f7q2JR
pCxvxtQlgGkm5p5CuaHUIeu6crEA/FpMRQGrPznQzhe9OQpySIP6rjw23napLwvQwI/qtEbeowUX
9Ngvo3V4P9Z/OfmHgCne5bbbpJaEJYzrjH8ROETedUJ3KENEwwsu9Q+hfWEZoRwU50enEhaU9ptJ
qjT1X5nCcmhRDkmlD3A3gskS7aUgChfYLRrXx/HvCPpA7RtI0aQjyNWS/I2WYE1GWHfIAowf1cQr
yKNH1pBdNPn6/Pph1N6RSiMouZPTco+6tf5WC2/jM5Jm0eREjXgcErzo48i2rS2QTlGZ1XPEr7vX
q+TmQ3MNXQqeFs6zB6Wv4uAdCODMeU/ssYwTayIitfAB3U+F6KWKLHPvF6Pz3i5fIaLuUMwP/rZV
2PcHCL8Q8kPYUKLIm89Ad+6SLkcwUMj7Fi3mZ72Koc6Ddv0eDN9bvbDYXB1TD6W5DfWcCqVymWm0
JGxOEcHOKGwrbo0UjKS99KPEuXhdzbvHSjnb6vDUEdTxbZCWhUjPfwebEAacV7w5ZczJQ4iX1XeU
ahJCOmvuY2d+ksIzW/Y4Gw2BlCNJ0hkBdDivh89AKjkNlDTcmwu9OeV8VsFAxf7vJnFGte7vMWOI
cfZB67dhjtEwRRtv9QJMrjq0r3g6rEwwtSFiqOwy5qR9M7rl5OggzBOExAD2tLGg+8+9HelotYYF
kVTPLOlXqiO4BajLtOxETdjALPi0iF3lhXgGNUB5HwH+4Ics5DvV3Nywct2OfRGChzBhJI7lPxDS
MdQoHR06ZHWYbDsJbIcDAT2db5W5kVJiGGX5z82VZXiCZIQyZlj69eVkisM4EtCgIUnk/gNn+wXZ
83YnJ4BDMm3vudFV9UKwwEFH4zC93RJegBq3j4d1JEnSIzIdvjl4YEJ7g7/1KkcRNnAaqy7K6G8e
OHRSFTiRZOxbac88GdH70vSxISVA7Wm4X4wm7tTr22bQUt1zMHE0dM93WK3jDWsgpKb9s85yaaZW
F3O8qw0iCL99aSG4MYVooUkTk+rAVm8YyB5QczSSnHbL82lq4y8DOIh/+UXawBoBZGMFs3S9xJXd
P2N7r5uVjUDp0zkTSt88ZI6X+QYNYDtd+8ZKbT+sxovrvb+cLxNAQf+b/KpMjR6waNrou7RnnJf1
1hdjAahiVIHQT93+DOmI95ixAaGjZCu4txh9gELT9/1nTdbqoBl+4S5M2dfCC/7R7y71xygt4OvO
+KQSa9co553hsx5nsSBLmTeDz4s5pdEQNEEEJPZcQMejlviPGsmENvxQpP6uEl7O500QXxPBIhAj
N2PGbifZTKwIcXEQbl4REL6y2OKFuObSKtWl1Wn4in0Jl4gc2QKEn0GGvtPCGM2Xfmviokb/O1zE
EZ0BBpT6cXwy2nff4poXSxVLIQUHTzqD4A/mJgggZ+izjzCzK9Xxo2DW3Lm0o1n4/q7qWnk4CQtF
KuJ1bGcBFDU7vnvMp8Cmu56EcV+m/5bybKd93t3I/f8xa/vyhR9IPTGe4w0jp/y5faQ5dwoM+ByF
dXL4FutoMgtngAGe7BkWKF3ABshGJ+Vhy2jz+VU4VopvJxmkOG+gYc7wLjSvWWNUwzmsV/WXrpvg
vRrNPu1d2ojFTmaJ3Jqje3Gc5fk8suP+pq1tKM2PvEmYjVBbWgokV+5UWQC7uHerOrB3GblW7etT
KdlcBPAKw4BOH069ptmi+V1sbQBYc//4eYBUpSyRskCbO2pbanrJt9g0xMkn+lQm59AKm/oN/V0c
0udUbvzrwB9XEKdOfN7rmLF5IirW8kkHR0f3+WY1EUJwge6hXXabMWUa5GiNNoXWx+DjVjYsJjXS
EW4Pf6imAtEawYS9mH7GJef8nv54UjDgekAxggVqorab+amcuB/abx8AdLJxOTd1aasXZeDpS/P7
7GGzf7mpu9tdGmCMcu28jyH6HzL6lZNvu1CmEt17JYWiVouIAzHt+vpOXkOY6X1AwSWY1DusRDKR
0oS5Fm4TnJXEszults5+gSZyyEaAhYqzXXsFuQHO+UuuC480Tio9BUSBnvFomM6WqwXKSIa0CEea
rxAuHVOg8ZuRLDe5+Z0mh9QG8HEqllsLDlrWAJ1IlnKNkdgKYKqUUcrseLKSnhHp00tu6MWTEs34
gAVlBHkiJ5oF05wflhujwVB3RPODmCNF73roTJ2eP8J0hWySm6QN0qhmsd7E0lOg65Tt/D12I5+N
dr7CORFMJ/7kZ1pTqJj3tPUOSCowNRIN0heuw+HSzJRegKVuSO8TiHiV103fMonqNquEY0G0UXVT
c00gaWY2IaVKBkyly90M3CaCcNbhjJc4N+dDhiwG4SDvpSleNhrVXfLvjCjfi1vItiB08mht2wQI
cDjwDkj/Cu2EwPOWDfXUhwNoQoTgOz8ium1A2xBBKB2QasmSfTeLhFGBagq3jGyNITMWpd/GC6nk
iAfoEI01ZKJTYRk7u3B+x6spsltxvXytaA7A47cVDHe8G2dgnK5wL0FEQRLZE0X6iVt/kEKDBwry
063oDWlVHepAudJEI7ERiYHDfXrdmRPwihIG8AWU8X1FntJOIYSSAC6EBjhwn7hPL50ANe9TTSIQ
75zmOCfmKyp6ZntmTXw9kXQuKDsFthGinooLhzxrMds15xhR4Zu5YLrJjDWrKxeNsYYNVRb08+Q2
z0WZM9rmrIgw/mMWb6pk2BOzwyvflI6Y0zRMZdpH7xTGLzS58yQgaZn2cmCm/Ctj33icsrTZIqEK
bJ3PFMUweHVY4x+xGClfNDEvpYQnSlos3fjSanZiFYR5Myy7AS8cUj84Bg0SgVC0u9ahXzE+JAG1
K2GH7c3ETdZ37P5UGG1rl6vhvG+dkabJgrQ+sVD/JUrHHWcndZEVCatfnsmHTAIfDUNQJdlApU+C
/slvG26mcsPThClO5+BCRFAN3AV0M+WBBUbrxQCWS3kX3XPgiv0QqstqA/Mp8oG1hgjmt/IiFcRH
09W+V+HuC+3ltUcEhIKNlJRMbxdlQnaXrq3SKP1U3eS92DJX7W/GAf9mW8thSQHMCXkuR+oWHVYI
Ue4GKdXHK9SAoSdJg/AkDKCuJAKiw7ezL7QFWf+5O4Vgw+sdaHhq2GGfVzH0NFoXZ7PMNBF+0iip
SFoVzaRZm0OvrlSEOmiJqvQHD7n8TlP/sbgDyL6AgI9/3yrloinqb3BsopUz1LSm1Sem+xMMICK/
3/SN1yQ0g6PN10K5tHYwsC3kwvWHIXgCd8Ck3mdzxiJ8MOUoiPzhg/hDBWimE+WuVG31u5L2OCY9
x2hWEikm7Em0haDMcfj/bnGMQwaEPDsW7p3oCvTi5Bb3PF/iQ7XaylUXoC8CcrFjBqvNAJZPmGNQ
8NJiXy7X8aSndaZZ7hDughQ9kZ2qZts/8Y6/6fNaDgKq3aNLx8m4W0KXT0gRu7K8cTAtPJ/GfUtA
16ReaTFC5hgowCm+oPk3D+VEkdH3+JpKFv10pZImA+8xeISb7d31RuYoxE2OdOfBkDx/dHRVhgdB
UWix2mFJ2Bxh2/trT69p65mWhoQcxrKlvhy8DJUG69SsmMcU429u7fxalf77mk2EM1YevPKalbH5
6yzDU2fyBOG6zj0TlpbNIZmW961XaHN6t666nJfkqz+RAvwxW49BHsC2cvBGRPEgJHVFaPxJd53y
yD0sXL7iPoNALUnYWLLIqijEPpKVvsfuQZiUIjXJdwXLfAMjA3bBE+P8zcl7FOjlCt6Andkswpvv
7CIAq9tct0NDcEn2ngWuCFq2KUCsOwQhAZi9/8bT1xzBJ1TOlkfyMxcqeVm1HLnBWNWIVgJU7Za5
hG0sMhQkpzKcfORuQSibu2fkL+vJzamwkcTy59AMWl3ARhsPe4SGU4GI4Tkv82v+iN0HgSoVdVr/
e/0miOIeFgPlqtKzft97/Bq7IfMZWRSpW0G9m2KEpn8WMqGkuJ3Xf5SIQEsLG0fNuuAn2IXor+3E
X4Jnsu53E/TmM5hlCXZP4336bjnyYtDk3gzj3c1ceibiSn46h3USSsiyeWIlZawRniK1XPyZ9Yme
8hYyswKbHh9Rk3cpZ1wmsQvlJKQe/oWBm+ECtHO9hqyseHqXxMwApHzkDY4AkPqD7o2sl+NiGbLA
17fcvA72dSbQuHVSmL3IgTq1FhwZQzTYCSHOgMxFNJ9MzNYDwf/W7vSrpFLBfR1EyqN5IXx9akBr
ZpUATkly3m0qPzR9OENKKKoZy4v5hVk+RdGnNgHwpeO5qX3YBuvhvcM27HoB8b35uFpXmoou+tJH
Q3Q/IXqP23A6KT8knQT5JEfy6WenQ7u/78x5LbM2EE5m+TOT1x4UxjjFOrsvXaIShs5ESCazHwhB
Jw3T7eGuZZ7RerD6+Nys94Ho7K4d98eYZw00DHv/4rAP+fKHxdmBe9dlK2xiHIAuDPEMSEhkIKWk
v26pPfvDAB05XARxTTJmbEO6HtVEhdFnRMAo/CNem77S24OtyT99hUKenlP4V/0lBR9+hG4oYuPd
ZDUr3zjhrkqcgWBoUVn4m2ErueUqRqZJkiMGP3yo7V8GbgNp8FWsWoCh/3pX4giQ05ohZuD91tQz
pdrYMR5P5zxko8sjmA0FaXosthPWJw3jdJ8ks/vgloKwCBs7OR4i/d6HtwyqcFx5aXra4yug+YDy
NJdk7JLViah48PCxTvZBJKHjt/8GKIlhu0DeBS+qhNdxVMe3I/LBHIUufaNBHGoppp4dB/z1Bk+/
HBcnZCb7Y7icgu4Oi0dpQhCmahTuzvTZmTe9MYrpm+QUZi6mNZAFN+qfmMTJ3ob3EgcNXRTBtHVA
Hd7861leRAEbSutncw0tPP/GJOqp4XCV3WxWxRxLwgY0/7sSocqIIeuvWehYVQ7xLgV4dzLM4sBF
nHNPukyX3D0sWNOzLm2S9z8cHRYHonHQc84rgNA+0BngdplPyG2qx1LV0LUUhaq6I8rVBi+jPCC0
6slJjNxEOB5G+Qc6d3ByEHJ91aUHw6/3Njqaw9fITqYOEbJgDMdjP64kzYUQr43gzPu82GX9CLR6
/6u7HocpLjbazqMMSa5ihmLyZRrA6V31UYT5XUSlJ2Gnrgmr0TkiT3P/afyImcDu5LI7ntBQduo7
ddaKt1H0LJgWVDr4dGK4Qfr7K31Db8huEeGXo4GN/S/yDb5h+pEK4nvoZml5Vjl+H43oyACkZVzD
ApVrO81RSV5c3Fut2Yt66sLbt1vNgoQQArJlgt8CHL7NzW0Di5CWbUkyRHSorOdQ0FzkPrLwTzqr
nRnaF+1RUX3qREUHOGcWdYUKWcsbSTgcs1qPwaeXY1R7ZoSpwBiYNlmflpmppfT1puPwhpkfX9my
D27v9Gw136+LsqIOl7GhSlAmWWc5f/2zFlURFsmrHeAhsugFudzHv+p2h+qprxJ6+2yYEB9tV/4y
umwZ0b5ooB6/03V+gtVnPvLeyxWG/yl5l+1fmwDp9+0cWiKwMwX7EAFYkfrdm5TIm/rUGPbwjraB
kJ2RSe2s6VPSdYEVAOgPmaZYNJJgtk20VAcrER1ltFWrPlCfqpGq30L+2CpJots6ebGKtjJZHQTK
pZMi2NNIZwRzNinRdXliCwja41FrQ/r7ESp1tHho8Tgw2/mdtMiCqHXIoO06pOaAs221E0JmNt7y
eW8lX774iS9kFrnEeB5J1AADSTXTEkSJrJuajW9tfZR+NzUEV1SdF4nFP+MeSg4PQDfRnW1fU6TZ
Zi468JV+5ovaZpTyEr7UBJBYyopy/O48bTt7wzbJ7hqeXsXREM/DE0qA/rg+HDGQOsls2+6AMttn
5rGxO3kIwjVT5i7ywUMdskUsXOlyINFfVt8oPoJTR5WAdTqc7My4aosRQPJ5rvZEOoptZL6skhNE
Su/oHCffHTbXaH4x/gVyIxZEgfh7ZTdvobWoFG3CE7G/7zb+10/xRFOnHEMXz8YgFAz2uizCh7vF
TJ7HH1cXl0ynWwLmb84T7B5NNUF9LC6rRxsbl/UDYXkznjxK5wudF34CXIaZo0ubUwDqBfRV8tNR
DeoHPK3+Nl8Mpq3jso+/PGzUByH9iZlwYZMFaChXBQlUoLcpBEGpNibFQAMeK11B5RYY5bxc005y
yBCKJamzj+e2sG8YE1/2YpjwT2Vkjv7hF52AsONEkphXb26ATeSGwoo0G4wtSMfRe5Wd1Phj7yIZ
TH7HUBnUuF1hq1CNvJfcbr250ag5lmwa5TZkmCsDNYrXrY3/zEUBmMd8A+uWKK61wqnXnRbxqgjW
npcmGOJgDyC8S7IrjesjOugr7Ky9/VnevjRdZzH3+DgdsAJ6xeu1peD80OCeR11r75g/010R4J9w
AY/HhCICdaQDWxCJOVHz6YFv480pKvr16JDcErodTQetV6D0pGXjNaWxvwAehFLbefsBj2Kxw/LA
fpjO/9kTk3gRJ5yyqYLn/eZbdm6p5+wtX4YvHXg3pzOAIk6BN6iYHpLU4EXYgRXajf8rW4r3y5X9
FektYfqbdk5Lr936NE9N6Y2CXTUmT5TKbZHJ8y3V6UmRSlvsKkDIdOxppvxOflz4NgeeHxvJbtLM
4v1hBnJtTt9H/55PcnuXME1feqyItUQTGMO7zVcwiEwvTnJXuGi3dBNIxLj+F0zmdJKKYXNsjlkM
ccuYdL/9vPCbQivNDb7aZKdpcLaK1fnchd9Y+gTnbO8fwHTDYanazWmfHSq7U3IsB4xLjnH1QN1Q
5OQfOJpUpdAI/6Q2bz0AtxVtPAlJ8H7hHp9BJtuoR2i9ny5WabNqNbIJFTbGr0jn8+TMAFcYs4+n
IqwiQg2yqOTd0N6+3WQnS3+gyd9UhA2DHN9NhBqJ4M7OBePYytgQh/CQJ2xkVoo4eA/AmkV3KuD8
wK1ng3+JuN3aff/PJ8YTWdKxJyherSYIbLcXsPsTe0+hxv90ID6t8KgbOMaCa9rYBPa+QbcFMDhM
RbQ5oWAzEbCvCVsAQZwb8fZQ6FzSwYfD6jAxFd4rE+7GChVXeSGf2u8J9nKMUWkN/YPBVHOOlIyN
4PGwCoOQull09DpJhnvKojqQOC++hAQAUTeV3FGFHl4I90DeLGWHRfH8z8wL/D45pdBPoLzkT/Fd
XPVErgwHlO0aNnxOHLB96F3P1osPRpFst+Go8VQvHL91QqHd9rRG9VqrB5Csstq8sGZPcPFJHRAo
QgoiQ1ZJIjD530a5+yFDsilAQzeXJ8Z5NQ0n/5YDvHEm1jWW49EOL7kcjE4/PRuEWFALX4qNMy76
88HPk1v9JfpYdLBk4yw/VgCVOykrK/Yx1fw2h9hiwsEkz72By+UzljqpZPBZXxPT/hQvaXnr9YKS
W2oZG4UdKdK5EHoS9oBnOpbtkpW10R1yOUShKGUky6gYgGSdtmOwpBQtRYSnswgDYr7/mwPmyvL7
d9F+rabFewh0bp6GFJyHQPcXXPmnCYs4hr8aeA2ZFx+JXa/SDx+D0s3ab7Beu6RZCH3TZ5u66CQC
BAIuS+W4MklV4+BmrHCBa0uzJi1vmiuuF4f6l25X5q83A0iFBdU/FdM7Tq95gsNEF6gcRTilwMYE
gDz+2vxqLCXyM5ghCUE9jTDyYsYTWYYWhwCrLrn/6y9/MtBFBZYCEzCabJkeEvyWPfnX9W+Kr8O/
F1l40fWwALVdYQPdQia2Icy1wleN0Ew83RgrtNFAaAX7oiovzBKbos5VjU7GmMpVkWbupQmz66zO
HdQKwjApbcFIwNjsweb/qoTWdFiyihzWv4EeGkYbKXY5oXVoFgZQ+WFOYsYCMdS17isixP3Ula1Z
3CQU7UQDphVKSd3nHI6ZBiT7tWrZNYkPuh7AH2NlWF7Ez9bJCZES6bIC1YSp3EGGS6VddB2NzyId
1OIzwxdLiuJeaOIFH75Zj4GmLpj+GWt4ZZw/UCSXX5YU7D810h7g2GNxsjjrEeNacJAKi8qIzJP7
ACxFP3XSBBKcqaxzeoHW6ZYGRlI/LbrWjOAJVrQCm9DpS2YH90UgdZhsQ8LjfMpCrZnqqp6AM65e
cJ7t2v0nbDiXnADwMzyXwAkizJKEcdl9lvyUHzLSiA54B+G5cVA256NnsE3Dxiyg3OpppdFhB854
4TbVrHe/bAkJUHAXkYKGzEFQa8YzueHRBe1QYgOeOwNT1duKSHNA1SFwVprc7QVDuoSbmBMjh6fX
D/IWB5AIda2H9NUNCyIzdlSevZB9/WgY/Qdzu45jS4H9KwV2xn4qCuR1AAVYYFxMa6pGTLtGO/GI
jWeb/b1wO26u2HlcmYKXnZi15x7Oga8w4acGmBTETkY4OkIkJh51G8/VpT4GUIPFuHtKBurZPeWJ
ZlX0wODWPJ+MGrusqIsgqrNACPMY9lEvf2r2p3cwQ3A0noeCUzh6tJt7T6d5jgjTU5b0MrFoBfsM
uC7a6RNpqquiee5K+CHyXxTpMj0m9pQrpTL53pUQzZCrBeeCQk9uwYeIbvl+A3BImORGWotJeZFN
UR7GXK/QstGM/oreoZWOOOeBhKzobew/MxVQw65ZjD1bNUhgsK7qg2N1Vu9FVaahzthWjTo2ArLM
gYb6S9tR7tlZqTg6Y/PqHYLpiHN30e+GWUCBKmsdrNV0nanWG+yE3k04lPsekmc6Jfmba4LbtH/h
BqpU4G7xtpUg8ni+nvOcVJTTIz1G+lxvGbcuK7BGw5LT7/f8+Q/f8uke6wlGGhT3ldmGbvu3i1sZ
Fmpbv4IC6xQnd9/kSDoqPJwI6fotkHI3DP6XRe/W5Lp3w/b3FjwjYJ1pQXXyvxWeoUcZDAWKZRxC
dlneZlHnT3IvRLzRVxklB1L5xMQ9NVU/jDE4kehJ/Y4oDSvo7guusyQnkcvADh6UHjvJ+xcrQ26u
FepsIVVQOnl58qLhjb7tlrCGef2kcXVf1WBOdExsENeYgwpavHuCIxYyWCsRMFkaqF/ITiZKTiVd
6JOQsyFPq/Ih1yvEELyj15+Q76yOoscYucV1B6mkzfUYGJZVPKIu9beV9VIPZU7EkF/SdulhlY4t
dk6K1XPcVeUzbeLRh213lOmEyjIr4avYC+LTDdMyQdf6eKuy9PpJRR5iPGxpuVwFsAzeXFArs+l+
HEEBwCdlqoWG2Pl+fBqWeKt2/U3vH4FIi3xLq/sDQfEvoDi08zTzz5E+AldYAC/VFlW00R1XhUrg
m7eBWOOsaY5G0I4xcbXwlq7tHf51O070++RDq4N3t/aBSHBlXlm1dQWI4UJhRLafFx2eMa5nmE++
0yGLOEIlJRI7IzP471SmHDfJ1d59tRTJUR2Ee32wO1+F6t35rb/4VuoF8gTmzMvc0yYQIIVZZCA6
tpk28feiby37ehgO26vThQLLvJNQWeMhx9glWPrY5xA17y364c+od7hu79pcds1k8tMjG357yO0X
dc8wPb9oiNzKzQrRM403eYgRP1uc9nVDy/a4jsE043jOvyLKveMGPlakalwfDVhpykVidT0knrOy
kVTs8K/0CPyAtmBvpd1MjGpmw3EhkMfpzgXBW8GprbCScfbtXqAM7l4mYqUGZII3ErxDSLGJRlns
4wlkpf9j1FEz2kOY/B0wPyeh7JwK6w/2sV/bl9qPDRfDbK8KifLf/EnggKIBVlXlZRZHs4V6TX6T
69sOKx0mT1Lx7P9S0mTl+E1MCztba7Hap/TRFOrVHXCSA7I2JGAjGSjMI+l/ROb9psvNdXiKF1Ew
HBJV7oP/igsq5HF5DhmjvYEDzzO76O7tXeQW4g3qeXn6SapX2hjqlexmPt/p6p4LPEK/0RKk4HGy
0JZZJLPqWmLKMnJDHJzeKnlSUJmchh2tJBJHTuynnOrldCNSw2POzTjOh7kRTskQTig7M10Oe2SX
LdUiP1BethgCXk/0xeRHPTZ+drnggNNDGsixE79sw/v3H+TzbsMaMNQTnYDKoV6/q3tJlDICyh3u
GAk8cVXnOiwzPFWs+0dIjnx7MsL/DQd7EwhYNNyxv6FGEHRJxEzBvAEd2E4p/ATfYM4Lm5JdZQNX
ikks8rrAKbCPrhrBMPnx3KM2FvFfOm9KXbo3r/Rsw4fzlvO+NnaoBOqFr99vWOJbKENP10mC0ONR
NkPplhI0vryvHl/lmYatJX3wcqdG+29IYsKy3qfCLKjTd3PdTf71nmnyB2xtCv+Kp+POVM6DhbSO
WSl1/vQopwKgB3QST5QANKzRi+TL5H5pi7mJhI4zhT9x7vxgfczmRbBYuPj7vQnP93eSzVyokXtw
wpWaeIwSddWwl5yOZfJf6clEjX5BSmqzcStOuWwkI40ocQBG6lobiA4Ue+3YUB7LMvEuGR08ZFjJ
Iwr6TbtrJAuf1sOZuYySqdBb43wffz/m6F8hc6ADnlXseAT2qbRWNbsKZ+bC0Hi+OfjJS1I7gT64
kqqJBPqlD7ZSQEp0SrQO6v3a/KNuNvCpSX1usZrONPXU7nnO2DDQtE2o8+CXCAqQQUKuEL412guh
A3RJH2AHhmTSxOJKilkjhnnYZ50K+Odc0whKyX7QOPYjy4kHoVrar5aSUYVaCc34Ziw5sj6iQYKF
iI+cEoOd1DhNsKRWZVWCSGo7W8dUNUd7rbCK+HSTn/HCe2WsB7IhQHSNC75x+uTR8wXnheh8zeRC
HQwjHmy5L08jC5ZD3VCE4VzEFXqA90GEI5wcE6Mr2tnPHwiOzxiQehw7bNY1tBauxhGa1Hx16h5J
nEiaaeUiXJfhKs/ZXvDqjJU2vhHyCs8XGhqgAoMdmPQbF9CmcYV6CFfpGEyef7msK4j7atgFKfde
wO44G3Df7I61bVegOYwQFltln6Z6U5hqF6Itb+cMOqkhEicKFZIcEH2m9gVDhydwvGtfgvcGgRKi
1aSrYuH1cCLvl2WMqopBDdGujLR1qZjnJyMNKcerbSZ2elEUSnMNmCnlUplJsB0RZKG6w9k4b3p1
FUOkuUFuwb5+vlWr9vP7iPBzOp1N2wWaDWHRIh6sb8JgexWY0LiFXMKKXZzn+Wu9rdp2JpP9ZEuM
L4PYIW/wsoseMOVrSbJwPslixazSFK8+pJ7leNgEyhW3mYdGQb9gfmvNNRj9k67dgCBoWqKY5McW
Y1Y7KxfJaC3E8GMDG91Y8ZjjtJDloLeErJ/Uhwx+ITtOLM/i/MBCB56hgfDFU9dI6qNocrJd00ea
h30WDYXwOHYCz6WSK7+4aWsXNA/1WbIDa4b6o/eYPNb2dpZZ7h6qV3FcfIeVEACxgn4HZJbqy43L
/+avE1mUIDUa3SsK4UB23d6P8OOEwbLxsNfWlb8fE5Zh6BNplhXTQS1dHtJvcKu434SEIozw3yTY
w/jRGUitwvM9plT9f6PfMtNEnfEAAbRKpgB8QKRj1zIz21I7J0mkw8o4TSjQzYlfUk13s+j4jenS
kxyYOkoUl0aI2llAYBjKYcGwHvbxvzZThx1ifnjSs6l/BmBiLWTLMETSmbQltFQBtAiPwnTj7rPD
Iqjs+QWiyarQxY8PR+BNjILUsYQVnomIaU5x38kRWnJBh7gOq8a0pQeXgXGAKBICWRs5tZf1PMK+
cO/2lbHXYVHoUKvtPJXLk6X12eeS1bh7y6MCWfkJCcJkwBGSrS2n+lpDl5T57ZbdIncxxbDj5gTn
mHDCymLiHBOI05s8SuG1i3D6j0cd9Ma4PH6LRAIt4sDWFGXT8CT/e7eUMPVOw39WMgx2s6mju7Vy
qRqxAPtPaakaCORgG4vuTWUkiS19GiLVIWqa4xXJNEj9Oyg9yxeWh6q0aYhmDIYA/TDXdCltRB/F
FJS5MhZhdYBOw43N2fQQFVo35CLNqk4GfxaMGIC2/V9kkkYyxJsEeGuCLsZ6zRZW4CqLYAoEGoVI
3gursQZuVuE7JcZWWqutrX/x6RhFolybTRfpThRTQOMzViY6pyrMV+MvrlsHtRdWAnmzquwmgcyx
p5VLMt7bexiLgGbLC6d5FfXVrSNf3ODehrML0rYz2Pl/golhcKM5P5MJNDKUDobhkLA8yCidbK4p
khyKhbesyiEVKoQ8Ujme5k5V4OzJG8muB1T557wRLc5FxEiRDzuC4cBPDfo4kJCKK38l1NY6D9z2
SX4gv6wUNXi8Wqirx8nd0W3Ddga7sPrIK1QOeOeU/G2wfILonb2AiANk8/ykQ8dpxD2dhWKlev0q
TRaT68czSUkaG2XeZ5PHcfoymmff6dCofFGKR0vALx5yEjyakgrW+d+gF0rZ31PZAitywNb6QgqD
rW8HzOfb7z3pXCNTwzxx4ZTz9LFic+gH64nyTWEx8cy3shn1FjeDo49HWjwf4Av/cgfQZDUg1roF
ctaNIUR/MVx2vggADC5pxZFwFQHbNvFHQZiJZJtwxEFtqKsPT53a7GtFANQ8Dhg1tRGf+b+m9RRG
7RDwg7RNdYney05MFcNJUM2q8qh6xWtTGZEf8bqUn7LzzXRB6BPNCR+hyVaEi/Q0c/4/NSPbIdAJ
Hiz5sEe0OiKcp3gzR4/XnX/DoJT8K4OYI357NVYDxKP1EEmM7cRDKwFgKpTEeG7GxIdk+v29pG6g
J2Ga3jUq/6w7qteQdzbmxe2WIa0d6dNbw054JQCqmIz1NRqynhoaN/tGKEXy1NKAH+SB4nQO/Yve
N6RX0mWrlKfN1bW+Tog5yjitwaNbx0xePVLEEK46h9hTrnI5WrbTEcuCkDkPMcTmFGibdLirEEgl
yQajR3jJXgMxzXiXCu7lxt3/3BydqQ7eQzQKEqUEjiggRBuT7gIAkWIOA8f+L94FPXTgMQtn7mCj
q79UQX3A77E7Y8/Id0tNi3M1rfYCB0JBxdDVab2by9N0iGYCQ2riAfyu0r1cLOgyTU48V7eKQGS0
DogE2HMSMnEfz9RTXWhvTcFfrgnQTclFdQT2EfNf33GnD3AGghqJtsWIZIc6oL0UKtjadgh7l1y+
N+CPiIHeYYwSdo/3zKXc0Gesmhhw4oj7dq65V/Gw+5OSJiXQjPbJHBATmvUSXXPkOAITymB84E4t
M15pbvb08QUUPNMaQj+gJlGXrtH6/0/c6XcEHHcLyHzL8dUgmhgHJa0GWKellYD9c2BjhPbmvNPa
RElX6L2tfQ14oWrCAxMfMRtDk3npKg4I5SWCbb8Nc/EDfd0G8eaNDTt6c2Y5qVNrB2RQXy1COOPb
E34L5sn0PDehfGxd5DSG9ZGF6cZVTOoNzmx+RCVCNwJ/YDeF0qBid1J8d9AqRWkSLYXo8yn0ZgnC
JY30l5H8LDlYzH+9khT/BZorY8TJCekBfv3eWgdbQZLbJMPgMLS9FBhyRX+pdAFGkhFdlMQkVgKn
SzYqXpX7i6FsNa9xoQjx8XVCE+mwvfbidZFyGdTiL6RtqT7BEIWsVbUEMS8tPP31Q+OBhS3YMcY1
fPzYqYGCitPdUcXA4rmh8WJHt+yvYuIDPc+kM/fYDIZUC6pkk2xlfIOkIsubgNeXgFcvZ3jHVe3z
NscGFRo+hb0ylPkrZoJSdGzVetW2Ag4hSDWp4OqukgRoeY4CostDZGaEXfAFzNlJZN7uEAaL2Dpb
JvIaYCQyLN5Dv071aBhMSDa3wUy8++j2pZEfh66mj2suRRXUz7wYOmt2cLQBIk4wSTQafU6yYgIZ
peozsx8nlybPBxlE/il52JFrNaKMXQhtVSWNbIA2VTkxJxq4mJjKfy3KVn4yvEH0bjWJnKhu0c6s
7c5qaevUMFZJ7mllJZo3oye8RhXkcNuuXUsjcmes69F/W9vBNJBOb13L+dCPuZnN36BdUiEue9JQ
MyDlHVAbbcl8hQ7+th8uX0B4/Hl2Zf98WXl8QMDu7wH7KxgvLdrWYEB+WGB6fLGxRyCsxpXFJODi
X07NHaOy3YD0bHsuFlFVgwD8lj94auNijenA9XGMit0f+CoNRabd7u4P6bl85EC8Aj3dOyBqXPmZ
KjgyPf7xnfg9XaBXKhk5KP5yTqqgQvCH6HG+Eag3yQcOT7Kd0MjwJGOhG8pqGLlG8vK7hxqs3pfQ
3lAlQH7T9fzY7BekNpgJsvMNJSdnSFDEisufMybOlv7BVM6kfuvJ6SkJZtVhTKYZQuekj1km3vX5
K1Ft3Sqv8LQCH0y5tb51PSJ9OM0fHwT7Pf+FoykwVoC7sHDu/GZ7oq5ZoOOgaY/WjyhnqJBKmkHy
rUcbH0MjL8OVKDQQdWHkMMkjdprv6UlHT+M96gwf30A6iDaZwebanTmsxfTqDVPrvwJ8bFPUQ8JC
GHpCemGQ4PpjrRKmIMuCI7Q1tiXzYWprr3r8P3LOR1Zm0k4jPA3mgIzzE7cuxwPuT9rnxqc9EVvx
f26cg/1p89CfUp1t4ywzyTYq7aSMkDAySmm+rXD91k8QHNE9c88nIyFpxplaLPL6HjJCYFzEJ6kF
5rFiJLvxQCYVBXlYo2qjm+FvPIu9Bely1H8cE78xeelfbEfX6X+hAX05GJZWPGeIAxupdysUcLq0
r/0VXwfeopWrmRyGNvQpnQ5NiwzR0ciXZN9DydjfeWNpv1iyj8xplEEhDLqd6Vzt8ZHjjOIlDDRz
G5oBcIwP2xKXEr06/s8FWGOpbEYe18YBKveDwGBzeOf87vc+mFta2srGha9xqB532Pf9snnijEkG
0b22nmINN8jf3wBfJx0SkIt9k3YvuZsytqh98efqr7bd6qevRy0Qvnf0aYTGv9rxcpy8dmpDYPG4
nD8MBo5YytO07sMU6ma025BEM1Z/iasPjkPq0h7S0roCjLcjPG6nWkeMovEplfMh0UINcTJICGY1
HByWAM+h2IU6KoNvMYStoMsdvoYqY0BgxYd8xeXH4E/+V2R13GLSBLy8EQx6znyvVZMSofLS76EH
DZkc55Wd8MZZQtucmGPSAJslnSAeoF/sn4npGBMVkulrf37SPlFs5rSZnIPQr1Gq8aMVFXv9l9+x
4YNIe/vjNkw70MTwP9maphReU/o1P3HnedX38UhhfhyHkC5Ctuil5K0uYQ3g0mgrnM74Sp6ieyN9
+0qI/bO1ab9Vt9relkLOM9IewFk4uSWDRoDSeCAbOEJboUvTzrGjQGLc5EzhjaB0paPBjAiZHbnw
A8xp1vCTOLOZd1sW+ZJtCzvc1TAKudY6lO5mJg4b7rpK1lRegssNtDPinKG1q1PIe16rcL2Oy6Ms
tgPBFKdcZPwJRzt/VL8yHIp1q1OEoNubYsSeIBVdSzSnE9p0g4zDkQFPdQ5hmGfXY3nf2BU35eE2
ut1HYdV+r1l8PmzQxe1JxM9GzAb4RlHPaNAne0NJkeV2EbKSL2EPMHTenXDOVoY5aEuKauNuG1Hs
GdnHho8YUo1hWL1LOzrqzV+bKKh7syt899nOw1GKdlZg0muZjTSk85mL6wYmcwPG2PGb+KBg8fF3
ww95l5aiovDJtRdy6iMwwb8qQCPTALsjDXnbgerRa+/UUcP9BI/jFVfL+spolnyUgMEp97GOItV+
JNv2fkeY1qP3JHyuKg9p34UFy/jerv/rmbvCdbTx9fWFVMvvC6HPSXd3XynnwRh+dKzrPxZDxQ/6
QGKfv6uvqgmY3PRGNK2L6WnsOi6jd4fN+q8a1aLDh6AMXV+jW7kIaepT2ibrnaPU/cDyMIrSXGAP
7fx/eFb+zKPVuCAGe2bjchs0Vxf6SlaHjJIvr8Oi4OKEMlxN7zg8tmJ6K6acB1yi4/vlp7D1isg4
46F8VQGyiUboXiOr5IpapIiN3YEJ5e+Ke9YTbZufLWrL3B//SfoX1M8FrpgHudsLbBgXwQp6/mXs
H/oUnExB2Dhpe2wU9U5evncXzayVX+CP2wTSGvfd7hdD2MwSbJT2bH+8FKfw+dkfflq+MOweS+Sq
rDf1Ido2Kza4zOWTUx8esM15YIeY428vzfgtPXLlzFjgFmtDgZdN2cs6ffqguu8JrljnzUnqwbbT
IhYAXSqR5wksZ3ClTWsacIxhzcUaNVzj8x7ezvQDS4AekVBIGcMfRoW8MCQYo8fJuYsz1IPLfUCe
s6L0bhpjJfLVlkkgyzmojoQM1P8EX3vymKb77E2awLRgRh2sAmF5a3ukqbbyoKh92N5ZLZmVysw8
mGe/kvi0DA9wCDBCjhpnCC0Rd6LICUH/dLYJPA1LnKJbnnMSgNza3FKkppyVlWXmpYLsDGAhyqKl
XPSEUVcfDTjXqPwLKWP/izT8qiQUnHcNkY913qpujpCcg7Xw9T+DZZpVVL/I6ISB3dmbN7QHfA34
1BvMMkyIwytNJNDlz+AnJhwQPtgIX1f42qjsbf4VrZNaT2r29ECZGXY0GL53jK0BimCmr5zXNJCC
zBC2piNmMFo071w7tdgPNSgXpQrd2z5mY5/YhTlJioGgRB6LSJo+g0gnHyf8Hbu3Hj+4Cq47n/MU
NMK0p4LrAxuDO4lsRdYKe1x5630RcKKDiK4abHVoFH8eiC9rMir9uOQumaHpY9LgWM07gtNTzS1I
XT29Aa9zS+S27RYzHZGO6lmGenheUltI3/cZGOYJnxT618BmsKDyUK+WYQcho6OpgVm0YvUbNPnA
8uf5bhGXZKTgt1qDmHrSfaNN5jHTNujkWIG8bof+JLXrfE1DUecCNgPbCakjvHsnvfJ2a0+zBL51
hxy1+V5dwHThfj3vqsZiavgLizjwtj+h8gir+zKgLuMfmhlDXrGz5OCwxEqJdTUB8wS4vFgbpiL5
RzG/TfkVfqusHRNROhUSw4u6RxwIcNNy6UJ3y+6+VDHTtIVCn88cP60GI9F+zyS/hfTa3/zLXw5z
j1uQcb3MUq7aN4IR75xrdyOBJJilUO6JMeFnMZtL8oQt2moydoXGpL1aXW8AWj3xT2vimrKgmWor
q6DPNxK7IZpi0m0DPtLsvKVaFnztl/xnFhZWK5VnCFzj51QC9Z2B/G08Ov/yE/L98gqn8m8moArV
XnZMZeFBIPz6u+T5AnC52zN6WbX9gxe3HGr0Dd43XGRvkOfrTbnH1A2lVCrcZQ37soK7+J3LUETV
cY6/sV9qNfsQlCCpe7bw9dKf5Zb/tJTlA7dLeoCGIHQnxDZTFIcnXilSnfbqaIVfuH6IZ8VOOyNW
P1XZb265nsYb2TMa2ETgybLIfU9Ypy2+0GNuuygafA8XfmDIWZ6WSJFj/ZxuTq5TtRKRwMh4Pv+V
S4BseVPUz+adg30mnthPSeJSX03xcqTJzRyNRoHdRIC33v+jwQEJSUzAKM6z+UBJR3FvvgJDXfA8
BWLd76G97BWwKUuxPKSD6mXKlV11e2NjPDdphRvHyfseTHXgHQG9S6cXobfyFN66MSVIJEKmrIEh
5KiLBaaALvW/sRLYj+nOgORTjr0VXSg5pfJwzERqH2RfBPd/yd3+KiwWwj/4gXoQeB+LI93wHj44
inzj9Q+giV8ZuAbDsyBX4p/+9p3757s1pavZep0/n1d/u3ZZX9atQvGeoeNV2YfhDNGPZMNjedeO
e0a6n2vhAos3u4Z9cfy+yP7w5RdS7BdE2J+Q8amNJdu2gqFIWWbXx7T6vmUEvNHDJF8+Kq2pne9X
YbnpwuBZAhfkY4UTtIlidypEU03tiytwIkbhgkAJdhcVhCoes0io29LgwoMtEmpTSboDCgGSbJX3
6weSsXY7zaDacl3Z8C6VC8NDZH8D/6wgjq9dV6VtF75SihUJexclvQVFhmhvW0cC0Ca0QIHe4nOR
Jy6ZAaMIC7AdLHV03ksaGlEkoyViuV0bxgd1q/twd33XmRxk8WXWQXyzi9hDpm62z5p26vrJrT/K
TsbrxOSWhwpENl9pxziNw9/+hw4S+uou3MsxfMG2eon7PorX46GfAGI6Yihrcc7uBPl9EWY1mDrw
cGVh+oJeMiCu6mjFMHYdT2ApbhkPqrd7PqJ8BjcpJnRbjSRpAoUqDdz0Q93Z0ZuxAuLApJkybYzq
XA4vDnbsarBVTKB3pDiYW8Zpd4TLb0gFgm1yxHTDKZFC/RypVp6ObybW//U8I7RamC19G4xCvwES
MWSPh6TJ5NdBHlj+uezh88txCTrdQhWLC7k4yhaiG1SuIx+xlCyuOUWvdu9r+ehSDuujESFzR/S7
wIhwj5Ao9aVPCdr+GdKlG8PJ9aX0iRQwosLDdc4kpT2SfM+Ech+o9tqwIpTJXre3Z/lbmQDeacks
+PUxOqppZ/4vhqd8uTBHmHtxP9Q9T8RFoomdJegOO+JgbKbH0GgrJm5saIbneNpCMAG8VvJzZreS
HcSevuPkYBu8X53seTvRK59x4GXWNA6r5rcQFqbCXBxBJ4g0lIDhPnLqx9RHFsdytUSIiXo54VSt
dMKUxWXNm7QRPALlnAYJJVa1efQffOKUO2ZGho3yg6D6YD7M8T23bRYPRQi3+/0NoVYvNmP5i5Es
Tje+zo1LfVOACWoZtH6MNoRDvh8w9GDhrw+dZw3hKP9U/Zu1BMGV/C0cyLw9FQNa8bBHbX9xMN5p
n1TO6jm/btBKLDSyPRmTaU4QFXObkFeEiOIMU3JUZNNB2VwwjPIaVC5DLL0UseBi1U0rzUV37ICT
DAeWyf037imO6dQ/h+N+f+56i3QPmvj0fF2rg4ErpPyP0Cci9rpvk1NonV5TzsEKRgNgzwVSgPA8
9TnkTB9wrIX6wrE2Ewwt+ZmKpPmcjpq2KDkk2k5jGhExvYNI5CEexkNyMED3uglnGWMKMgeRiGMe
1PXcUqKZpF2+xVGakS3rrtNCf5tsKfQwCwdPrHpHgo8aCJKv2FQw060Z5mnbfSgnC4RdyrhXdWM6
PW2+PuFwFthvSCPSmQymVV14Ot1gb9B3p/fQO6ynt6nhQ/IAknhS/IEhTvPkQVXyWXk9FZvoF21V
MZVHS89Uqp7nCkxoWly53dVoTJ6ScpTfPc34llA4dezDug1iBXkCyRYRb9N9nFYj451HdKQhEUJD
P4Qgeod5wEbLTVtLsfR+Qc1ZMerAUlSkiqH2GxKPppALiKQZ8AKS8Pyxd9CaWJVaomIp+uyISl8S
c5+PqmpB+agy52MBmSr1ilF6/DR5krGSwDznSVxzCpByHqPZuUME4NISfqIBFOFti1Vnw9u+DBCU
ILaVnZygjDybzbUSEpt4jWKQ7/tZZ0QawQLfpzxbaL3w88lMUSqU+BrNPt1EkS7I48A7q3Kp9pxG
i6xkKXKg9ekgXY0OtuSaghDB/s5bLuZhSHsqFmAzg4SqXzOgFlnQz47tuPIlGoXoUkoL6UHdbvLr
+Kvn4Zn3O1wgMk9cILc0GJcWC0G+LV0EUatbnAPgtdB1o53+q6VRyyVHkuBagyLpAqh7gzhyb92K
TpE42AkASjBH9xDtAsOwfzOUfVxvraeuI9pZ8KVkNeXCBh4saSx12P8/8NPj2ffSVDCjbEQ4wBfd
wE1LKVEp0JkSwz0Op9BueKLIjChfRJfX+73w4UtGXCobR4BsiDGdta28M8yBV/592moiUdKfOWgi
yc5cNyruJv/2kZJ5Y0eJoEFQuNiPRs3epwk+I75dJ3vcwjEQyjK7+GuWF0mTUhMJ6Eizmreh+LBw
wgYJcnu8JXsfFvYS8jgtQdZjVBbDTU4P61zPKplZKNnSwRkBBRrGyiddXVxUWlWLuHpuAc2vS7W5
yTfkoTEthmsTAAiYjjQsWkeyvc5IhBWUkZ62P7v2Hwj3BbrcoTFg0/j10nmkoe2vqMlGezg6fvt3
pz3XriLbmtURnQWtw6GhrjTvL+HCDi7DvR0Nz38OCaAscl1faKsgJiWBBzyfcl69v9RTDNEwjgQc
l33o4Cn/Si4/wplH44HnbvhaJ36EhHw8o6uPoF1rGmerOkZs1cvkhJXvxIWQXsUJOsuDbRT+eQ0k
J07V+gW6qSMc7Cg5j0SARcOK8keitY/63KGu6FEDSjGs3LjPxUaFNqn4sa26qaPLuxZR/flRXgos
jRLDaZuzqxXmw+ZDAxOUg2JME26fe1SjCe1FLyFLZzL1dBmsfv98Jitc9ctyb7rOIEEUT+23GQWh
XLmoVxiKW3T3mYxutr/C6x2r0I42/xtwJc1husszHlXIDI3owxBuYu35UrlCFFzlBg6XblJy0LGH
alzKZX1ypk3cfIqcB59xmLa/HujBO7PyM7CyvoNCg6w8nHO5k2L1uCSoXDP7rv5CLGcWWzwnqru+
76DM/Lk+tTfSK+y3VWbJ6eG/A8ftjKY2Ln1ZqZeOXz/OmD1DKBKXvyThsf00xFHMt3OY3Z+Jtf3n
nZoU3vfIjGgCdY7PkvL5yK+NO6tBUHAB089RP1hBrGfBSwTtN962e62OmWOKzcCUeuMnCetk572c
NyD+sD5AVyB114R5SobOpW/nKK01Ms8b7VVt+vCIpeVCh/YcGfRWuMFNcuTO1/JrM9LGXQx6YbCz
F69jusJ35Rt7dZMw6qpG29uPlyuLf0sukOIKJsxQCyeGTk9p5kQBsAgxXpEi5a169sEXHJI4GRgq
6uAneOrvrwUTYzXPNixtt6EjQyfTMbZL8d5BdYAkbTvWX/ZEimnpKRts/uzpxfUkqc75h1ERWlCS
ysCiOMX6iQ2CHPOelMTmt8r/et/Udbg9a1cN4Y5Ln3zv41V9CqIt84JHZI6QbNAUomA/sclT6m+A
lhgy34pC5Na7cTusZ7lB2ybPPuo3Odc/eMa1AgIAlP3qXw7kRek6sL6G48lIwU8tbxeYO+N+PvhG
s4MjTLzwu5ylnUPxiLH4f2BlR0t+Uu14c81ddidbEQDYPfbi21idBCasDiV0kc4dTqFEG2hl4QU/
QdWzjOVHpIsbV1RstmcLVPpncXJLHOWc/fIw/7LdtiSTqOUzKWGVdaqd36wOLLpnzQbAXsA5UV/Q
NFjN0zP9DhCiAEucQGTt60wzm2/fDZm05T60UZ2aP4SUI/vNiDZI5CQliiVT3gxe4iN7OXXVX9p1
8xHh4tfELadsGoWunc7QZl4icdK6ECv7tHoyj6YwS/OUz/zDVKNtmX6UZqcVn4lF7FolLFOEREec
qes9MROm15GE3DClLH/RZCrwxzk0qtaeVkuG0SojhZfaSu65yucqiE6Dff7bgCJEQFwrywbGFD2I
ndpGHADaojbJ4L5beyaUAy2TTO8EinZKXi0fJ0AO743d+tc2mpIjcyHkYSt4584chlBQWcRUNFp9
80hubkz0kezmzpkWqYt0FEvBeT3vCEQDQYxNWY6jE7EHscC2fT6eXkgzRDZDrzUaYmvY6Rg01Tw+
nKBRKeluPW+ux8uLED4EPFsUdKIJo3Cl+CGNeemstKqRAGJZMRTBSx6cmDOHT8h8LHkmGUbm0gN2
Pttn0TJEr9kg/Wxh5EGqjONZdKbVTxAVfmt4EwP5KQXG1peg6dH77F39AjRtY9zvfwoFsCFSKF7h
I6thEnq5DmccNd54FXWHi+MbxyqeodhsPm0bbIwRg2NQYiJ+TCF31EJIwUsaUxpZj0923p3a958W
DIE1/tBKaQN/LFxVYEasEWAghrL4HYn7jKtNsDikSX14czovJpgint1wUw6G/jjjaZ4ySpYTR/2a
VABrEZoMZTcPl4FhG62dA4npM8Q8Xep2vUkGcfjqGGdzT/PRG6D13ldHJN9AcUsf/irIrvHxo2+O
kWM98eziHhd1RstbRqbhUh20VEsy03pBiuLZebm0N5+POLyNC7/c6Tuhhttyrq4DWf2+dIRiDMeD
/eXMAmE4YW9DY85G+y3Xoanldd77Lmn3bFH6sW/YBmeHsPUrHsEvXP/8p2FdkKeGS4WmwvlEJgVq
KavWD0rSPYYpEcH4URNxSuTzhFMVS/+Y6lj++nS6k2FvDAEj5w1OZPGQxD8nkuhheJtHGZz+JcrP
NvMHkgPEt2zt17+L3KvMpHRI1nrjl8LNetxLNxArVQJ4V+kgZPeRhsH3bKoaKwxCScabwf1hI5K9
WUY/IPLJgxiH6k5m80wrQ3/Z9ni3BTZuOSFdxM6Bk8avb9ZWMfGALAC19oNePMZaumxCXLUnKx8K
qn0K0+EWHd+6qtmxQXhcItRVpwJ/bEeIGNAfyKen2mzaxo+ke1IJgHVDmATLFM5ykdREFoYk+37Y
NjgYu1f3UxBwv/6Cc/X8MKJigNRLib26SFbWlkQwsfnPHjGdrTu8ujMaKaUajcRppKwelZcBlma8
+Q1f/0kzm+I3F4kSFp3V8QgVvi1jXfbFMzelAGM851S5Nt+KXfd+hUCXuwdE7Q39/AuTZCKEoxdv
B4YJrw+9zYS6k8JQxIUDNckCD6bAXsJSSPQoZvu9S9XOn/zv6KBz0nQ8gmT23OYu5hRhOdB/jchI
v8dZHrK+NJaoLH5HLPxuWL3ik1tlQDJx1GB8tTH3FTtcMzDKW/YiTsjM3Dg8cee1OTsbiflk9cmd
dZvOd/GCrKkA8Lg02vLg8fXs0zSwRpJXlbirnwOAFBx6LoCRtNNPva1S0icujia10ZzT745r3Rbc
2W2Wm/t21zkGsz/3CI4jioNfjgYxaO+dq5nyebZa1uthz7AKBwV69/OKT4BR74gWHPBXqC0TfdJw
iPeMpZEPq7m8N9i6GZqVPMRL0g17InYVOQoOqNzqyY45WEjb0MYTPm1ixNo+v063CxUWYQqNLigx
Ie8fsyW/hZ3BOes+1SNyXFhPTGf1Q410J+G8cBziWermEK1SPvE4lY7Iu1spIr00E3YeSgkXqWJ4
w+MwXKkqf2OzOF6HjbdRemi+16rah2x/biXw5nWSqhQmFoyRM20tr5frreBXr5iYyTQLl0rRXZsS
ohEOtrGZ0AfMoadLAsRSTTxb7Fu9+cc2i2QxcS0UEt6h9L2AX9fytOqoOnFaBQpIR7lugBrXLNdj
8CSrg4hKRopIVD53Aav+/7MALK4wNOi1DNyuChbM4KFIIuxMbu3mjKP57EyjKH/MbNjK9n01JSkQ
OMOp6rrv65lBvHcS5X/12Q29rlz4iULShvi97Iv3KNG84YqpmfD0MMa1WNnQlnGQYgdgZaLbNRh8
XMouyoH6ZJe5beUeLq1hR4IcXIOIiCBbcRx7kN/l3jyn+3yrdJXesawhKV8ddMiUY11Dao03uARE
URsonCMWTWdDA5OtUwkdO0RLPZWdan5auWXLKzlhjp8to5D/JDPE80GsDSVk8Sxea8wSKBDwJ+xK
nJlEnIm1Q4dhNwpUq13L/+J/fB8heuXsSFS+4bEKv00erV9dPtGhG/Y1BPUv2SrDAcVlLGt486GI
HZy72gkU/MTbIGDMlV00+y014Jqpa/khRI9kyzoVLlF+KdsR3ddZZbtrTwfuCfc6X7EtYf/Y+d2S
GPPgaqK42UCfEdbKenwPGqxjCsfcyi250mcTjceSMfkgnR1SGpb5gNhIVIdQIYd/LrQ8eF/JyCt3
qP0dFDFZgAQtqvgnE+fEuKN+ivDkAL5qpZuHIt5abAkORSeHPxKgU6wp2VYkn2ZqcPmvbdUQDXWo
uYXHAYbdMqjm/OqWu6ga0Qqv+KfazQy5zdLaNTZHLnKaLKrg1BMr5fJxFFyn0m4srHnpSofq6IQx
l4O5xZ5SdCkOpinGqz82yNYh7fy476NK7ISkSAYzkIe38DIOSdLdoZCJemxDudTk+Craj7TLO8+1
/TktTZqZn/t8Yz1s7CL71rOUEyiYHou4qtO598Bqzn9LsCmYfta/3sAWhkeOyJTqBJvxOcDw9ryH
sVIFMeiCm2Cz5yzFkS5k1jeYaAp+/vTUy2hfTrIIyq7weyZqErY0U7mOulU2wy0K3RTObYtbSbtB
K3bnsKcuaQOYn8pbDi5dL1kZC8wHb7U/zRtmsHWzqv5TAMO0WUohzUvNb9QLbHN6xmG1+Gajryml
JzrkcTrGeN3tU6T4+UQDmWTMSv2hTBRSECAox37RIGBbsBuHYy/whbXU/w/Hvl1rLepd9ACpH+TA
vue+AVbbhCPyr8gTLYMWal8lE2N1OhRwjQ/Jdr7fgyFiZ4MwqFXZhJml9/Odxrx8ifDlT/DLbGO4
yscCyL2GBkw4GAWpDg77jyjH0UyMWp/DCOx0aP3CWcV5flszLba/ZkjZkjbY4ixxb0g52OxesYKy
ZU6u5xKK1TWyDJWHE0esdIolLo7uJHVOoGrtvFdKkGxl14Rudk1lIxfU3F54a0TgE8u23C2iseDM
ECeghx6M7c1hEKktMpJjWddTUBymki7TRJilnngBJnXFNfefFiPcjpXhGcEDFzISNBJl+X0Q3v02
fipCmFYo+ep54IY1O79ZcqW5gh6UMLvCpwLsrVjhEbqeHwa64eKKl7NPXmwa+u72zSqpLEVDzadu
NFh8wpvcB3oCyW87eiCgylnpXzKa18Wj1uzR12O1Xtr0/NnQwiMn/ogeJxIv0chLGdDvpK0ZPls/
Bl6iBnvyZY0x5rV+7whVJk/vfYTC2cY4/CVP22hxUoln9sF6AwUDlDpgamTIEsXG21LONSflTuFb
nr8HaZuVoxZRuRM4z3SoQOdd75ijmaLJfnYvQ/HHI6qbaqmvLLbGPlHXpzvjmvcu5Kt7uuu8Y2ip
/CpIY9229hnDPgvFnPT52Q4ajoaaY/3ZWsJK7R/oNLwM4K7eMi4w8lrsmFbag7Np8AdV8KsbH+OV
KPhYzeiKSzD+RE42ltME2Za6iYV+YcZ3Eyr8xy+la3Cqfqd4ueLIvLO0sOQpy1qeVfcu3dNd753/
ZC8mv0Gkkj+yRCvSkRP1Hox4yeSv7a1NFEb2gu4YO9VTawdEQ52jdwyYDYNppOUdurYtyuQWfL3E
d2OsxMKJORdj28TBd9iP1wIQX2M7YiR5a3MXE37/sGk5XydHRK2d8bD7GRcySrv+reCHSJH1oRDS
2WiuPELXKvkFv9mzHiOpfq/yXEIVx4/ZhCTo5WHD6epkLU4MN6Bs5rxxKd9y/S90e0eUfdrzNZHd
oek8DCxUhj0LiS8Q4iipvePV801qZrtv54sic13POpJB6DQczv3SGY03+q7q6Jae8X8hmXpJvKCm
gZ/HPq4jR1n3o6ol/DgLo1QIbRQdi5NinuQQym130tWbC+1V4rtRaMpPbFCJqy2T1OrrziyfaB6V
YE/+0asghBaSc2Khk0+FS3mLAv8J5siyF/XHuBp1QQ1dcA3sVm6mYvdcTn2gIQhgusEWleu4p69C
SH+WQKxW4diBr4UazzIToHqVX7v6WpHKxu0GPPTPipfW0AeWffMZjY3WuIy8wBB7rp1ySL3fZUqt
c9yc5Jk2XKE9QWhCwRJ8IA24izDY0w8lNqJ0Mu6lvZV/kBpLQYGe4NSROuo/IRKpZleyWy9amE19
dyoZKSMhMqNtv99ruDHbvCgBLto8RXGijQgNQF/fEYHA99MtACZyJzXnpuVeNo/7rmu6Mj+uXNUD
8rhU67VkUudAXKQlcpHWxoA+jdR8VT0iffoTbCvxghAorewctbtoTQt8W3pMvQdYt6lGhvHXgjS7
4NTbWqI1VXUQk+L1qYgazqzODM9SFmiMhxg++N+QhwiV/55+wG7FYxLhNGsmeElRfKg/IBYfuRRu
wco6gqTLWdgvqZ68LhVX9rUrbn85JqLV+OpIKlbtfNy3G4USzOy5cxqUN0SHO+MEhlQ1c2Wj6JN/
upuB5q1qoejxexS2U0MO7ZP5n6YF4rUozcCgAPBzsAnxEU21G+CLwiQTUXu5hJ6112g7uVIw19zl
bFc3q2p/PYqiHALbOCp8ToPZFSPU58QZmrKEaa2nqg9hGXOsAyq7rwwyHTRZ9cfkPT+iI5631t55
87GipFSio5nXDztH7e9r1831d7lJB8G9p00R5hzisshYq3bPdWG8S6Ig5rJ92DsK4XtDxlOzzbu7
Fi4L6S+1OpHGY+eBG5/wVDEme8gfbnOz2xuJ8KpACKn8UpQnkoHzyBwj1nTpNg1tXtSXuzbEQ4Nk
2qJ2h/0H5o1V3d4dY/2R5+4KMd4CONdOn8UPhAETLjnwJRKaoIjdmuY4qfHjfgpMNOe4JcVefCPe
ORlT82kFHhRpX7SR5OTSpk7j7i+vP2DIsG2U32dO2P6gYcgjc00Z47GK2jk3zhoHeIiA7xfS360o
ZALLFmBow7mA4qLvkGyfkD8GqIkDBUcDfNyAiAX4bsvuOTNTYt9wzjPf+J50HXOa+ih+x1c/TnLk
egM8orPzCtCAUeTH72RnvMK4khidDscVCYRbwRE3GJiiJCT+3a137iwskHpJCpxd4kedt4TdawDs
X5Za3wFePofb0au0klpA17ZdkPrGyizE6nh3c1XYHat8bG27IRImLya4ypVixWJUtl+pj/w7o3Q5
VSjKBu+oMQc6uJHhwDty0PuMgjn3EZA3ubVCzXlfdhvuz4H+qojPbNXnW2YjPklmcunSHVDpNbQ2
1ExfiQ22HeFBjcFOVVGfLzW2urrRX3M/toFxLLHeBl+IoAbiKig7A+YSrGTOPgjzUaYcGdRQTeHl
f8G6GT66ZYd65tHD4r2+6Dw6FPjaeimVu23g9lsyq2iQizHs1VqoUQcnRL8ICxoiUkcrVOCDoOK2
6w1Pdv6ZluyUvy7iniDzFZ8ouNOB1jWFUMX7etAsqlYeNgWwuNSNBRNaZSgIanjuEIfpD4NPJnrr
E89Z46ArWxdtj+FPOU3O7kJL3NIX5xcWXFbpuC+HindgVPnij7v5yA7gnPT+4jr/oIZuz02vDSX1
7kZIwmdzUlxLKwJ+srQn6S8T/ZpaPdJXUfzs5wg9BA6hU50cJFEBj6iO7dfvMsR9vIlFsQrY8uS9
Mgr+JOsEN6z/b4QPL7r3l3t5VfKnsAuxoIUPBLrEgNKDVBkk6u7FlwMrl2eRH4zuF7BM+cPkO7wF
31uxYtgoF0PKk7HA/QrNnEt0i6GMa1pvHowHXt/xKNt4yGTfD5xOcjXstKEpxs0EwwVmuLYC7xr8
luj4uxVqks2Nkik0tr0yOBb6eYHVQlghSOxIHL+TiLmUwLM/GbUdZ0fI2NTPA7AFAiz2EBTaPW1x
k0qz6nJ7OMUlwjAz0dJQCz0fjkxGAo/VHNAhKJiiN2n1ghUK4Sp6tYBMA3tcp9jp+/Hsc+GA4F5K
zIlQhyobKsGYy2przurBd9Mlh0/PzU7WdrACrBu0G5gfPJfHGHWjcvsKVcWlVt+mwWU2K5XVu+5m
QX/eF35ZiEMRBuDgw+snyct3Z41Zcu1yWk3785iLXKLOKNNTwT+fcsqBmFELpV21G2UZflbYYKdW
31/jR9ZADhCabHmD4gxOFy08s810rqZPk82X+ltiMPckQ9xz+VOHKO+im067BdZRm3CDaLFGlOYo
MTt+KStSrZToLrFFvIN0NQp9ItprixCl1csv6GPw0pSPQCRqjwh0kiM+5OBBwhzmveN3iok00hZQ
wDM6wNvqR293VCK8MV0ASL4BAm94GJb1k2NbTHAWE3HZlzRoXvUFFclPvgKs7BjAINU4jG1RyxNx
Vpn6uBdboAJBD0QfxJQn79hokXqtn/BZ5H4e0teeb6n/OvyWOYUn9w2x8QlNU3TfZ88t0opGbWuK
XePUEIp0MuPDaMAePADyoDu1UGGK85Lz+/3RUv1KHZ6BHA44Nuoy+t/CTqR8k42hpcSJEga9yUYz
l1x1Ssc6EFiBFx9SEn6ySqNKR95MVhchb4enM0i7tP62VMmHAXSEHDxAUTzSUQACxpHTyj9679Wq
FFuoPveWSM3550A9FEOlCcgkRf/0PwcFsDA4YVZu2N86Smi4rdrVUBAg4egLVcsmMl1WABKw3+YB
YoX2v8fl/XMsxN/Kc7dpsIlSt4om6P9H4aWYdHEldVYuT/xM1+SU587tOUB7F61L3S6XdX+d48gI
2ERtboABLqQZXF+x3CDNH4n+B5Vz8gJ5hgYnXABZcmtgf7fI97WEVsKoG1P7Y9VUtj88U34xaG8o
qBrNsO9eXZDTOFZolA8mFG790I7ub2JmE1qZI0ygIWGiBqQypH/TKIX/2VvSmCa8VQaZkEiob6Qu
wln0apMATn6x93I3eJtCUqk6P4Yx2iwVjSyNTB1p2Dg3w0IDHndIo5X/rcuR2djK5SfeC/npwfgB
bvzlyUhQ34XPSAt3ati+Mz1Eec4aOk6e75FQjQjoC3akzyIGjsFB3SNA+TlJcthRfSZZzc338HQ7
RAYtC8dySeqt2yMVWHaPpTUyQgxtnRtkjGCKR31lUan3D3oAJzClja4lbHbW3WGdGahks+F5Dhk9
Gtr0S2WUw35+FDWsINrsARRF/2otH7Z8FRM+nrtT0Hpm6hC4vfYDelimRvgF0LjxPg5kRbKZwAcR
hkdBaoiZdsPJ7xCh1uwp7POP7R6QEZXayRKcPBaN9BQRWyGj26zXRL89M1VN+jy+OlOpfkIWgH6V
ZHvkkWqn/XlN80mhf1hY0Xmg+isDZNU9DOGzYciDkDRGiNesAbbj71EZ1AxG6vrRvf4V5kLOnPe6
EwPcRLShC824ZKxwm92hTRHRT4IURMMLdfq4Yvy5xKPOuvGKoZcRXCMIK1LYnaRHiF0rifbvH3Wu
ncpgaTxQsAGTkGSf0we563Hy/VlkTon7xu9W1W1wHPSDE0LZ6r3cOiFQMqPRr1wSh5qDIuf/aaJv
t8753N+Jrt+YbSu9LcDH9eEuAeztDN74y35PAKjxJKEk+EMZJriyHHc6cm3t7jMZ3UdBSGoe3V6S
CCizSn3jp7dj4NBh8Sf7Q9ofLF/jDCXNZe/xO24MlzRnMjhukTUiFL2cEs9jDT+X9wH2f1c87RTR
L3+qBzSctFTi6crUVcEbJxnCSt/O3QqVmY3MiXeXnB2v2GMuiqdCVYQ3yIfa+19sZHi7I8oxaBuV
vea6WcB9oaZVCJlwmJQTVNX39aW2QbIHkGl7yRNYC8R4Mw2lZk0kkkFc6xmC/1INGC1eYF/1D08t
bXMi2uR787FaEEoGm6cd3Aa/1lCx/jKcKkH9gbTcGJ1wl4UcPi46yTHri1nBHa6FeOagTcUmCalE
7/+iC5APY/KK08+7OIISoEAYG8mldnPyyeZTcSZKfwTrBsV/vVNq2pYiy7MovrcGIV9L/FHn8GTR
kGAb8tpkza3PkPW90Eb1mUKDLXpFwYXfnp54v9PPvvgR3o+yNWWlZjq66FQgjd6hwYRIKyoGPaJH
YOGSfDOHS0aWC/fmC8YDE4XsLryTTZkO+FJTsZUFhqxjjccAQidgX+vRx2vrskteEss0tnFB9mG9
nWmBsvYkPu/vxtJz6tL8y+cCaeP02WwOEs8BbT2pMB/kBgn/Z6qKpFVIzSGTNatd45oKgkjDEVyn
r3EYDMTDQ3w1nOkk1WOeZJyDVoC30Ic965abZAivOaCEKmSB1YPj7aHBLUxdyFQ+lWH1ZBCIrnni
LpzbhiudbJq2Hew2ta6rwzxuEn/YYPSRglRWBS2z/GFhsp92zsKsgr9Nip40JHEFmFsFMdHYg36E
bt/EDILuAdqEayqBMxUnTM14d/jOMBxEe1s4WlhsEZLRsdoyJkpw3roz1isO6uKcaJKELOZ3KuCS
WzHr+yefNj94dQj92MsSDxs2wysh20SrJA+gCE7wnx14u8JuXkACzdqoFrfWtV6KyoaHLKT+fuMl
zBKpzOMx/jTG3yM2rOXarYEWxCZRAfugN8X5wCKr/PXhBZS+xzlbI5tfEy6EBRYurs/9rNvL+unO
7Uzg1djXjbZeVXq6drvnavY3XVVi2cETBNvQnohY3ef3ihcNlogNH9x9CQQRnuESN2ApKfJMRF+r
8sV9/ADHweHyf2Y7BOH3jVQq+gD8DKpmob0gtZ0Sz9Pl8/B95T9uz42jyNT98xLg+q9WmNHXPJ7H
gtAX29XZvrX7pSZBBdpn/QUytjCB4HeMWHw1N+UmtJPq/CRoBr3SspkqH89E9aF1DTEserlrpNqU
K1EWspmW5mvXBK5n6n4uM1xLI8ne7uUsibg0hQ5nn1Z9/ldUORVN/qjW5VuRsK0vT94mxXLugLwC
oxfuDJIIGW/bF77y8wVy8sVu+0TR+NJtW9QE4Ijp8ZXYVCu11GX7rKefaeftDN8ybtZvgczqTuPA
a83FgMaYUmJzwmJlG1XucHhd0Pl4egH+21wKyHNGTMeNO8KWqCHIk2i3ocClSb9sx1YlOdP6maB/
gXJmhLfdISoJ/BagdEqIH2AxqmbMcaMrANLvqUU6Zkb42h6ccM7abl/eaa8muoivnI+quaOTj7Lh
gm+lbDfORGYL9RkSsiZe6dUkprRAhYxx7oKr+TotDp/igFMV8Kag599kazIpyYegdLPu/XYddNrX
CGVrSjKpLyeIh2VCEeNACa+YUktHjvaKfRcNqXsBzjL/rRHhMhTXdbY7wRFuvWcjwlwo1HoGrVJn
lbD/qKXSskSNhyL0QgxC4DMjdUvb0wbkarIG/JPqtKCz8JAFb/8uprqpidsIf3jDelIVcQAl9PHi
Qv4yyL+++nxFIAfhAn1/RcB/+v7Py7hvVLVDZbAtP1MIuL4f2lXzLlJiTlm3iwEZkVz6Ce+2W8Zp
YH9JNukp5w5zu0Q26KccOiDileu/a8vlOkKRUEqEUxu/1QA/jt7ap048VFcEjVqMSdvkLve6FK3d
8yz2nA1akM+MvaaCQTtsHCSHKZIgiAspkGO4/Nl/+xIK1SXzKl220POI4VgOJ2JtibEV9t+nz3AX
H+i76vC4GQdTQsPH6wNTtdPbYHD/uLKZwebr7RrA06NG7tMalNhWJPN0L1TwAfmi8NsBcPiuASnR
1tagSZiij55Tb4doKuQYNjjPLZGPH9goONDmcHuU6IFM/h7inrogbxjiuJRC3HhQCorfGFc+jGTV
MVsEL1iexnMAb2a4/o8M1GDui2lRAmAMb2umZhuzL9LFXMI0KaJ1kRiMGqigX6zecL5Y8zk78/vt
QJPBn0NInD5NhAj2aSqfSKoIdmYun3vh/1FVjJOrU3Jp3HnurnFDL1QSnsGQqZSFqEKgIZcoUY2v
ptmfXtbMrArTCHWXQxjO30a0JOGXeofgQB+/uR/D/k/2V4ESsoHLgK7/SrtCaHWBnIYFSDTfcAeT
rBcyRw0h0HzhiZIOz6DpehDp3FVQEdt4TkIpt19GblEFxUdBaLfDVjQ82qws8+pFdxbVCjJjiPD1
ic6F1CHp+COnlnskTt7VuZRsK3h9ng71aYXrWK2r/2eqxwJiD+7J9RNFcg/JinK1sy4uiJHcBBuG
sLlwiS8NXrE7SiGj/N1lYf/rEeoenPNYEIWj5R8J1trhfA3Y5vaDYHtYIBbCtmHCuBA3L3EIinHT
2IFB6Y+tHerdUMUhky5cZ8TDjeCr5Yki9WmalghRH5w686igmaVYjul6h306YHQ9LqA9t6xpqzu4
4BpZ36gX+oX0wxTBTjyx7ig8m6EwWF62JWFJjL3rGfYZzFB1L82Pgx6j4rwOXnHIEFMG6vnCIWLL
cdAdOPFsvIHif9v8hcDF1P2MMaO5qIjyiSN9A2SOImTqmM9txOeb9cDMKZwSI/9YbzluI8VPN/pt
jAjW2x3IdEKnJ7Xeumh0YlBeWnMHNPjQ1/wbM0RISaqVSfi/P3FSfJe4dU9WyeEbPP735i5bhXXR
0YWnQ62IiSZWpX+lh3zJXRo8MLXIBWWq2E5aK4DRcqud26wZSwUN1jj/WX03JU3DB8xvAGOeJRsQ
c70GZfqk1nrwl8TwGIxbiOE5DjYBuNcO917371E03heCfxYY1LQKpGNIz6AK2xwdzg+61nS5Z4Od
EvVxsx3d9RSBcxp7uuV8AWLxazhaCAbJUEIO3UMhUWvLq0GPe5grF/xp0QtTMmuh5wNBu5KPRuo7
XBfj136SBT1UcdburFS4AcPgd37ZXEXygaSTPezH8xzLM7h3HbOM9kmgHaqEtNKGizDA2YAUcArl
Mni6D7i+Lm2qBEgBFuGE3r2MeLqATmBC5YhRcUyf56LBgQl3EhCEYUiSp1FeAIgnZOW1XL5Ug9X9
xwburwP/lV3Atl5MiRPRZyH+vYAC+pi1ehn75sq1nTWaKgtBQviKLPBoHKmlTODKuVcJVbYuJ6NO
dnLBzjsUq+m+rM3gbOxzI66i+hFeMK/JkX27u339bRDbXwkJ3b/yoArAXvFwbDQbHmPObWoZQMRE
s39CAFqQih7pvPi35shpTibslMwuySPpNzxsBN4UhPx4aUMGHxKZHVxbFSheDfAU32114lOuc70u
E/5NkrlbQxRNKiyikcrGKpXF+Ziw2MYyzdlNNBa+cTVzHUB4aCPINqqJciP9hc9yx9/vpEXJqNui
x56FQcTmJqYAuzd79hzffDGQuwiDequNoPlpGE8gq7NyoNBR6h6NrNzwvlGsPkQf14+xN1d4DKIS
vcVWJwaGaVfGyqfO1dIBnyTb0gbT45IUWDe8g+M7FBv7gyPXpZSBNENvNEGwM8lh/9BeucCZR8sw
akg9m79bGsO+oL4HdBipOuwrrQNi7/XKh+VEq9SEEfsnE3K5VUm2z1dgz8IbV+CXZTkipKhmpKqf
04ywXJAAGovDgDFhq0WLf/j/Xoy6xTFVljcUFRKYNk+ww+pm5RbR2irc0BJKhXV8gUyTxWbJWfZO
q5nQuv5ZxaMSVnm4S04IVlRPGVAZlYd3mf2o55KNp0m9+5dZ8dduWmIXs9CUjcwfLZQ7NYUOADHh
jQ/81wIwegrLPUaMx0fTN2zLn49glbF0O65jP3RGQK212LQkLJ5XtF19ouc180XFoL6aNRYWLO1L
WtZm1Ktn8wIAhgUbMR317nLIFnr3FDoPZ2FLk5PoSTYHVS4PtJoA/Gs4z9LSSp2VjsDq830GcE4n
bWWkRAPRK+2m2uosV8VMnzjmrDbN7ZZL+mUSwX5GNmnupM5xOAxOCg/kIXZi7lGZ4GbYe9ZbQ33X
wBp8hWQMdxY16Pg/oSBxpvVT4u9chjL1dfr3SLhFOra2JZ/GupXPaqkkS6FdiYO8MQ9EnIt9QQuH
xT0HjNRoTCzqkLU5v+ijlhwEKbE5gT8KakYE64TzB7P932ojXyTM+O0eAe3vXuTSKb86ArdH0uqY
47spdj2ES2ElvINaiIXMZsmP5/yfUWeJFZ4l83nzLsGFuss34lzHsGyzpOzXzTvDFgRsMtuc3Ril
gUfcv8W1Gj6gTFWFAs6apgMzY1xulOjVyURiGwf+tvQXQiFaAbNJNF3DvAjFMiDMX5G9l5C1iNAu
Ww9nHZHqGMWmKLykjZ54OYB/hxQGwyJ6duRAxgrGH3UAQ4HIFZIV2I/rkDkSMcjW4MR+0djSxZ3o
wpxysV270PdoOmQQRi6TFny//NBDCIj9AqMX2w8mEOSTMIUuIsJELrO5zoNM3NhdHBjp7b4c6IJ7
DV5JN9LW0XoOVoc5D+Tp19BThX9CB/kfaUaW0xFvlTPxiR5XF3l+4Ke2hSfKCDZRoNg4tgiQs9ki
AQg/W0HVoqNLyC4R72mJvdOnDGYXxKuk74cPBCKF26K9ffGUCmsHH1hDs9OQ2B5biMo8o3RlwjXF
HeUdbo8Vb/HCxP06JYMg0JDYTcp7OlvIfHa2aZ1kF7Usxu0n0NgEcMIPMZCxS3icOr8pD+R1HwEQ
tjGXbEqesrm9cGjrqAo+ALk6TRaWV8OFqqMvc/2ptVBYR+gjgNDvoNFB3RHbsPdKWQYrQK8F6QYT
pBS9Iw928kJUU1/1AmIJGzF0VARc35iZEMgR/rQfM4kixzhVgCGQIW8/VOVQ7jET6BzHwDPO6hp/
z9h3kmQdgJD3D50O5jFL2SHrDIR1SaBeCVlCjwDn49nohe1xcYgB3uIfEZP4FrJ71K+76HaXEu8F
Baxs6FAQWovG913YHBmmPmWonPwmRDwtH5A4LuecgE+l7pPYNLjtanWDkmMiHOAKQrwfuE/oMI89
A7lLiIGZEegjHLaVvFeBjgOKzDJxzopx9+0tqTfGbUJKK5mFANTcIFl0QL1x4lJKLIa4F6wCAYjU
1ykfVZrHTGVKlShF3otNJidC44ofC+b/z7TvYsqILG8TsHiFn7w9LC0kdKjCp6eL8bcQWZXAbNQm
//tKuvJhEcOwnHu1oI8jeMgNvLFfSPUZdmjsCJXxA5IGoDak2/ZiNHOzkabTJE01gLmlC8xGf/Ev
XVB/YJqTKWoedeIFRJZIC7OqYNCw6w4S9OWwBwz3EGG9AH1udE1DCXbH9RZYAT0MLpVmPIhPO7c2
HQN8El2k7EXxndrNIO65zLUWWYiLo/XtvMBImvtrP/2dL/qr+nF16707Pf4QWnqpprZM+x5Vk4SF
G4tcjQ6mxOV4czeCJASMlZE1IhXr7bCUh+JC33OgFBM7RvBprmF0eEtz2QfFMQSQaKxTULSqeeWQ
mSbzjrUL0gWsRMfOSXE/RU0oVNTfbo8FuBxmX6DbD846XKSpZ9CT5nF6jgVgIlGmCZs06elyRwfa
lwVAkUzmr4HwAgc0ecmGbK8ZxybGFZiSCNsuMgsjmOmjKaKBwqiaFi+JVjI5L7+B2OQHL9VoWdUQ
LSQ9jdGkdh/BzeyNAK1FmKbUWxnyPrKxCTyhjb/dp/x8eVVVmBILgNKoDCEJ7nDp7Bq+BTOmV9Rr
fYGOzx/aw++wCjd2APN/LuQH+xgwJmMq0wypS1aSVjZE3/E2C7YgXxK9aERfcs9x8LLrWMJ7rOyp
C+l/mlm6FQd3wxSxMx7h7DJfqTMMhh4h3c/xzApJ7X8+1f1dH3iRQvd3a9zENHd3Qwk7LYddLE/J
oGnpwTQJDPwv4ZZQzEyhqyWJfUgXmDlprvyQTFDGrMOdEck8B4U8fjM0AenQewhefoQ8r2MXrkqa
LDJ2Xk0jjmBZVw1sLskLV2dv2LutOIctDHRkeIl6zWqQUrWLLW1HPtDCjb2VRSMBGvfmKt4V6DBg
yzofnKukSeNhskfHFT59tElZPifGkSLqy6zAwMTqOynFtd9AqFe1Up0B182TSKW227fO5G/qu53z
GYrsFipkOPUjY5W4kED9PWrhV1GzYkTv5Jto00p8gpvbes8g9O4sBTAQE+0a1gO7fWT16+1WLg0x
h6VcidyxbviKvtOndr5m+ctIUVr1qufIW4QI58FlV/NEXrKA8mQAGAj1Al/9kjRf3kIssN58ExVJ
ZIxOrIHEAWqKz1Yi41wvXkHemDMQIOKLvF9gJUIzm2wDx2iYftGbKXuNgjZb+oi2MqSoSuppMa2j
fHCViRgLfhAgqFMFXdN38ztY32fKJyQoYup8wo18YfAI1OFAF5tmk7sDZO4gpjpqkXa5Uq8Vy2tr
IaaUFivgnHl2zxsiJZw1MkYlAwdL3fVP49xc76yTLAW4I9bczZ0FguRWQQjbGQvB+zMgj1gfZ4Hh
ynxq5yZcvfc2VDjUR3RMu2EaDnh7VJi6w2bz4yXqgqEQ3QmeiNVbgkYw9GpEqClDQeBS+PJ3j9u6
zOF0tLNfvMy8gtyjUDGVjbFqixu2EQGAUySVp70uY88iTtZfLdTrikTrjzzCH3VbKiLl85iwOADM
sfaw8PwVOlGntXSFv1tSzHWMJCW4rCzus6sRi9iQyD+tOR6TkzeoT5RAmH0Z45X93gXl1X0xKDeB
Vp495YOJIUuaH2PewIlYHLv30s1tEcfO2BTXTB/eLD8hHf+L5Q9ypNR8lywzhENAUbAkU5ri+2fH
BxSuXxOvtgTkTzzsoraboGxWJkjI7tzfR9KzECQ8Ko7q5o85cCS+UZwiEM0QO1MlmjEJew1plvyu
UhehynY/v2gEZPWNF6kRLQnRwFGQJc6CfUywXowdLnZPmXE2MtEG+YnscvG9X9X4b4baJU4WVvGR
DeS8goqggSJGQloPcJRaysPg7/grxi8Vl96K0mjRiLyuiEmgwSJaA7TL+1Swukswj9c6PsITlahF
I8/38DSpz/CffbNnT5RhYHfpEDs+/q080o07xxM6hbrZYhMPMVOjI7xcSBg3nLConqtOJGet4oEj
YVKNJ7whGknnVsnnczhzqZp/CdK5StN9Ae5mq53sToJ2AsqoAyHACSjM7WWohHGNiT52xQUL3OtV
Pn+kbTk8ZQZfcigHXtLv7Sw9Z0PO2bbgLVJ0BNboDJytRq9JFhyb0RQAzFQHWptuvkt/1XrKp4TO
YhQ6UV43pFd/yqJ9DXoyIjP3gZCeAo6cVV0185EIc8RdEIu0r9Rk2b6HjEcOeSgd5nrOAj7i4TzW
8IlVPHslGQlXuy6miRYZ+lscLWj9TAboWTpbweOFAmaKv4B0Cyq/7xc6T4zHPRpd/Q+t1DTQ5Twp
OBiBs8D5ELeWSltfaQQAy5X8HGQ5kPEOTI8NMyu3CB8mM1M02yNvUDbhBXaOIO1fXCmDEwwjs/zV
aLFHvDBBgguI3SvT3zWevOSPL5wR91Z6OnVeyzOPsSSHhQYwHUIEzUt3j94/KTbSUGemNvlY1P4f
bjAj7NxhDmMn35f+wMZUXrhz6OvWFTFzR/Vchk6kwdUJP7Ni/3u0IkjqhnM8ZbtBQMALtLzeLKy8
D+CVU4lFDYLOd9RWEjsP6OuS/iFqFvE1nS5g+PhUD3T0601rTpQQS9l0Y4zDaBhcs2u+f+Fv/Mcc
Sit7rBZyYp5eKHTQIz+I1A+QHHmTkkw5pRiH232oCLe73kDd17Gq2/c8HVX6hH7Hhle0zFOJzOON
r0yqw194jF0jtyqfjrdI/9gN1naDbI0xs1IQnlU5SL8D+tvn8xmQ2SViGHQWR4IsbF3ItNfPDuAU
IxDgcQkG1tEPdb2QW8COO6KFCXgUF0zxkYtL86uZfIjmzdFIiplPfv6yJc5mNcKzafGFLYEmKH0Q
5RDmWQxgFfW4xZx90/d/+za/7flo6DV0IL9ZZvNAjKtKjH6ZI0R6tEr9Ywgtpx68tQzZ/uufkkSb
xQ0l7QH1ApksZ/hXy4ou4IU8ZZB9vPHrJ25emjrWE0KRnv4v5zmw69bQ7pCKiDIMCiyQeQXDYygI
yrndh8Y0r5xj0m8pErrScfRbGHG6lZRM0XSjBOYPl+xCwaH2QhO69JiNUYNZmD4XbYtiQTT+camu
roofmeNLH7s+XZop5DtljfvEoslpDD7pVGOPumlojZ3SdBgi4Ig+hy5QOMu89xQprHAxINmx4bLl
PnwMNG8NApGNBSxzEG3aSBs7oj9q9B7fmUR448WoYHTuj6gTBlX8YncnEsJKBRHkDqvzxSmxOxzo
83z8JQ/THJDKyiEwrpUQfLsjw+3+us/iSxuALcLSO+BXSUwkyxmOAk+OxtOfQWuM0MXf3KHlFahx
yxGBvhIDNg4W8PVQA3MmzLH6CI5MvhoSd5aIrLdbwClxKlpc8eLfLhtITc2Fyzrk4w/cNFPrVgtT
b58Ym8fELhFnbTvaPgGmDDZV9exy4ZUknjdgLsJMqONOaHJPy4mEoLn/lzjGdJrxHJLYv5Vni/4z
6Jvjfs0b1fK8hE5b2Et92vz6/8G+UZQUQJf3RAevbg9mi/REYqBFGY4o9yKDPbi8ZFBBocstKzA5
hEgSbFYY5rJKdUuNm2SX7qW50fnq2mMJ+N6rwcG6TW6Fjz9jDLe4GhbtU+af2zZc2AHoYQMogMXl
OKiB9Gu9Gai4CDoy7L1pbMOyMUHD9LLDxfreP7QbxoTEnUsQFGpChbhqLrzgie6cr0jWqkpEavFX
dMhNKDMiyrU+EBmYvEWhpBBdW9RpeKbv28BHBIAm3aUGO/RS5hoxOk7Mc+ag7q1GrJda+h3TcbTu
9d7gF7Fl4VOkjau0xR+I1er0gEYV9ARiTytpH/ZO2d9U2A8C0GN6YpHBlkSpUajNgwFVyjbXF5FP
XFT/eYCprupc6U8qb2tkJ4LgtJhSYHxhfsgbXqfiTy6m21EOlAcUfqXR+YBitxO2RHp0HfJOC/Kh
yXXOQ2URuj/5cmm3RDYAs1R+u12DtLe4LUNP0sJhsWZX4t1QHFsXtEfONTvdAcTLgVm+1QC+k3yu
54eIOGXUjpJAX7Bk+fsk5Ia3t0N+lteqc6dLEV2b1uVSfte87t+beJKzV/r+l8f3HOsqxj8NBJFP
epm3xgA+QwklGhJmiwCauzHw6nEVMCuAbMvz0cH3caoH7LTS4gsuEO8/OC8O+A0Nk6zujAzEhtKr
B+VorXj+tUTX6DNh/kHxicbWkzadh+cp6hMG2PK2jvPsNkMGys1II94XpP62eFde6gtM8+5D93Nx
mVt53xznJXhxnnIthPOHCTQUJc+inuBq/2top7T2Y5Qam7+3jqfeP0LxwNorjxd26r8WlgN8bUQz
EmNp902i70hEKrp0CCGlxmSJIF83xH2QyOWm94rKp1CZQiPvVqOAFAsSoFebg1WqM42GcaRlfRSq
bFXL01hK3hbaHYD7apoVgkwNJZ3LYkxSOO6iObxtTjfXHdq6OjfKIi1nJzcg6ujMwTN8JgNUTjam
wHJi9O5aHE/74nWcJz/1omRCEySPQTJcM6dixiYaDBv3vf7So8mUu5jviHh3SuRQfXw5gppv8B7r
3gwSmKZcTU1zC7WebMwiiHCfyVbasJRFyELpOs3KUbMfEGnwHtDXk3RNBVBlOaQ3npF5ghF+GS+M
JttKu6ItroJafTJHYy/4qZBrnR1OucFxOEPSLTFwut4Tfxxjfmn2f09q5ebuc2f3BNhpUQHfpobf
a7tX/nI53+3/LqUjaWg90bImAFRFSH/bxcs7C3gUqdco4WZ7+kQK/2II/hwAdUDdeGcbNtlLMoSa
5VbwaKWQc/XifI2ssudsq9bIy/a2SoX6ZCfQITLu3p0O0wuDqmT0D7Fb8OgSJ8l7nhmSHhYcsBZz
nk5kujlpJfXz7BuIgtfzL0yjeBVPAHi9egmhVZhNbJcgroXHi60BfWvjjqwlgtWING/jZmDqSyVe
uS0yvsikHt1hpYyiXdxfYsdhCI/NsUKewD63Kza9rlHq6s55RGCi4FXy9z+0jPQMwY2/3CWdGKPV
ayLvNGkCO0B1eJhJnCLTCu90oJdl0ieJeb+tDnAmYoZMKh1GVRAmGXmu/7j9pqr3K8GCdtXrga1L
EzprxFDnh4FifdHY1NVayGmnqQ/YixA3qVEla1MiLGnNL3Dl8kV1A4xEbnXo3BDEdkKOZgz2hQnv
Uq5dq7MqsTpc3V5f9DL1yHEMoowdPXARj5L0BdV9d7+2zZ3AZERJk4m8AEeG6le1QNeZtWeygPy5
cokbwM/x7dTl24D2qM6oqMwCKvNSrFLI0qCsNy58yZISXT0I3X4nVz4jW/5gihcDJ4ugzoIceRax
4RXfVPoW3WCxq1q9weyRMFbOauq9HWEU4M2iGZUg037B5hvcDuc+eKhNAGgSESFRnhDw85xh1IK/
IpNq52YynYNZ81Zkv/8pnG7zCGAks76CDNnVkInRtmOw4EjmrT3SfK7hv36WXmvDMeGS/D3YNnzO
SjooOBapJ6zLjxluEvJPb4PkIZ2xMoxDtDUvxSfmTnaf8molQyB5Rq5/a71JfoR86gesM7FCGkQb
Nkfwxr4kh/WUyHKb8njXPOyStRPJ9+mtqn7zHdIdC8Bdz43Onn0t532geXAoBsPgMcqahZx5dfVD
CT84BOMqvrDyOIgNS18EWWftTvHiQT7Ela/zZPjgUGg8feAfzYvGJXlPRlUtQUEitLqT6ImBiHFl
L1Y/Td0le9jhBHyWIXzC2UND7RFKCTd73FLZGimxRdN/rhoyR0iBagNhWNlggPAqs2JLIU9/0l7T
TbRuRv6qMEzjC9HzjIcrUnBMiVpyoEsNRCd1+tpFVsSv5imvm++ss5kcnDEtqmiW/IiuNgA2THef
amyJV1zvew33d5jXyjshHBJt4PlbnK+r35y1VJ7op/jTKSRoVhlPAIi69D8IMHHF4sXEIsZLBccf
uV1IEX1208LeCASlaCU2MIiM5phuf9d6BAzo5TBllTXTl80tnLFVImLbJq3LoaMfpPloqtkoLMJt
I2PfNY0wnkU+MA9V717FfP54TZu9Y6ip5BAWXpsOXIU7y3tvzFGRiTQxT2YfFtCUCUiBT6IUbun1
M00bqVHW7MARC1OfwnUsW2coUiaufHWF786V6mJ7CAOsaWkCl3HgNO1RTz6q83KqR8InrpM1Nbed
ICqYdlzwDaFUG+z4t6phZN5VRlj2Wx7ogTjJepUVwl7B0yR7J2lY0aoNlkW+cQPO9HdiAUDbXpF5
/yXPL2fE1HwWCV/bJ72tRlqImQhdXumeBQXgA8ZU/W08M0/FaUwJ2scRRd7Jhok1DmIMl7YRtOD1
X1SzBSyv+D2UJYc1WZxgiokv5n/cZ85R4o4HRjBChzI2docsCgRK/KlRw2EG9Jy9WS+9WoMwT9yX
pbJTLy9wgZ3ZlpYS2Uk5YJIWIQlfrvAaprBAO7Lh+mTAUf7QiQ5zY7W4Q14mbr3oY2ZtSQ2SW3bM
Vc0meUvBRRWQMLodVupTndY8CQXqb/owNuqDKbp+3bfbPkwPpb8sJwqJIhED3lci5gLiwbpbFjj2
FWHCRCl1EN68OmSzY9Rsqp1MrFViH34G/CTtzWL/rhP7MLktetnkvg66FdN0e79hFdxCfpTdK9vx
RuZ6bx6x5LEdA5bbSNZTV6LisIEk6OUToN0XFNHsuQpywksZdV+N7Mbl9F3j9qjb0Yv9Uj9xJf+z
rrZhX1bjYQGaLsJdCD5eGk7zUgkiiH1/4vj3LCuJw46Drs9NIejHk2BE5wHH0eE2mozcdilaxGE7
aoZ6gYq3K7XPJh4kUfKOziKBRIwzmCV85pASIes5AgJmi8m9RIigs/jrSSjLqQLBkT1cnkn0e6tK
9zDpYvaUXtEQe9zUJ62vhmCbR19OZSqCSWS3dLzZ+7gaEPXpsoq2CQFVFgLgli21L8g3YTdgQBb+
N/Dwnw2OIxkkngFULGUEdzyEApaRHiVNMM+Ape1VGCIijoYJmE4rCzT57d9pLVnrK9s+RU5Msx6t
qh8AXKg9HUdkr4OL85TreN+IQcpJe5qKG0fAoImiaV0Avb+h4q8abtGaolrDhYgGpZqgFXahVYEE
0qbw/DsicIAfKXnp7VaAAnxA1/Wv38yJKC7ql7NKD/LfY8/wFQeSRCAaPRPHy0VwHVbdQaoyMFjX
HsrmfBuIIPm8oxeiDSevmICdxN2o3nAofyDmuLpBmTq8zO/QYGFtLSI5cV2zAe6lM37qOu+kZk3O
D3jCtpgHaZpm56kh/SHLrrak3hVPrabMZbva4XFsKSAGUfmyZbdwMI2Ki1TfBopgB2/x226h60as
SllqEEFX72A+vuwJou74PA5VL917pwZYWh8xgVZemJGhe53idsAeGJI/Tqe+peSJqSiRGtbD1HTl
jtKCAmBFB/KN31pbS9vJ3wFVk1pWMlYo3nR/7mV6Yg2SZ0Za6WOmVcKMYex1XyO+8Vu3v0eM2JDp
vRm2FoRnCTbMR6ToHgYcnO7E65hJHJASyDX1kzUWp1Kn1cGN38cLQY2gO2BqHoIpmgjVMv0nkP+v
IS3mNGTCraleMsstFnKSDbNs2YyhS00UpBEBeA8e2DTC7IAmRSrfYn/GSXo122hiRoSa9KZICXkY
1mLz62/aAk/uTV23O39Bf6DWrYuxqnao6Bj0zkqcxHU+zHyLWOF4cLrVvAljnhjesTPbSHDwHhur
soi64MRMzeKj7Ly6hklqGB/BEBgqQcB/BlfanJBAPH9GglXP+xKhGCQ5z5E3bJ4GMGJWRfVDm/xU
3nI86PCxnwOuRw1EySHf3d1CW1TmNN4ZBdBa/8Zol0qXG9AvxBhV+A8y2/oJwYAPsFwUQ1m10eK1
a0oLvm5lLs1LvpbxYgdidlAhJ0x0UxrDO9Fw9g7X68BuVkmGPCmWSRCAFBzpgWdWe+OZ18DGHbF3
gC4QwDxf1xBxayH182VpYTR04dE3qJ0/hciEZWmQm3ZXVSaMgyjHrO2nKt6cbq7no8isjs4R9jaD
z30x+eKTsNBvBxXoRCv/GQ8sg7hwweM9JJSWEtYxqZbSC3uVZgstQW6S+6upioUHRH976j7xZFnN
xIkj24EqDQIyEifYeDLDiHt85/+6yJFNdowYVHE12S+4lnmP/sbvqCs6c+vtvQKpgByg9CLu3Fm1
tw3LSGX9ALkRsLWfLP6EAdQM2PbPoJtqe0JCKf8I8+R8u5DaVOjnxBFuj+XlPU30SNbp43i5LmLd
f6SQF4zdLxit4UDl2XzgmL2Qv4bMTFx6VZvxgEpHtdkOIUtb3ugQFFbSsfZpOY6w8ZkhUhuftMKI
sAgsU0F3q+jxrK+v767FgDGHrRYA+6ezAhjnUESenKQTJLnBbCDXJLEoxjQG9hijD7IFcocpmjRb
8fqafUjgJ2zQgFhSGjrk6YPHv1aRTLE4fQXR1AsszYSXnFNYvLOfiNykN7PX3AcPVo9ndy5pd8HK
2fJLlC0ALzzCWM7hgbQp3anU7wZ+Haf5sInbrc3G7aWBN/Q3jLR7uEiZ7ZEs/0gKfADE7kf4isHa
c6qDZ5vBgWFRLF6GlWLP/9vAY3Co0dxbw0RvLhyT1l/LbViXkpmyslZ/poEz8OpkbhEUc+hG9RKa
aRMVC3LkDOoyFYnL1yafgCZ4b8uG4Xedffaxn3Dff86sldfZi/B4exXyjEpYxAgXGREBnUP2X+Ti
fO2EKzEJWY7lA2nYjyg4rNtM6hcfeng4S9JcfUZD3iuAmZdnq5S4AyfbldRSkLWLa3vyMyCFbJrV
IGdNqOeDG68CleypJgwAsQeVjMVTGkCqaf44O2X1+B50M7mGyvlp3y7iidoF1k6g+ZpuvKgZzqrG
h7z7sdxBR91jWl9Od3PfL0GmVI/S71Id2BYM8myfm5HEdYkvKsTvG0vSDeg2o4asK7NOgHI+5ldq
dTMwSDFw4X+nZABR2LvhPIkfLBpUk/RchqMcfzXlB4cNLLuXpifjKDJkXaW9TxJHb4egQDYl/0KV
+23pRhvHJXShJpEvg7gMAWyONzJC/RzBHwvRI5NLTd0iFrWnA0RQg1jjAVklbY4U6RSCdy34a97b
xro4bU4GEFamUy94dwVc9smkJlPJxplQVlxw5NMkeEZFB3g9oxioP1vMlc4g4pwgmWbWS6wOK5kL
Vf9SNFP2f1YJndI10HV2Ujyk7GknVWciDXDb2o3bFUwTjSUwVChCxbRvoN+iJIVfalSa6ybmAWmW
zBVNaibuIeR6HMBRyZIhFSEewCbgFhfDUfW7/HpeSXOhBSlL9xdK99+3/gNnPleXRgDXIVJR3OYe
Ow9Rs0R7Zq3IhosM4Ng8cbKeUmEt15e3ny5T8Ki7qhnyTEAyVI3q//dj9aRb1qBxvUZRnQuJ2yHl
zSiFlx5cBgcVoo04DmJx/AQjl7kgtGy8hfinvymmSWlwax8AGHUa9zbSsyEp8SsOq/g1R+m+hEy2
DC2mVCLqrzsnQ57OprpzVaJBlNtKLgrjO/9wcfRVFkLsQHqU9JLs7pOLyG32dtuR9hYvZiAcqYZM
Ti9FfV5dsfaMvOwyU2PyFTUBf9eSbk3en39W2K7CDFQkxfG9f3Hb2SxfI6sqyEQje5Yg3tfXoFEK
CkzRHx3fCWSODqeHUtrkmzUA1Feb2s0mE1OS730LcL+kB1MH1hap4xW+xJtr/hDG+GbYsi2iVUtV
P+uDfoHij6zBEVeTNbE0VcPZqYJyxY4XrvQ3R9gWrZnIoo6OsL2O4aN5yWFRH5Z+2zUMEnio7oXI
ZcDATsqroCUS5Y4AEN6WCV44/nS6usE49Itd+X4cu7LZyfs+AHTjSA6wML0XeP8Me5g/sh8xoId9
8heMyarAEH0dmHqUbFht86wrMimMzJkOU+yuthYFzksGkMKexd7eIx/U74/ABpwkkm3sjFYF3Zag
cHBGgp4XP6Gb/hnN1s1G6EjF5zwfAju8LnYhUNJIo2k8PEzWi1GblATpi8IiWAIg3kbsexRBcMis
8JRtWVUOxGdRiTCldJXDK4GDqKWcQyo4gp1XIkCH2pLOVHlEsWREjNTcgbRz4nW82uYVBdOdZ+1B
PDEHB2riEbjl4hjUelEF/mPC/R611tz2xymwsNbgvziOXOnM5jw0Dp4BnZMyHktYwHdAqvjz7DD8
kGPHvwTYwKrhZBWfqVJMBQUqf/rYtUdDM0B5eaIw7S5kxwb6jQ2nhs1/dQ/216tjjXZ6it1no/jt
xjLNTT5201rrUNHjrRp/oj1hDFLXQpyL5FYGbeM/Jk6krmqKKTEzSASnHOmodr26mtIJuqq0FkND
B2WZMX3qzWGCu0PIB/si1yYJHvMUAfZqzuk7KrfRVHXxQuMe5wSBUGz7OaN+t1FJTFEaWFr4GzUK
Rg/kXZ+1rVukkYCn8L0KjvHCE7Fj0k+WmtRTNPI0WQ3mkL8V75d3g4lj13zUfq+L3Bk2UCc5d64j
GKL4qAfPFNqqiaxQQZ74q8QoGvpb0lRF++Z6jIwHLnPq7CJAlx/Qn+tO357kmyNZRRu2LKZRujYw
LGx5STKCEOBBzvVsT83mZNmBOA3/3zZFIUaHslNE3NyaaTw3Y+DUR6aFce6PSaECNtJMDwo6CSAq
7+jxTJ5DMPWxTnDewoe1N5GVTu3U71tcB6FUGPZYEz7kDy8uOBFSBvhkyhTo/VTQb15r5juH6LmY
2eLuhfAim1TTv/3CTaxo//GZXBqkvx57tv79sYHZvMjVoAY/sGSaDlWvWdH3s0TXNBGx9NyQnPmR
WFbptL616YA2kVJa5scly5OCc6hg2jTkul5KarUAsNjtr5F85InpgRPi+sxORwnBKGEtwjZdFL+Z
EGQpSa6YqV0z7RTeIH+zYo78fygfx9a4Mmkfo9oKrJre7p6Vz3s+pydiOWTapE/0eABvGOz1OET8
+vkfmogi9IkHVHeOOMeaDg4utr4YDgFU1WNN/yEmR1wUn8sC+HONMleKrU7rTJftekniB6ZMuSTQ
+QfkEnI4e1nhF4O7/lAmr5ikXyyzYorwrlLLluBlP7/PzdRWjNG+Olxre/mHplsDDPieyLnNfq6S
LsT1iLxOv8zadgBcpF+BR6sFDuB3/Mgi7AKhVxpiqQyRPWDzdT6R7TuGihKD48U6Ez91twV9+bNj
HmWnLcIi8V8u09Loqgyvl4jJJcQPWa32Od7zhcVx33zDspU6SwS3f7/F8WFD2SNqHhEqy5m+dFDv
AB0WV1tAm8+2HrPryk5QBV+YVcLb3F+HhBdHbxsV50H6R9SSdgo/hA/f9tDLANyUWoFAHj4xTVfL
SKvZqBoxiXj+y/JvICH864pCt1SXgb2jn+7UWU74vCuXzIBvatxPb3sP8XlSY+LgI+jB6MhPVeIR
rOAFkDeAxe7NcCoUw+sp6Im0MkPHGWu3fBsIdxpPDUSRtNYVEsfoLK08Xf9pUKs5djGiUeyzZHAa
OcAjeKWNJHa5f0Kh5ElhwbkcQ8JlENzERxhsxK4COOF+sZ+DQRnCYkYNdL+HQZwMdloX80UmZ5gV
uKfvT8e/6zG3jiFtxzzqN2c1T/ChQu+UOx3opxcZucfVAnhdoL/esq2corHQkt5b6JML44dXVmdW
0LWM5XCy9QAgLtHfFrmE/Y7JbwG9SfnJPJszDiX6w0o8hqmKud/taX862z2wepZLggmcEiKASYsG
ENQLkkhhsvf1L2WziRsCtqumGvRrb2eWsZ8IWQeYBZjT9TsW8L3etEU26thFzEeF2nFSvItqwawU
KTFjYcm9LcpVk6Vf72gVotoN5cBFniZSa8xLpttYPfAAAh/bFzipjteRuoy+8ks+TeBx/aMUn0ol
KCwcz9uu/90CFnIFM4tWRsbiUEQ4bfCy4/P5QnfyOJYsI9unIpgqPe8GLPmvhKRDYLDU5nCmHxDX
utfGg626HMtH+kDLfm4aGnJjMyA5YnEJNY2nh1szWP3oaxnl9r/0Kx6xWVHMQcS5JGmaXEncNByw
zI1GpJVkgMGrFQXcshzWccc+NPD6K5xdtpRt1bgRBBxIR2LKDT5+RZU/sBkp7A6yrsk+u3CoTmBm
0TJI2QY2xBRxlaT2dx6XWfV3k0zQUYy4eUwP/0+rh5UgxBzsLnimD/7IoSwXdTbg24gBlejIPlwF
b/z+fQWg8AuSXg6s6NdyXVJaajITxrHGBU46N0TfzNShRLGQ5E/Nbg9saA0lbvezF6+4jXyyy3Z/
4rv0kl5ZmFzR2aFIu3JPeyMWCVmC4KkMFFim7/3fp20WF1zqXIN0hXuP5hlM2bD2d9GcVzixtSVm
YLRpaBupa/ppSDEF1a/sMWxYQiWcO6XZF28LNz1B+FktL7jI1/XmD+jKkfsZRuxMD1s6P3YgfBMU
XaAAA8qG5isAdkrIbM9uml+AX7R1GwgP7FkrIw4KN5/u+7UueS1/rBPKdFPHZgK48FNFQitBAx+1
jl3y9lDMWowGjhLEAmwAlTw2IoK6rRZ2uFUvGK++7UvmW3At2ft0aqjC5AtJmo0mdmmG//Q33RKn
2Mi6n8NUTftflXfFNfeFTVjjLbjQnhKgOBXnQOA3B8OHloRcf1Kcw1uZkbdtzh4lQm+gUKaIfD4+
ARXFyWm00QjfpityMnGIZXHaNroNmcbbmzmLofyugU4kHO5LgfCWuxkNR7mX4hpgukU8luWWkbnE
VGUk/fnYBhfrGzPooF6AQ7eCpxu/5Yib+D5RQL8Zsihz3Wgpl1MaWZ31PwJnFUhQlgQahIQ5GP5w
F6JqQuRKmaUf8JCsZA5eu0Od3bZpOK7h5jqG4h+VnmFh9/8ABaLHgsuLNC5jcJp1FbLFkEAxx7/0
2l0CiBKMHM03PPkBfgU1t/HDJzK53heJ1BbgCdWlHFiv2OxZYnaXtET4BX2Os1WVGM/hEaaXptEW
6/jA5sJvHKow1HApJSOO0bp1eoTF4KV4Zf40oVaZ6TKCVbk7v8FZ54Jm0jaFN0lnR6DTLjmG6/CS
/9tR/BNi3UdX2yWbnBmrzglBeFQoQGd5vQyVqoy4tLoWNuYd4+b4XXO8UayLSbszXNpBEnPda5I2
t/aAqgnOA7IzGbZF3aKwiCPZqtvwjqWtJQurqtZ6nwgcQoaIel4VLEgng/83qcdBmLkhaV6zzG1E
9LRapNJtGLfWGOn+yoyjuXIaYYlVYZIJ8aoBkkRTTlDkXofSumCuTNV5LBofjLwxjjS9gPIqzhvx
KhGM+MAcZMnU5ULGXdFHmxpBpoj7AkiBZdEwl1A0b/VvQcHwG/bVbnxOscLuPPrPzMtbli2IMmMf
agRxZ5LD38SrFdWcAcWzVuW3G+lcoYewY1XMkQf3gJL/ujFvr9Dimj201NB+1PY59K0JR3O8YtOZ
CFcnyE85J8RUl94bvMXFjLiuO0a5EbT/wRM7tL97ObH10gIGr0/hXUYTAPIqnZyaG7AD8Uw68Nw9
dEK5UHOt6m4dm/EwrZ7Ho88cZ4iJB6+J+nuyZL79LtRNkciNkt7cQdoru+JqukkrITci8IGKWwWC
WBUZehKuCd7lqEMskHrTC4ruPxejcwy9p9ZLWCvlMuwE9cNVSg5+hkQ+dmVNeeOOw2FaEs92yaX5
0kzX4Mr7bssWz7COFgAUeLogCPYr2Qx0ijpjcyJLl86/liCgki4YSKZ8BV3hZENuj/tGZc1+d/6y
b3+3dqDv/RfJ97m3G0BrgCHwAtU2VLUnQN2y/2qPHYgLL+hjgLdRE0TV2dJ4FL9Efu5lh92m+Stx
VaeUiR/fcnJajYjtDSTVhY+IQc+aMWFHw7jp4BCtdWZj4jwZE7a9tXVBrnxBi2tpIxdZKs0X3j4z
M7bvgcsE8dvBxmT02JLOPcjsZ/QKTiRCABGSZeUmxgf4CmElN8wnKooOGfNH5kwy8RqPzb35BABq
vZ7NhyPiHvIFlo2+fTHYNXcpOSeFeUTNRHK7FOD6T1zkqL88Y7rMXBdVU6P5AJUHR9ZspJqQHXx1
DFt/1LwYt0aYpqOlqSIqJDc7Q4psSKwdY2H0XDqHGyFhoIJ4G3uKec3lTgdtbUzlCRqj67ENinvY
TYb+BgIYK8NYVtkTCIaSJH+Vvm1U92CjpPQjEJtWSHHT3UUC3d9oIQbIIHHXWzR52GRevb4MjXpz
xSOmjq1MuX7iS+TOs1bZ4rLgNt8t0EQq5ezQwfd6TrHBOCGlLnWGXkRUpzmgALhD9BeLB3qGXzgc
fuEljNqBhfJmPUqhnWXf2/GNkE5kOKtVR6BWpOeNSV5moXPJd/GRRbS91CHFwLH1Cxe81uZJzGWb
0lmAWXhe6fLFHbx05szyOlDgBdor4/Drq6u3D6k7pAJbWUARqNZpJZPSg/fi/HI1ePTqLUwYWgzb
ScJgxgK3g/Xq+FNWzYr4zzw4lyj5vBZs2onwEhSY8WN2buomKCYkx2Cn9tBZ4RTk1I+jxrR88Vg5
gasugEkjXoKyMs7gfjCgHSy8FLz8xdJYU0YR38MkU85K0PaE6rJE9mDkaq8EC+fFceiHpnJuTY/y
JgJoePlrJh5Nq3eg8mReU/sqM1Sc8hr+SEIg7+4yMVnzOWxu4IoFYMg725UUngEDjQOflb0pHnfK
icxxVTQYV3/Hop/WWPCJuh546/lJwoJ1ekjpceI0wbmFuRR5OL9DozQNW2g6lJ8PnJniNYAyCj+M
LfOySHNbD+svU47KIFm0Vx5+NndkzYCLjJvOC8QDY3bMLDwffvcXR0EkOQL9im1IcQqUoWo4wznc
fnWuiYXAmUJWAB+15q2TZXHMj1MSYHzZro0l4WmfqOF4ZVFPNgJizuAmJaZyeMG+EW0LXlrq8LDs
rc+HTcJxrUdSMRP00BdKHPNAXkoxQwnLFpxCOMvN1A4KjmMKzKIE8342HUZ3krZluZa00xAqbibr
XfgOBxx76Pr0cHyinpsuKylc44hQADXfA9VL2Jv2GxiGnrFLofMs1tfJt3+dwvYEZJ/CKQCpftut
+nRe1C2j0mkXgoVFP+/HZ/tp+JaFiEIdBe9U3JmDAG3grxx3AJEuE9ubxChI6v2xgWX6Fcg6t84H
pcK5K5U6671bJgEZMXKXzcnL3s92hwNCPYhSW0ZuQ6DOmFagBdudzQB0LrisstRB0L9S0FfI2WCT
f9vxTxOuBjw2aTz8OXZhd96+Lq6x8PEnBrozorDLFzdVNFbd0ZzKeI/Pj7i7Ie8Atb3vGzRqTgB+
3yDdiY0LrfOHAm0B/Q2obEns0w3/d6BQNMoVR1Jshw0XY4z2yDGPxzRhv3i4uyC7ASwrfUzh+7bR
SIkWMrA4PoGn68GN/pH7/hnjC01MTDSigHkaOJFTK7ygL7INd+dvdui6zssyGFJCPxrUM90r99mP
jetbZfWcH6l5US6i1Ow/Moijf9V+S776CjnSkaWGTOJC3Keq5lqexDF5VnhoaY1mba05kHaP+NcW
MjlDr2SHzWGJtLE+p545WVZua8Y/r/ghEPUA4KAvLgq54lDmLY1Op7NPJ5e+dAm5mNPt7JacgTzC
YX/WMLSy8ziyYPjcwQSCCqsu+vi/s/y4C1wc0DywNNYFxa4AoWNxX2KifzFSMmbfKTUjALEcJHm5
dsAnjbFvjmUa0czxbjBRGHv1uWfE8FTftAIsXZgYy7zGnhz2PTX8yymVi5x+A3P9OWYfTzg4KOsB
pk2Vr080ZqwJxmy6wjx5g4DO0sfgH4n+8g+S7yqBqtv/J1XvGKLXlsNcK/mEhvTxyW9o4I+A6loZ
CNAjgajzgLZflSRxLdHSdr4HX1xhefpi1dV8d5eF/M2PAH/VZMFBblZ0u0zOwUi0NSwCJIYxgRpt
eARyAWmC6ACus+xT2YP72oex81fCI8YlwR8JNGP6OJ+bvjBw08z/kf8khlpQpC+dOBxDrgbEG5/z
aUhGoY5aweWsZzC5hc2De55wmROPwnl/nkBBZHEbFEih0qcIR7M3yWSOPNXOymdyQ6glWxwfrd17
OmGGR4lp5mXmYkwrw4Yzg7ChfasHNWsYp/feee1D3gK86qcgCCNx6LnmHWKLZLRh5Cr/BFVdFfIp
zrQo7fC9R8vv8WlXJS4D66Xeed/DS4IWkzHm9pwiQXEOWXQDGKUuFlX3MAiRj7RhooMY+F3YEtWj
iRxC8r71J+Vy9d9eXL3C9NFPM75HdDrzwrCKCzoEt/Qq6eiBq1SKcY3XkMekzwbyhaGuv+W7ehJQ
czBQ9Khl1XZiPLgURFq78ghnmpWHGHhhT/g/mYFQhapcOWEmLD6kB6zGwJvifGt5jpD/G1BbATBD
fo+fTTgrcwHTtwdlHIi0yC37erEW0yuPIZyiaCTeZK202rAZ2zGDbHgL8bFUTFtYCAaAZEInYtKc
bemudEFpswsCyGBNrGZD2vVHJ3OgS3Yx4fZ5u118Lvy1UXGoV4X3kYRjIjAGsJjqu5zgsihjLCSh
LrQcNQCHEQaVDpHY8115fpawUsHub3D0swbM0T5mvulIr8C5qn1DrwWvGS6wgGWLrR/Yk1Ac0z5h
t7xyH8tuPnCCSyqoExI6V+iNpFgOhEzrzW71677Y1isb+lgLDObnVnWmYdwlNKK+dGuT/eqVlN8b
bNjMnvzrnBK7m+R1lrOMSqBjNCVt6MN3vBfwR+8E9+hzsGVMN1ia5tyidMz7wBB5YlP/79upAzpy
l5JhPOfMxsTmg2O2voKrapCJTi0+G0FfMHNR6GTEwK+TbND4731QNEaYDS3TBHd0sEi23rXeRI/m
IeH2bPt22Z7cA2lkDt/sgELX4zjUk4CT8odIi5AqhQi0GUCd+NXAHeMSY4kS/AcRQqPD2HsoPjKS
yDRmLRNSNEnE/cpZM0IZh2EqV3cSGrbWEnkmtgxJIrbBQj74Lz0W8WgIRSAFTqysckWLWwm/RWtV
CIWIZ0nsPRyMUIl4ZLxyNhyjDq7QeZ9FS8+L8ADFblA8J17jL0REfS2hXn6WVVZVsFrCDKSsQKX1
Q5FmoT70X9aP8v6rsAEXUbhsVhmfJoNrxuH/oRdrsNYm2xv/aIz5iBXvjtqNvaALe4mksdcH0e3i
tKY6Jg4kavYD6NEFpj/hEFqHBay7pKLp+XwFSjN6q5936fCEyGhYkLHcJfY+W9TrR1FeQe5NSPo+
vx60VjKHEx955n8fbSeENV4X4jx3WxX3qVpee1yRgDyZ0Z+f2p+DjbkDW+S0sECcoVYw3y1kryCR
0zlAT08KUlQrV3zVvxC8pgh50ah7nrJY1cHUYyCf4wqDagDrUYQps8EQwBImDuvO+Fp+L5OsR8/K
HVGuixHc25z+ZDFQcl8zttBOttul5zuxXY0QfO/RTQIRBQyU4oo5zWgsGQ6THWu+1s4QHVK4ohbK
p+jNNwNkQ0fdgdLHm9Y7xdL+auRP06bpaTioyWz5URnkw5drOUikr6P9cBYrW/enwml53wpVvSXx
612BiwkojxMfdM41pOrUOUdHT9PfsP8JJPA1LBSSps+5bPVPpfETZf4grftTloCxhn4n7xguF3+g
3WVuqgwhMW5JPhhoFJmnWtRbGbQcpcpcumtVuw7+f3FLd77MPAUrRiJaSNo7PmvK5a0DmRkxF/RM
JdkhPMFi/F7+TsoCUANHBaQWlAbX3DFocrZ2LfVxNH2iUwXr1dgdwBNixocV/WDHx3R0cyqbEqlV
XgjMGoHDIRB/p/iyEKkGYd2PtjQNGZS+G/iaqUUfTWfP2FMXQpul5l7Zh/39lyI4PYb+kwkqD+LF
HP3HsHnmbtgAFJ/eaZ6wqfh0zIfoKg/Y5JeLMQ2I2GNFWMm/IHvQdeO7EFI33VY6teK+EEeyiqDo
mutVfpGZZOoHdAXGbqUIemiMEvY5g/05XSWmN4Bx1gIfMcWVsurdUejaPv+G/QsiNe81ilE4W9Bi
xdivBKbbVzecuDWHlVjzIiZ6bFmVya/PF4cnsSm8Qb50IVgmu6QacKwVV9s6SB+rtShjCqhbsl36
lPdDFgtlUgAe+UqJhkTK3sVaDisqRVu3BDKhD7vjEyyaPiU39OHRT4bWL9a3jDxK1v3Hym1k2YEq
ZcAVrd90tawdp9D0HxSkLZGPIqzPjYW9feCrC66lAcFiGuTe976l6MoR1tdJBzcgplijMkaqtMnY
7EzWarZQGuqDiSODimHWKi6+diw6NoSaSKFlTQ9TknEUbdmNBuKYrJX3JFrFTXmD8vvi3uJIS/Ni
lOJy2WQ7b+ZirztRXPlB02gHkBPlmVOk3C5jio9eYSfExHllB7IkeMyjeZs9k5jKxejkhF+jqKFj
lh4nsgI9ecdkEcnk9AaOql2Bt6QtOs4He7aEkd7rDzNEi/s/PKLwX/bmeVLn6LB5ysEJzRp4CXn3
8Gk5GQq9wSSMej3bzWrf0MIvYHNfHD5NPlm9f8/i8PbODkJwnoYuNYOSma3aaq6UzTbtfIdG6Lo5
XAA5pCXK4gUoMpWQ6c+Xu6MyJtjs0pkmq1X9cL30/EqNUl2UGX1oV6JyQ1tuoAZgUcEerTGXKSwv
FVm6GcB3MVgd8z0PUxAJN8NC1VgYSAZKAfFuJF6AR7k23Dlo1yBsHqN5NlViDWQ21yuzeGA835dV
b0V3g0hIi3hOYFFmL9ElV5GCEt77s4afIr7MKGkQaK/4zcsbpH64PvuOH2K8dqBq9xSvQbDFNxwa
qOvMwLkWjyUFuf38MkyQg3JRyml6pJsh5Nk4NMTJ/Jl0OGwiiizPsBmVdMHP1H17cDCXrDB9202h
cWbsrjilRNP0u3yPhRxJImgMM7b8QiyCqkbVKL3ppl1nKLQRTxT1UyIkqTwKvAOBTj9zFwiqleBO
/sh8iQ4NRtZusMX/yeWZenHjkUYXNYU4kn7dIKkcLL+kOzztA1JaduOpOQZvoPZ4Te2gTtz6FhV/
ANqIK5sj4FKm9pJNmKabADLHTzf+lfoNzU/49vnf0ldwheQbBWctsT11WlqUQPknMgxAVOq+GM2H
E8RRPB0Xkz/AkhkFcZkU/FRUdBue1neblxWQzMDamXg9IjUEKR/MSVbeTkQYyp2hewRHZQuV5Rl/
L/WMleLkm1XBazTyVSUsVlQye0gsmLJVXqeM31bHLlZdMPXFUTX4fPXWJVoHqHEnOZzstjSaMjYx
64WckiE5DzSXCfbI6pNlkj/y5YT6PrbwVxBcAq/Q/pnvmovW+HZ0YURMMIsrHzHELe/c9AxHV0Ef
/KyYVXVT6baWDNaWCUQW82VzpS2ZHTgod3iRc0AvSgtwTNar/t2wxgFxnK2DLHUots2Ov73JOGPw
+d5kOv0WRufpy1A0A1yRUOaDQSMKbfMDmmyswyneH/5UypF/Qi9RysVoJ+KVp3l6STqSNfrJhEYo
YlYc5d2Eq9Iag9J9Xo0x8YkDewt+UeWImwz0G0V+ZsJiwjhyZmP5zxBpp68qANPN6izVhPM5n+7Z
qdRJQhg1j5B08iov58wKt0P9qBdeSZmqVq/cjzwO+W67jI9rzZBVD8ucvPuyVZG4s7Aoy+yoEpWc
IvW8Qv047Lz7ksB3ZsIWpztoGWEuDHz5OoRGlY7Xt8NiuV+41hCzRxw66ACT8WM7rlnmUuFxX/3k
xlxVSyYQNFUuuHPrmGKiw99TInwGOYjrO+t7d9RE9SWNs+ZhduC1/xMnb+LGB0Nz2y1is7cj4Bgw
Crg3gYK0FygYptq5PM8Q1ckE48PUBPXoTr91l2HNLcHh929bXMOO9I8OOMVun3/87xYdxXux3yzr
s19Bj4pM3NwBmSL2KHXVPRGY4zuj5Nq7YyyFlbGVx5+vrUOoA2CzFuMBY/UKZpmFOzsdfL4EYOol
jldmJIfVIrUFoUMP1tZkvfBBWGS4rJsA3VfrDN3FHsBiLQEl16eoEZdjyqNRlYB8TAj2zblZn2Ox
WXS6XQGgCHCEWij/ZtzhIG3V8goNH0GHhXWRSSXIab02Y0sP9/p+sa+CfDHvCuaooBWoDZRq0qJJ
KVedjT/OCYsQB+nP6ihoedTZDHFeA25T/e7o+E0gOOXMxhQvx+ZWUC2uqbsTUc9x9v9MgtEjAwA5
9mUT5K1fur/PUx3FYPfhrKhlk8kIjbjGGLuIxJN4rIXl2iZqLbYIShI7A5lkKTWgQJgZPOUxeKQI
g48P+qYSgcbFKJdydo19q3tCq0rGlHxnNqdSorU1AfX0gmuRDMMU/43I9V/lxlasZ1SkWRLahsIA
MCLAjFC/5Iml4XKdms3+hYd5yDDuZ6avN5T/DPU8fpAPkbDTFnijYV3tTAxgMrMZ8KnDNn73Go6N
wJT7B1eC9TMl/pzITTaKQoM78f5tHSKUyLIZNhHkR9GUfRemzGIGGbrHQDAT/EKoY6GQ5kbt7VPw
2dyZL9W2JkKuBN3HDFEbwB7fVsTcCzc6pCm9kJeVoNp9yI2h6yto7/xrtNGqRi3Z79EzjNzkHvjU
lAK2vYRPrcaPS7MBzzup4HRdMaQRt31X8d9oYVWJ0Q2FA232OibbjimspfwxsLhajZnbwO2lNxID
H5XLMCeMV6EYc7JgvLfzV2TGPv+1XLNyuykHc4ZgOfLmP8p2QQgN4rzQoVkMRsGiU6biheng9ytz
+V844FDe6IT8E6h/b2/OTyM1RZ7LGIP8bcvvj7YRqkI8E5C4m2c+8kOuPiSBHiGwdzgWBbw4wMtH
fSIkESvxwv14xXulpWbJJR+l0GGYpnGQiBZ1mi0t2MUePcIlkxt0881isWsEsZ66OnJdpo1US5z+
92POStXVpRQSVH8QWmo1jiRcgXM0A7z2WUquksMo2r52ml/yVCjzU1+x8q6JIIhIJdAhoyJU4D0+
swXm2i9cN89XbnjFC3lQ4uBNRj8Ik2X7LMnpsQImGHQx4yRaWVNKtguqKl3dalPqyX+4G+DD7GCf
grZILQqhhABWhNxADVOmcZUEQdiNR/l3ZxNCEwJV+Bu61IUrhIXGZdB8ghSmw6aI0sQPOMSEfAkD
OgrfbeP9xoCKL+ukfL1ic8xWxmgg7ammFkugeur35cOxgmDuW+DNIgYKBXYPS9uEHEkYjhO/GxoP
wMjU0Apfcb4pcYsP0d0OaaFmUkv3n8auLOxKeX7J5OnKUA9SKAHSQx7huxlYMxdqxthaEJWDao5g
DbttCI1nbqLxwNeKueYDZu8H43l2rBTtkMNrGekcUucSTZrkLuOlNnVe6WTnbS5H9XJKV+NCWDe2
AlMYuzqJz9bG3ohZt0sYJD2JgZTmP5WuskvCQpTcgnemRTnOYDeZmHaRdrkgJ6SnZ4MHkaw6Xnms
RsFzGsZQazp0TS367X+EEBFU5W3dBdE0InP0ND6P2iu45cUrbaqoklzlTtmkx4RjCTR4fFxN98bC
l2YMBQYM4nnwazc+wUiaBEM+52+beY0u9diRkN7sRRnYHaP0xczBSbztzkLKREDhzKVY+0kF2E2D
+kUynHbYvunckgOmBqRcZMKMNZUMfXWkf5vVkn7BSQqno36U3GkIDjnvwq/U+l56Xl/kItcEUmaX
QxAkLKUMp0MKUUN2SiQvsWPZ01L8YvKwF6budlT6ctsLz7JY7bsEzxFvkh35xsCsglRVt73L0tTG
8SMwxutK/0Grex9nFIZmFu408TZL76nD/Y6Z/C+EFOb61MQwsaMhd7NRzoaf6ZLUuEi1XTjHvIVS
as+wbtpPx0cTDTm/oy6mFvDTsLAqHnD0jyqyX87a7oCA3w0T3WZhAogkY0ttmpkKzk75CYm9yFgs
TjLSLO7VUYDo3csTvssgFZ3kHQRtn+J6T2DUDS8rq1PRc2y4Oclfi9kaLD9zPTV/EOuZOWZSMiHe
wdU6DzCTVLwfj3+OhkAwnZFOZLiVXZowwAnHSe1CT5alB0qY3sP5L11afDMB9mqBcaumFxH6W8On
lPRL9LI14VmdxL5eLiH6nEMb7vnjXeB3IW8HereK5YP0DTX8GGcYQIRgLKelFay1qi1zCXnZcwgS
3zS3MV3WRowhMoQGthh/PWzZbg78/SpowCCXJf6ddBJKyNY2hDuWIaZUfBQ36gTYNuMNBiqnLqxP
E4hg9rGOcD6uSlwPgFH0W11AOjMqH7m/w2ai9hLD2Jg+nBT+BaSMuW0zM2NLwSxs8zAHm/3q4bND
xmURv2bVCLd5zJoACCtSqzRP3xh7ow2WCMKO5dYRMVCaWWg+U5H/C85JI2HPzLJrPy3LbdVUqY0Q
yt68leKmC0K8BQvwIcSY+R8lguw0X/zGPW0asEFW9RCp1DN55nMS9TI28r7FvH4yiYA0ruUZbB8b
KSfAuRJiQL5vH74Sz6MnI8dXJK1sUSdvzfvW6MsrzQFWDXuIGGmq05jcdITvhtc3EjE/XkD41m3r
1jSuGCwBdKk27hOzhnzWGjo3XnW8MfPRUj0eimOhxbjvfoWHtSupFdLpU5Kbz0eB+t0AW3BoJAxc
PveILrjvq+2JV0Wt9bLasIGxPZHu0DCLDz039kqhGOxHdS+8vYeyodRavlOTnNxP744yZfg9NHlT
yXDE86lu5qJZDcbaNh3b2v1z+jXbK5Pum39qtiFdFlXqtPU/QPvDiXZ4khO8z0aQFfKOQiv3ujgZ
fqTHAk8QSaFkypkiBaNQsnQskZFR/PgGVy8vmR12cdiBQsJA+PRWGi/uI74QADHc4sEKRgGMWum5
ZnkC8N49dWxtW137Yu4TflX/2RB+TmHR1Uoytc7L7981hR0bxdAly3MsapTua9Z/afLDz3VAuBnf
Qd5fv7nBmDpKIHjFe+pC0JELOu4LUAuh3UMFwdxOj4HqZDvHhO9hkNs4IeZM2fOyIAIQRlyaYPZH
cDfcfl2lePU3mMJfdfPRBYfw/qpJP3K3jwdnI0VUS8h3zAopQ7Jzd5dbsDvN0xPgzellGuu3I+JY
BIQIieHBhx+j8DKP6UTXWxofOxOreLkUSUx1kWcIU5iLuSiwyUKAoygZ/5S9s4OJPaO6WnI354uM
hIwkW40PMG8Cd1mOmvRiuMpdg7GZkADrJY0rjdIHEK+GKUbyQ+y9Ibvl+1B1DMW4fEHdYcvvsT/D
7sf1SqrVKzJTomyFp3n0SmvZP7FssZLRJaiira8fYqLrSD+uPYbjq0QcGGsheLYLTXSV4aZAuVh+
/Wwxw2ANJ7Tgb4ejwUXQtp1zYIjCc84nYs/urScCArvBDqodaYg/RtQvJ1JkUvQgKT9bcrw+rpBO
3alj/VN3BEweTnWbce6YvU+qVKA8zzh4gLm2DpuE91HYp4RLaqC22220Fn+hMYomrFWYX0JhEa3t
R6hCfkowDZvJqIoXEL4EDmp439IgJuLIgWsTKsY54EXv+BcdpK2L+B8BCSUBYeKoGnz/c46yH+gt
6koPyeJbJo5jOydrisNjsy34NsM7ag4aj0x/zY4luW7Uc+ZGff+fVEMWMp/3lUkh331ZvreHGDoS
EHvLuCuJM1H84cWwsrgec0kfaMtNVUC9I7i+wQoK/oxkUoJUGZ2fTCL8r15cdLVQq7V+P5a/UyLx
HRfM3EnoaUE/hIsf9wPxb62UGJmTPfDBSLgxkyLiBzjz9KUG42whjd+gG5DDvQUiiJnbO5iJM6XI
5VRjb8YWFrE4gjmC/r1ca1nxeEvIqKFLNINrRfjvF+lQbirIxyJMPM8EGzXJAsK8NpllWuYmw+5T
B82vX9+8Yr6jcSAp2s1uKPfRTxuj1dCnmwTrxc5hbQMtPZaHuCy2rZo8s2Y6R0nL4y97/53nI345
cxoS63uW42hB7ToBegCxhELzVOTPM4vI/g2ET8yWgLYvrPj2LYH/cOuEtmptRyw42/Bzei785M7c
ZdUJLOz7/l8e1A9U+NiY4IXiGdxb6MLPfInXn3K8AKOqr32EH2fIYfOcUvN1N/IXEqHkqrUFgPJJ
SuUPCYsKKi1uN5bgoEDiORQw02grB/QGlux15H3Iv3WynLKJZLQYrRTF58xLgAAeALqH6WkwW279
mBT9Y4GYDIqIFg5D4h9lsBK4lNFd3sdxDhMX63nEdM7m+j/3H57Zb+IiG0Mpb1Bcg+Ms8w5dsWKv
gTefFy6KCibhVOWj5PawRQqhcvMvxBfvVn4TjCixkMs9OkQidtTEERSvNl4rsX6yt/+6hD1jSp50
Dgeo+z88FiQheF238DwmB+rf3zl4cuvCVZi4a7kMqZ9IJdpo7BFbhcmtCE6aAC76cMHCfLQ+2R9N
tbjj0VdwOCzCjWYhAFumf/2+8j7ulfoyuniz2qXJT4Tnwdv83dbwUkdCHhjAdbpTC06Akfd6PeSU
FGRsD/W+KKEwvekBs46dclXds/HuJa+Pabvhg1oAqXspWzwfXSeDUfiaRauU69RpV/oNgmXRZdJy
ayWchKSYE1E4ntcIubx4BO3kRSm9Qdq8gye7aMRshBFCJEj0n5+Fxww6MHjkUkQxyxhmi5ivoc5R
zN8e8pbw5u8xThBGGHcxWp33iNwn5nP9dtuo0Ku7KyeqJDe+84Riikc9m5NjIGPmX3FEPYNHTzMN
n+mBzf+9zh94sJggDe6wjNkug51cwulhPNNzQwldGi2KHRuxPwBUEqaJP3QJH1l4czFEQ5sjdGDp
lfhi9EN7miG6mBEk0G2bWz9hscNmV8uZk24Bf1SYB0goZIWRDUsKtvQ1cWASodPmetKEOugUfWZc
ar1t1s7X0FyYIBthGnB+eVpVE4Djsd3AIXTBSJhqfr6//L5ESCW1Vo5YoS0Y+l0TUoCj+pT9KE9C
2L9n6tMaqIMYOMzNyQhzkKClxBgjyj1yawFlWzcyxXGFupXZOzXtSMX7gtEbNNR/9qxM6+bxNmKQ
ugf8DvRkVYfWlnFTsXth2lO/zuCFq8R0EyQjrVbHeTzAMZ1Wf+DjfwIlU6FED7UQeI4fkrkT+XDz
Y1FRlCzrIBP3oD1FoDkUuxbVfNDnbHkAtyG7Ew9z1SMe8uovKKQ56B0GYSTEMGazxEcZuUpbSu69
F9hpQX3I4Vgdrkmee7PcrU77mMJC1qomwqkNewUxdbxKwRzan5EejcDg3oeUxstm++8sXFpkdu0F
f/5hTHcn0kzsz4euBh3NzRrcsor1svD5B1rO38ql0L0G4rmWZgJ9lmfZbRtz59U6BfacRDdDcrIQ
4kCUNIfd7EXs8DqXBKKeBHdQdNbKHjwD8B9rbUsyhnpUXnRrnd+dfToDvip4O2vll+UDhd2c7r4a
cTm4wlvStpsV8x/MyzBmjKx4vIzg79SAd3RXSB+LUZKZvQ0vhSV698MvxF5REWN+M69i04xqCfH9
k0iED4Qpi+Bqol7ZeWMYzEDlDfXgX+KmA5ifiPMrVSJxgs7mSvdm11+89p7ntO7RSA+pQ6rDew+d
1mqIw0n8pVyfmaUKw2Dq204RL37bHKz/TXP4jJKlmWn4kHo78VjjOkKj+jESYA3Fs9gLkC6kQUFL
szONRwwtO3Pvu7q64ZpfVE5S6vv5lEpEihWTtm4mLzaw8muX0rz6gVezawbqMSD1O1SZ3oNAeXmD
BIJfGPBzRgCPddxAe+dJGoSTwcytFzjizfmK1w6r0T0RorAHgCKF0yHYTKOmyJSy/pjaBm0/1USU
mSmawIjBd7gliKsanGO5v/mre+JDDB5j//XnQLSdI3xp66rb1ObX1UYR8W1MCutVVXYUiPB4jBOs
McWrappD5HAGWvmUKTFwQ/lSfpSKY0/smp0JzFNgdpoz7FpxomEZz9mujomfSplZyx2R3Q57liZW
b+cZ4G1f18qXDBC7duKsXRgXZe+djeW9QeDJx+d6MeO4H6uo0+1kp7CTCIsDYomHakG3PuldleFF
GedGizi8RopMg0OW00xh4ZVQAFquP9R8UrK+jqeq5qRQ5A+nb7n7IB43rwya/76w6MlV/FXYVkQG
Q4L1coNO81dLz5Si3wS8526/hDh7NLLocZlayr4unVHUP2Nb7nj34mRrCghf1T8FQMZyCXONXMn9
vQutXgshrcRCsoiXoxbOwTX75amYICs9Z0MRDLEg2pl7TIldPXmZSXsQR2fzHoXMB8ULaibRu2Hz
LH51zBP64oPuCd53CfRH3tSlJxIquDDVc0lbL4/QxNIb+IhycWHjOSHsD2gT55217MbFz3vqYPJS
IvQPRQvnMWxnelI/v6oIYDRW79GZBfu8gaHXf+Fk+rBTl8ipII0S8/jkB0HfyZIIRrGufdKko+p/
83ZHc+2QfgR1zW+cVK8WihrqhQuCLkYDV85Ff8D4BjfoTAo94eCOXQ4TJD8P0z9gE0In/Yr/JyHr
WEnMpyAKBNkvN3tx84m7vKAzQbJZk/4og5kLS/oJIUv87RjZXegdjPA+kSEaFqNvBNbhqi/tGeD2
316UyfBnB4E3pPgLWL4wE2mmiO520wFHk10yfNK7HYhQkgtb9wGjGwx+k1xBhnOiskF4IZCuA4c9
OwikYGD8LqZQiELdzxo+XWFRhUtJ9Qz0NLG7TLr8v5oeFGAvuF8qR0PBlA192aKWcOQEWSgLGNcW
kXxC6UA9ypzLMfE/gxb1+prRp9HN4cPRckhnZEfI94gxBJjrDxd6kXObL6cLnzZQjRPKMtUyb3Kj
53qKNBKv+tLlEQsTFvEsWXVTNtFkjU5G8lEPrQuNjDOkorqikkJH8c9EYS2Oy0aQRLSOkpaBkBhf
/2R3xpZEQLvYCmBdbQPqQo+cSuh08CdDPBWh8kEvCgElWMzqIfm5lNzgMnSWuYT/Pxy9U9sj7jlR
Bb4RLkvZFHrR0WkU4HkOW5Bn0bcSqqUt8j+5dhdosW6cE7+TW4XP8qvbARo2gORR4JdL+xK4CJ3C
h7HF/N3O42cKPJM9i1NYceisen+DdS3UeJqYb7SO3zjbknDJFM9cr3UPv5vxv6JlqpZLwyWNJnB9
PUc8ibbhvPrlG6Df/WBRbFE/X11GJWFNR8JuRZg7/T53gZEfz7Os1p/7mjr38RMm0GVM0dkyBUvC
PNJlp71es4SjSA5SsI/C4NB60BFsm2Z83cftdzLIAwfGXv/XgzMH8SYZ91vSvJ6W5ihTRw7tyhe1
sfwdEP0SfK7qrMFt+4PGh2Ccd2us37itTXKX7gySWB/fRPbrRwl/9CxO5mSX7zLzNa5vDdvKFk7z
3Cd6toXgT+H/3QrxNEimQWD+RQcrWSCIxIxaryg86X2dybc6OJ03Vfm5E5oncyMN+DByJiV/8VxX
/LA1DcpN3mwfQSKstt+LnH9j6ksWKTBeVNQYMXo4GLFP+AqstmwcjHR6VsE6gniDU8XfpkWB8oSS
7TifhviC3FWfZ5ml2FNriSuiJfN8T+JF4ZQ0j8HH5TrY2spGP8aK0UdnQ58xjhHWrwbMU6odS1vd
oOmw9O0CaWDanSpNaG5ZVIse+bpuIb4mue24QVcsM5zNo2bZ1tQH0IlwF+y88DMVUiDUYgu19o9f
wAdakYd1K3Ffix8rnjrbdsMbZFOQXhVw6UFsw20lhPC+vih9M8XL5wIh32o5SL9krsxNup6d5IpI
1ab6rEWmlz7Y4dIj9skuIvtDIAWlwNt50ExCAbwI0V1lFNFUSBV2RqG+no0jXq2OJo651ZQK8TDm
hYT0lXOqdw9wntzkSzviXYUYM6hMMI3QoHPcjXlbYQc/NPJy9YpDvN+E+jg8gtHPuuggiG24onfZ
kmznSue3eClWLIiB3ajxuGFtpObwECNIw6kVam3Tbya3+b43y0o3EU02E7iVcGpZUgyTJpLbOB1n
zsHiSqUBF9u7q2FfdsnK6jmGb4jMVbe92cnZ9c0y2uCeMiv2UV0QsqdL0ATTWAMY40gM6t6xC8sF
lmBf+PtmH4ZI7/D6gwEabawxjz+ZANGx71InBNX5180BoIsj3KRV2JraURA/TKFXisePLsRqvrtr
Cq3/gHRuvtHVUa9e810Gqj8WSZ2q/mXUM+s3vsYBiEQYZkZInLGMFK3+Z2s0sOJY1PTXOmgE52M/
68GhskPAYx/RiUMDFZBmoLf/HE5IBEkh/rHdSKuZ8olXSy4Hy1E6fmN5K4k//Qlzdw9JjhuhfohM
NRfnyfW6lE+3Y8kYP9LPCVeqHLMa1cPhDc+9PP9db1fdIgC8yPpoD50ZxxGOLXSpbU1zgF4Isrjk
XlFqrBmJAJBrSAtrI3/4YYMFXEeUWPQ4gjyB7llkDQB4Jt+9hbg1xHkXVaUi0CAKDqd4hJU2do/7
jv1msiz6KpBTy+c4zJRiEpFEQJKuthCpBpv7yPQvpyJCLOBV+FY12CRM/UJ8d3krRObLHTcM2mpF
ZSDq2wSOcZtLqAwSdJC9BsoeV1ZmodZ0CyevditeauiUpFy05TPI/QI1T6LBC2nGGk3zI8vQGQ8K
wkTnKgwUfnoB+9OM1Y9BDXcFCE6olpJZMb4GMUC7CCaZwfOs7NltSzX8bSG9Eg2vR3bxTLReOlPd
AHKIet3YmVeKdWC2GRhLrK29RywhB0f38fSX5/AyL/fjW5h9J2yeZjrddb6glCRqygwjIQeg3ru8
C6QpLX5Vju8T7EDI5faLGS9J9kC9i1D0b0YGoFZw4dvZ2w2Cdr7xMbLCH1C6yEGWWWyH6o+H1TSo
aYWH5jYjNDcwhi+bw50/JrGQodgwiXVK5pT+cAFZ+xe3sIAWkPXLwn8pLYkLDtW/OX6UBkDFzPXN
yZFcgmE/kemA3doTz4v+HRoGEJCIRsmtdrG5Slb8f787g6rj6fre64k8WF6XPOsjQP3D1XqPU08c
V6krcN9N6Knuf3ENvcagyQeLgAze6Sb6xPPrqJy4RIcdzk563RxoWYW4iAlScEMwvdthek8ST5fY
vUTQ5/syHn4y/biQHvUT6pVAbNgICDDo2vl4kulaKqRZG4/O2yFa75WsbCXy9b0jzneh9moojCQi
BaS20s+ruOEflnCziNk1lFAEFFJcNhA3wInMr+st/zRCUdAepcNTMhHJn0ifS5y3w2LyjoVBZqCk
Bby7ukbGIlexnpFrfJCKCD+p4WYkFoHkWwNcpZRIQ3eywF9mW6d/OnmksR8q42/xZQnaYqLAJgpj
M2MvDzDq6UOFl530v+7s6GkmNHmGQ/mv3E/RomTnfH5tcOnFlM4kgNVoAqLO5/haPxJqoA7Dun0n
cuWKyxOznYordpc0CF+uE0/WoqbWCe0vqUetSnJfZepjFPok5aJarRWx0Z1ZHtdv1LPFpsVEkGly
RX2L2KNYawLp7BTfIKIK9cljHD9A+fXsG6mt7bNo9I+7biH9KBA1QBfkuoYMrhMTvfSL8KeH9ztJ
kwxT/J31lZkvoQkFBw439ttat3sfBOOQ71naEFwPIpBzUyf3CI8mkAABEhltVH8BlBJZ5Y4Wn/5z
f0xGbnRFnME82/aQV+cjoGl9Drr3/coSRFXabAkeXfByOLkw7sdmYNFJbDASqwRZIm8i7NDuJptH
dCdsw7imoKV/ycFDL1RusKQfEPnWp2aCncbPYg/oFO/zerHrJmebWdf/Ho85yFaBQAOAJzmPmd+b
7qpVGgAib67SWorMy/Q/idw1GGD+jMeiW628IAYSlkpP/PJThJdbkPEV8xSv/Zfng9Fk9suBbasW
zah/8S1Kr4tsoe2TwqvBc+SnPOeZHydPQO8wOyVZ1J/BchzDeYzrbzDHwr3YXE2QQbyEZyjfgPoT
XV4cAo5GfLV5c9wCrdQTeRoXdVUtF4WoVWaWdkJS8uaAgHJ3wvm41qqaIDb+pZVwOeaYaRjUU1Wd
PvEv62E5QfgHZvihkt5Mw/gD5myAeOHgG+gT0O9p48BZZAye+T4O3/B2wBd83ytatMn+IyDI2Tdm
VzpUQ7XjYqGWv0K192oUj85he7KJcwEDnf2KIGCncc5889apNqRdcu+WZUbjVpiI6gmBXyB+pVXH
sL+SFkJtePEUOj60xV73guUbM/uEQ9sOEbZeOGWHRAemoOb+l8WUglOh6LjIIgSjBqmC0z5bmdiU
DkM8GiKjhz0f5Wuj/mLTKU3i9kpaW9etBbLc+6ilslCh4UEe7AZUa6Ic+mO8fiKBvqZiCodX3VTs
In8NAx3iujiv3rg/jtw1RooFQzAAysvK4YpdLTpc/1ETSDdIhwM3jH24zgUcOT/9S+VPjwc8juxT
2zCCPhhJihtD+/b7SxLMKKUdaaXnWOkbYEtZgc3AMk+qlKqejplEpztaxrJcOb/WasovAHAOptil
itTIW9yNWyOcrR24p5asvWSSe9q2nX4p9L8xod6BaG9UO/O3/DUOWYdkNBFRqIGaxOwfMwyYajZ5
3y8rnawXMreocTvFqoLweMDHDPllu8s7SaYkDRDKBkQuwBmSrneM1iNe39GrBubEzwkwAVBvMrRA
0FCzWWJCpjBPQiW3c9YHsWTjPyfwe/RqP54n71ZH4A9LQ5/rUk8AWFireH5JdEhT6p1/dvB/fR1D
6p7HIYmFnHMKwJYgTZtNOv06nRxraNKgdZrJHBdVADlNeM0a+jowPwIHNo75BBwmyE4t2lgKbp74
0Bqjli7pmOYiK0i84f3wmo3FnNZVXhWHfv1I+eVltFtzlfMj4jq8Ndo/m1HIUKKFfJMes6fKItlM
2Mp1bA7IEMTZXYZMC+RMov2NosyPiT/oeMKMM0n3Iowpvva2K7wo6bn65GP4lezzL45fSm1Iuwbu
EaO/S6u5LNvIcIw8c0KHXwpPD7CGtD6lPur93Da7WQAvhAHrbolcoADV7PxuAujAZZoCdwRcAqyL
yL3ZKucyTEo3pHHEuKR7YGX5E5Ge15GHP8GspjUjs2GcPqk8QIe6FwcChEFvYv+lHHmy/mGOnJqZ
jY/pfd85WaED2sXCLzB0DQCWwd3GpRwLC8+XMDKDPi+tMXFB0A/NRBZprYQcfbhw0IX1kpf1sBMR
Brol6OO9YujcIVZmhHAmoQFa1Mg/fYPNpe9ETG2+l84vZv9p4Ac5sXXpTqs1e+b5T6Kv0/wmEYwi
Fbk6PfqQBJ/ZazG7anGSwwd9HGvLyJKqtp3N8oaFYmI2hhKlhTC/UZD8hEsJA67YsvCxbqQE0W2O
6cg/9V39J+0PUO9eyjNxQB/ez3owjfFckBR4V9SaANooi7jh3OnuE8SvHoWcWQM1hQkspJkOUHVx
wDHrcF5NwbDcl7alEKb4GvulDUOIe72ndKRW3e2U3UoE7mkQFs8X9qjVk3SlsJ1OBeLlKqWPx7rs
WQXhirKcVuXY8I7j0IEO5ZItjo7ImGUYNpMvklHx96CrmZEwbvjDf1m9UYHT0ni6yAugM8b0CQ46
urr7SSWF+Hzg+/kF6Ov52JL0ktsCAX+g90k4aeXYzDIteNzr1tYsY4P+8XyYGipRcUNkoozpFn1+
nRBHE/TaNoR30xrcQ4oiE73tTxYiGA0ONPU8RAmgrgIBVkoaEunew4qDraTTpMFXhk5/pmqkFv74
CIToJvsAIyJP6Y8yNyEKn3JRU8O+m01TdeesVxyaiOyUtJGfVAlwQezHk2KE3yv624buLvjM6uZI
ZXlfO5TDqQipCJDp7S8W9fqsOtL1q+V/uoBGgKP9BfGanCXqLsNMJyEVxpocHw3R3YBlHgPp33R/
wDwhvmFX1yvujpId7bml7lg0yqjdjdLggjHeCx7hpMw1JErmguw80DmLtcl2JiqevctLlKAfjLc5
4WoLEwTtO/E/lk/PAkMwtFRbS4J5rmABZEJpoerghEcxnA4BES63RazW3lganldj+GHEpOAzTADf
wkhSLr72Dt6s5tyhbyjneoaQWOVWzK5WB5zv7mtf5fUis8FHugsqUp9u9zKbYidH8oXESx54GdL4
5UPalgZHYk/Kc1zPnKBLGfUEktZn+YzygZtOy47bVR3mnyKlwYTQ0YgGKyMPdZvGfLTCZW7pdK/J
6YVjuvxh1AQMQh6XqRsTkJrVPJiU/JxOfFzcm/vH7oIWp0tVkgEwAZXhnWc++iZn9JM4ocsnj9vB
dn4tXVAM/hqb76zPs5dxXU0RxL09vVIEG6TrPm1csvUG80dI0w4DTxyMa7TZxi3Z9TDkTcCSnCdp
KZZUA8nb0PTI28i4DLcqvxnIR0pUMO8TcHcYmnmtvwO8UqV2a4vO6Pl3+24EgBpnlsCZkNqLGs/J
GtGMpjtBctB3KeA3vYDwWb83x1Vdyzog7lPKPZrasdlxMjQfEJxXryLYDQk94A3MwaQs1jv3dDNk
jEO16V6vht58BMp4avCaNn/tGiLJEwi/k43gkez6sUqsTvtP2O8uDdxXJQ7fMSkmDz1NIBIxRIQ5
hf1+QAjw07UAizkUvYQVzfGVrWPFb5OuuQWlsRkgEn5MnjRoKxHfPJF/zRKAHJcnyRjz2kv/air8
tx4jppHLs7ozLzaqAuHvNeTbwNB3PRG7hJdAlp4CwfaRHoteSXAb93IXf6/I51jhHyjtvFi9HFCs
OE8WgmN8paRAmGUV7ePszVBDk2ikoIKAVWUUvALFcD5N/n2W+4R8DG1jzebYiEFr2z46+xh2lDmy
ZfQjt6dodoNj8w0/sOtMqPKWqOljRm7GK22Y7tJ5k7i6dm3yc/0mhrc813jQz+QwCLol4fwKjenT
3ykcrv26WTgeplRwaELheEdLhJz+C5qXLfwTx3CcGstKR5n1a+WvjCf9U4pX8YMFA90HK1d7zRa2
cmm7YCrpkZskOlH/NLsgGs/jddjev9/glyD9Izxf77YgHu/UgUuR8ZssCr6FbgYe7iTmWtkiESs2
KCK/chilS6Eh4etvKAdavcIPccCOAQ67R/CdKzpP0InWsDVv0Ph6Pzq0swapDBRHEL0TWjUPo7J5
T31s1Q6vieFTrbf+TAuAgfaAUdkyHgr14VqiUFM1Yhr7Rm6Bq44UyMEV1osCuXwBKrpu0at5T35h
8B9UhhCU2KaDM2mA2N3+kksuik1XBTM2WARjPXVN5PA8dRR5bHeXQWGPBs0JD74fWZPhvFUxANwW
aTKgivyfh8CJYObSpne54eX8uui+3Ijszhs+e9tlLOXZXAFN5tiqMv7mSfa/u54Mt95//pWXaR+t
G4l0dd9SikJ1uFRbgmrdsmisRNND/VEEfSKypNsnOWSP30IyTWQjlcEow5n2fdREKebQABI+S2oI
jbkbjjN7oHFm9STs2q1s8sQH+GfOHlZqXXJZO2u1LCCCENC10VTNsUB82le1+o95OjRwbpC7NmCf
4pY5xQYENlgMSY8ZjKj0gtKHmx3O26+aY5g9kl+RFcHFmILsDNY7wxOyWRImBH1ejbViLUv4dWgx
UsL8CM1aW4+xQliUWi+dgbNsxUJCBBRzRRO56aggWouDItrN8v1v1PVHqSP1aTo3gbBuFlCR7lu3
1mz5TzOC0R0G2QatO+W4mtAjIAP20dHIQzloV3N5ID0j7T6BnRQwpRkmMlCcJGR3NNOlNNref/oh
MU50YoTv6Sbk6l1IMe0RVGxoHhiUfkfR8U2lHL4k4Ft5A2RjjMTguDaPdQ0qaacpNXz9HCmPr02+
F+2xDYRN20b4UIv1TZpiSdGeQMnEP+3jslnK78D6A35Mdi8AoaYGYG54B/rE8IwDbCDeuiNpi5cm
XJd07LCTC/JEYcwJU9YhiMpc/C31t2vCEecEXXgIltSC+Pc/+PYU+ROfnacXAh5KzPzjtSfLC7Xv
xhOrWqhdJblkB3t+KlsEzGB9gtrXgAdEm+i40VHmEB/y5y3A54WNydiW4JsYdhIfIdhNL9CQSh5G
NcZXtDUUo6uEtPqqBBUjfBef2leMNBFJA3vfn+5qvbuKBNgva0gHhwI9uma/NbMl32N2borZSeI6
wVcCp752u1CkOyNWpNnempnUHyu1h0AsBBZRm5M6wUw2J27de+zjRq9n2wvJPHKeVSrp4QlfMVtf
vl2lyaxj4mnh+FX4NeA/66EffJmjMppaOMXMVKI3CtWKSxwZnwdoj23sMd6N+pI/VBQ4HK8krBfr
ljUXGUhW0R15+1Z8+bbUEJiGWoJo8osBiT3jJwCo8vtfCR31ZfFB3DX7F58tVTdpyOCrCH+cMWnt
uDgE97iJMo6geSQ3x93Iz81LSKrW5toQERZvvuUsD1LQ8bX8YnjBOZfvjUpmszw4FX+pCMUxakba
vw5nA0BTEhC/QWzPGKuCl9oNYv3PuuiFMzh9f6eHswMLy1HuouuKxXorVl5w5/szNjw+AHKcgClG
hXfeZvNZ26eZaSu9lxGRvP9cHN/EH37SWO0LQnh0d0QEHl2YmaOfuAeL/OOVp7B9RO/DriRR1KY2
1V92+8UVFFHBhrvSWtHMfXkf7cQ2mPGTkZWDkymU72DD87rkr++aQFaKwWJGPipZjq63DjneZOA1
DVg4VeDLhG8NYhec4XljXIFC8IFxV7cuiedzwK9XEHznx4ik2FKaTdx9ZC/++bz1EmJaEwz+dIEY
CN0TjR1TLFz8vFQrMfDoS6Te0lzZUHe6d0HSbH80xxnooEg0ob0grpPRYa3qId/3HXQ2xDjnm+rg
N4K4mRQYOgzQR2FyBz9wfOAZSkvC9DuzZ92C2Y+DOgdZKA8Zz05ROjyKqkFUabWXNM5puFmS5Jj7
vK61g4vznE1EC9UBq6Htl8yp/EUMBjB4HqGSTHUVNMG+FmtJ8YZ7tEgi+Tph1tEITG5yGlnOmF0b
kRzu1Xc2cxbmltLKKpAVbHW/jmFR3BLK5CaDnqEMpo4EZlNjM+BEnE3eJZlVXkpZFt209e7V2mE5
xVZFJ6gxIkIFTd2ecj93ChIKjSYW7BAEOlm0rU2PaxSuVQ4Jvh4JXfaVeWWB1DDMmtaJDB8xLTpz
MyCml9FDOgSFQZMXQpBc+Os9yeFAyl9iEz13aXCZFlVkJFw9Y4n9JFq7Q5HO6PKufV1xEpTY4cMq
XSo0DDbjNGsrQ7pdyUzrf5mGFzNrm8pu3kbVn3DjYH1UTWdEqO5tVgYQslj+8L7ul8pm5HJQoDMP
0Lsg47URI0sY1Jdh69BtfiMB/vDt1HrrtWeOBlX7XCBcDqxfxIRoEiMIypkYNUrbwaOzkgv2R401
MymG3QSXfoq2IDPZRrIur7uCS0ZKI2zmAS25lVHnFY5oTxrFKjPXM/MGM8han6qDGBy8gCSvRrux
IIo3fPybf4C0BenRL0q3D6VtRpnRVJ+WYIfNLhl7DkD6ZyUU/7BV+wwE1a94KCN2IYsIOrKP9WzE
zX+DDwubANgu4QCnyVaNgqDitIhsxkh9iFied6Yf+lKyPTwwmH96Q3TGEMSjR1zoCtcL9g+mnB4V
fScnl2HJeYhJE98iXn0uuN1nyTe5X0k91h8g1YHgqPqc/uRRjaqS+mMnSm/cBDr4yp9H0pSp0bLy
svI7pX3BAbGPr6YhtkCKNOkfM91eLQyicY9mQg3MQjHViT4r/VfT47V8eUC6Oibgd9arl3Rq5iq4
MKu0i+pKtbvAqrZio58MvL5nb31msQ9XkrvnP29CWK5TXqSjJwwIey8iCiNxtIIMWl55DwjQAnpX
VTk6O5ZHB08iuhunl0t3qer855OvXTVMpNCuhpOGA5aXh6zC8ecoOdxVHO/uH2ris7XWd43+8MK+
b6vvX4BZULlslowpeyVX2ELzcEiM+AyOusxSAB4ufSP1HJp33lD6jdrL8BYg0++CSFiyyAJEQ9zf
Bim8dRXWOswnwaNnXBTjTlBHYDhwB/AZEN+8ZV8QpU3CKYOxek/85P5IkZ/CUcBPbVJWBn8n5Tvt
AX+paMHSk6DAExrQnNW/NoSRXRUFY+Q3xmOFmnM6u7CLUx1oMaa5zWj9J5eMPvsiatK849aRiY+i
KBBnKe1lnlXgkYfS5G95erWQeS+TaD+/6UQ8lWUF9rFoz40wQFpO1lr7efVJZ7eM+ed1r7qqIx53
ih3ekifqEf+N549gzxg1EQkH2qZZb1sq1MhblJ+7zyrVXuhPorY3OndnE0iePYAovx2bXItoZav9
cKDpEkII4YFCwGWL5m3PpV8uzu98eLuJiaMwpCKbXjceSVZXBLOz0H9um4d7uwrzWq54Z+P91CXB
0uJxx4X5puC+s9BXdDUroVhrJwz88QqVN3XE84ZbEDtDjxr4SFzpWXxNy84RWDF3oghuf9FkoB/e
lepzc16iXOG9W29nBlTlLGR9kAEqR3i+Sy37x3eMrU9BE3UE5mixbOBU5mYghJJdx6/EykBBhaYl
MqDBRnnYUw8lan0V3Ikoe4AVzLDrL1+f1O0SdZiGOabmqSR1vy8x3Jg7jcepM/M0t/iI7253HHsy
RXIuudbxzr9CMJdBbu1iUywSeiNTl8aF+pgbpHs42lOf/eRs/wLdmZj/+KaqHK6ZnyObS6fpmeAe
B356MyAfmJMYcgo0xwYwg20RR5c1a0vEqLIXuvyZBDMazZnfD2eV5Pb72VlmbUKN+6A7IGxBccX5
PErs2q7V6oY4SVmh1Ak6JG9rp1WkjnBvulP+zEx1CaesONUqWvZrRmiZ4pSMMZAL9EcIYwpK1DSr
wt4+wnMODLNqqcS1TigifDinMhM0MW8ejY0YhjjHaCeRlvE8fvXr+wzbMhZQTZbj6e62xrm6IPLl
5dyqrHhe9doRW9MIsQ1u+4BC+g9gpa4vsy0SmQ5ae58iZ7O0KVDprFAkDygO+zkG0APiGnnnpWKt
k2hSgx68jInPH2kS2rXLNK9WyvL2JxPea0QW2cdf13v9KjiBgq9jTtWJMuL+pfDDQMAZbnqys4RK
6PRd78k/DXCC1yjZEYOXN5vGYK3oBXrDrJwy9yVTKVPVixHQpP4vtAEfYcCKDHILTgAbUmfJPKMc
qd8qcqmZGcWEkYKVK2EvZo8Lry28vbVAqSgW2nTBgc4tX8zzoRBqt0GNLd47jklY5/WMpUZX25uH
urGYypsQkOtUhP7WRF51BI5wAz8+9qJ6+8FykTTKD8dpBPUEleIj1xIAn2rlsEYfA1kuPQGLWrE1
unto2vVM5/AvxFy1a1d3W0/1NAEvXUTJrAg+Ktykaf19Y65K25LXSNoon+gPAHJdbvrC+8NhyhLj
4j76LbADTfZYMNo+qrGZxXvrUY21Il5c9iRPQYmxLo8rmTrvhn7UbUip6mVCiV3nRExdxAbe4fdZ
kPMBw5eL2hlpFnpVmhlsNH4q5V8ocVh8BLrRcq8/+EEPltWlLbRG93XzqJfimqGFdlkZMxNQkBuh
XYLm7LiA2FUkOaOabCh9k3R/vhKyBGsYvng4Km8oeEXqnD2KtxhsDFmqPRx5b6nQjRXNKQYq/O4v
kjO2wVG8Gib4qqd1fyzarEhPDOvdy+6JC462y6vRTE1NhAOFjkS22hV8Qz1LRDZvMMYzvnECuggP
9jLXAHuerIMBBGzMSLfU9jJooBGRqfczbUiX+XVuKb2HwRAnN/Q9JvVVEbOA/wWeF5YojZHwEBg8
ewLFKbrn7GtVYuRNMp01+xcg1qSszevyEKcKEDujLmxYnO6DTOgOvnltDN0E6HqtFn5grJJUIzbF
fuD1Ims3/3dlJmL5R4TGbTZY2jTE/LxeMbgAGMXkyFvSDwIEiWIwLfg/Ta+vdhgeS1WY3PXFYtES
VbCNE3sMwCtSQHr58mrND+ZJOQu5fEEUG8lFRYoLaCWtWjybPyyxyOa++X6CfK7n40otpUOUOLko
qgIVjk+ZOuwqRucyKtpTeauUscDFrd6N2AbMiuX8b/sLqFiYarsLCYEtwCFi2ixfPDH1hxc+tURR
DLmJeFxDNJZG7RtarqP6g76OP985GDxATnJknW2NlHPFn2M3ePyzN0lsGbTeN4JXD/5twNWwDzhj
HoMDS9o1MOJVCVA4SUIlUZZ3BwddMH9ZB+44QBFmy70HELtRYN4bLxAoEgaJDCTx6A2UFietkiEa
djnwxdk2i1Obj3gKZkCKZdH/lzoa7PwIR7uuV77+SmjL8vehc9RjvIA/IXDOAAIaIajFIOL/LFGu
WKROpDSiwl/GgYTr6AeSgUXxN6i0NnbeUy479dLxBmX2kaz9G/3Ma/7fSfSmJ67vgGgtLLDaTcAs
DrhIZFFhlLcVTjQQuZ1c3VlajgFHzWzJqLOInxSZyGVCqgJDD3W1dF3aPy/JVhfSYmHk6iC/di7l
k2lA/FO3SqvANWweMBGviJrpHZ+zJzVT+NwWvEKDbgrWwzv3vrnmdBZxbD2+JIFFMO0sdzpMn3KT
xo+iyAOwv/1onwUPxhyBG5oII0berfpnP1fEDwTwaPp04NnNFz5e5FuxVnRBu1WjF99ShG7AHDrv
mLC9GC4RFcuJVKVJ20BOsOX0kwQFKiu50EYXuNK8e3f59bKRd9CumUmA4gTTFvboMNBnccA1/yJX
2A1MEqOdNVIw4HCYxs29iYaPPxT0qgUDKKiAlsuibUvHsaiwLsZY7EgViGYr1doJHcIyXqhZ2GQ2
gE7qGOt56ctPLHU2lQq4yh2/wraLtLSocIujQL5/OEIPToW/tXLpLVO+OprZ8T/Ke9q69lZx0TWe
P4LrIk0WOGfdFVyYaKce6KyVZdhgSRhdscRlqaCO3KH6+dQEeUBcTV7bSFXMAc6befEUs/cXM3Tl
bp7xMIEe4h+P4zFxX8IDCDJWCrRcVic0ttRP0FTU+LjXiyquJjsyfyWIagsIcERUYUP9ueK8ObWh
xhcHciDQbZHOllegS2E7CQZFWIo206jeKKXNlnqiFX89nCbb257vMKkawSRUK8MQQqK56hUNTj0K
ubQVwDhvXEojUUDfvpsD0cKdQ2JoVhfm7ZZ88ytYhNjQQWms/fuRDDRdobhVyX0IoUF+2X/MZSn5
b3RrlL97UJ+3d/df3RiP9iQtzo6U0AousBjoGmMUMD8b2jpckU1QO+XElMRuBomCYZKKb91Vppxh
0XFSyVcRWNJPv+BXwY5X4pGRUSGJ2uMuyFDJ04E5yG/7G0OpkzjxdZ73B2jc0BzlPdRR79LPmwvf
sZKW1AZM83kDXh3Kr4hYKkBE2LFGCbCZmuZ3ESi7E7+YD2UppEDbp4aSBuV2Y2ktnFt4+MyWX7sT
p/MIE8MBDoa3VLiKrdt/lLGbNnrmraJbFq0kkdZjJY3NVsH9C5m46ZpZuhwFtH/CvWOY9cRJ3KJt
ESX7cBIeXCWhi70nUhG9ak/h53i/4WGJnUhOYX9OLsp3qYxEjc/v0B/+fNY04qrmy62O/s/fkjY5
deH+rodzbhzSgUxtZ6y8elbnDPKPtn8x2m7U98BkNP2h9caAkx/e6U/7iILND2W2mudSCQxCFAS1
7iHnu6xw5WswCbo1/Cy3n3ISE33Cvj+zoVCxYUw370BjEAjigehQXv/kJLDsxi439+T5u1VBNOUf
GKUah2BnJ0ALuN26wniEC4SKQvOCKOiqdz6KAB5U4Y9xS8HW1lQV4nJBwIe+/MknmsKugxuphta9
Xm+1sW3aTvienxqdaszje2RZgQHWGvXToRDpZJRN5I/MylyZbh7c4empD+RFa1PAmik1fibEQ5WE
BmNkul6zwaF1xGDpiysb2VjnbTuAQM9gTCq+z6dlJzl5SI9f2vypTItbzhXPNEjWn7aIMzlRCk1k
1q6cyN/fGCxsl5sajd9Dt0dJ5CxJsoWXgE+Gpc8otYqilQ1gXfVYuF/Ps8/LRGzP4OLIljhsEZs/
BXSvYDbhTWtpBoVls+vlCTk7gZkSeCILv+3sM1NvkXBaSP3mkIHf3Xqqer4W9jRSj3ZCIwyVHGj5
VWSUZV4So7qZQ01XeE55t/C2OdZzSjtdGh7VjFIuXBokMqZuJq8+PDN1Ci6owx6d1imgItfDFqWd
cjA/7TjcSvsfKEaljrdULdRVZrqam0htWvI5ttZxQtsduaKAVZguf+oQOzngqt+GWcUPRNJXkLIV
i/xvjgUA5/45WG6teS3saD+PiUihHpy9zQKQUt5oq+LG8Pf4RXMsqXYbhQaWR+KiwEXWx63tHg2B
wHADfkq/iyzuSiVf9NxUKIhwycO6zHXnUeq5S9uXRr4zGVLHmtUem1yWQw4Tgu/Dj7zXeCCtLMAk
SbBi6OgPdN8ZmjScFUvsA0n4dt7DBKWUHg5nj+0+MC8xsW8lcTeLswjT8mEYDpEKsn3c/nfU9HTY
BmcvfcepRuFmZL7aJzyW0XP0Wye6YyQGNZORa3lNb5qfKNtWGAoc+j4knZZE0j97yOBQb19P62+8
IRHi72AfgOtM9Sw2ylZS3RHz0GmStAj/zKIfGgyVgaWVcIu6ayMQ03yFxDOuJhnvG/aEUAK14GYR
cL8B+FRmXURfZTbavhGG3RFwj1MwwdC77QnQrZQuz36fYpp0dq9CoXA84P2DQWa+R6QfoYrGKkz6
CAk7SrWcEiSry58l8GKSc6o0DlepZHLVr/SZymIt1Q5CJruDN7ZD3Tvz8Wceg8LukKFJg5vEkSOO
xfe/VlrmwoR3XglmQS3WzO5SFi+8EfVRUzvoVoc8UUI+6NawCDAeJv4n0SdJubYgf4nj7+otEdfk
WitbTsLJ1slDpwu4JoTUw/VJWjyGxxwjsG23NZbl1EQgQy2OGy2UFnjbBwbdJVmyE1smwiTnJUqG
dMdcLyf6a9sv1MfSHFr6B2M+HZQxnPboDaP86Vj8jAv8TCpVlfQjX0BxzERVY7cAz7t56vBd4Hgh
f4fyd/BPkTPtK8PKuCORyYRsrAPHQu5wQfJFMinkU+JTs267QWzPirkgcNK7ciC2kNKlJ8SJMg9G
F6JeQHLlU5XYxNDHdwblJeBEQCQ16hIFGoaMaV2xBIT2ox2VIHi9sRoryoOWjWHVR60SBzSZZZMd
TwNuZTnZfOnoyv4oGxoN2p68VxJc26ov1VxSwUnUbxTrlIpMeyxxq7MwOWNO6l4bhPiMTqMX2JF+
DA87NCG0yFV7J8wLYhvbdX9WGgFErJbQCY+NSJx/+0vDnwbVXhpcX8sHEwSohvC5WUGVM9AMe6ql
PT8sMLRlk7VI9bGUZAD6cZY/TcHPykKyiIJmCxO4cLPllEwcwmsm3ucGbKNNlaD5q8mbQHWeogoQ
wUt6eBp5cgNnbFoT5JmDzRQS2tgOkbAM2oEe6IcCfUNGe5CKJxQZ94JwgQFNaIBWBay6MoAsPjjx
t2P9g3pCKB0VEoqXD3vctF/pwiRQO9GDng3VS7VvjWSaZSvKWhvOQOH4M2RHtIj7WtDYqxMglBO9
fQNJ8lEbRFo5lMYmp/YUx4jLzdj1vc2CbxBsmi+qJcnUWzD+dN9Q72yDMUf6o6Iea/SW3zt/ONfP
Qro79jTEkl3YNVdaCbUO4p7XTZEYjD+ORT1Pt6HvYEn5iHBDd3f+aFjIgCkFzIhSDwCrNlur0JZT
ymIqckrOCkEjoU/osGV3RTW5VgpqiPmjzqJhzEVg+YKvKGnQLNU+jbhhoaJ16Ko1jxM0IF127UOi
+VEfA3Oy7vv7g0Vin0DntQBsgq068UhzfN+7VJFJwlujOK/GKPyeUbWus7O4xbDMT8pXplDZ3ZGj
S1ExoCnX0dB5NndaoCN7wSQZc/6P9aYmpFP/7R8+kt5oXOOEKxvn/jQXSOjWycKtdn9WC3uYN6a/
t+mGOmSoXPhNcjdIyAwC0Sj1F4BAHmYqhTKACGVrkm5X8XjBPHgmK1ejpx11li173kFCeFcqO9RN
BzlaYTUPWXx8gO5LztV+l/iT3LWOJQ0OmcoHFX8bHNuqx94xszJlimtuuQ0Xbke4N4p1Bhjr37B0
Vet9mxtSChKyNEq1JjD2b1mLlKKlxFAkRCQAO1N7ZyE0K8RTBuigDLO6N5CewjU90kKlwo2nGMER
v1qCgsn91I3A3ZvAAjHAwuAnRWIQCp6MAQ2t7KmInwTnDXxkxIfFMa8spkAGecpUhkIfBa/gcg3i
tnX7iAiDtRR6P0iVzXqlaOlDJx3J2jDFKz26/z2fGUG5SeIlvmao/cTN8/mFmItkcRmN9zuDb1qI
bSL+hVmgWQ0/179R2vfWK0PZOFPK3vSvg4Zu9NNVlGyTCs6XDTlqiikgp1U5Ob7J77xjXxNy445w
Nf3lt2L0okH7KomeZM++8xLLnb2JZvXYLiPhudLYtvgEBTG4tQwGRFyYnpw1UKmOQpseaLL+6tIa
CcRM078A5Fa7C3/hIo8TMaDWnJuh0kQrk9r3cY3StiCOmIy6RbPQktE1CqAxprgJL/jah/jS+zEo
RNPatDXD352XmzA6E+n3AyQ3sRmOfUkC9Yf3Pb0vkD8e6px8VHSEonoGH5dD6YDCiTJ8C9fpL7vS
Lb5OmdkApWTiC6d8JBP73bdTkAp0el+YbFTsfh4MJyadZ2jVFtiI8BEOk+LTtgujNDPHbagZ3YcC
jQ/PJ6Sa+/Ccqlr5inw8EdPCbXk5e9EnrbSCMy9J5QJ7v55D+HpzqpmaO/C7ZzL25yN9DH6R6y51
JtpnqXY5pqajO7LM7I8Dxz3ci8y40uJRJgaoc5/XHInnllHWySia4vOAzfJUF5iaWxQKzBzCJW6h
m3F7ezMyfX1gWDPOpdloWMnviPNcAwdvnzuPa8WH3Hcw5gvJ6PHgF+RQcGeFootaaW1bq6EJYAeV
/+fWtY1OMUn+zgwcICqaPSeQDLgqVaXG2d6ryuynnyIhEOmhE49GMNueXTcqqE/q6mqtJP+DJDtc
HUQSHiRsygK+qi+eJ09tWEr5tP8EV/jnkD8w3M7oskTN3hWwCHPBe1rPAC76LXcQbB9/BZf9XhWi
5yCqP7eY/rJu14A2w8taO3zTJ6+4FdW+C/QhOpdE6eR6dkf4++bt8ET9v2HnjbCJar6+OL6zVrAh
GRkzhZL6zpd4qNj0sxt5sjodc4p35bWdqn5lXE40uI+Ps08QZ4szINL2aUNAwy2qizs8XPIQpsE9
R2JqM/s+ohXHmC/op6QLteia+5Q3DhL68r4f4pQl9WOVoPndaO0X3FePqqrZfWGzN8tZ10XArVit
t746YviPNyf+fcICssNyEpPdojZkho+1KdoaYL9ZMGXJZbyg9QGO1wpRJoWO0qJZ+MZK7X1FhZJi
MafiFSYI/lepWDTliFju+GhTCC5GqYjhjm3086We7jYgo8BGQRxdjgrNc38O7zo7OMNN+dKkUASJ
CQPuwcOjmQSrmutYaSaw7QxJkASKI6/fYiIdllVX/ojyMoUyOYX2sYBMHWeqYE1s+00/wrjBUbgg
V0h0Rinb7AqNqhaczIZQKLqBZ7sv/SGbSWUBDZONZRHO7mPD6W7FPPjNXtIOkjT0HswIxHgZKRAY
BI28OVfzlXgr8XuK9rElr3N2GoOzLq6lSSVH6ML39arpYXwMm0i9j+scB/M3qVIXDCFV8A7nF6MQ
1U0pF83CYAB1g3EsJ5Y3yre/oKqmEI0SS1DSJa6UhllA5HR73rSsRH8QSADIWN/wawVOrTWbk3aI
3xYJw4mZQqEOZUXwF65Gc8FhaLIPztehuFpyIomgP0lRYK70W/x8zsIUmjyZBG/rXSUkn7byxN1H
eOEJGbkh5W4gLdKZfWX5ot0ZrOkb5hMUKKiozVsBJBFXUqbichLZmUA4GPDIJfHymBh0g81w8iIs
ZmJzQwlxHtwn6rNgjVo0zuBrhA3PU2x61gl0Z/EiFoANo3C9AH6qW+uGxOjzR5a0/tACC+FhCuHc
E6wCo52fDPSu1j7yK2IGVVPbdoQuiHMAS6Asc+9oI9M6gc9NqLdobowUuE7qSmkepG1wGln5wCMs
c9p/eGl2deSsmIfC6J8ccaBjKmsHIQ0iyi6ggd1K9yYwY15ZpysJyODUGQtmLeR53YYsh2fMM5TG
efzypvApt8vcKKqSQ6Vk4ofVlVOVLI6cQY7KC2lr9gSKYq/n564hy5gIsQbsLzldHMkeqNZd3HCZ
cxvIZAgwzPxUhq/GDy9pHWOXp4UGvAjP14JI5Dejst04T9MoqYYGqTdqYhii4NG12SdsIql29CJl
RpFK+aeDaY+PJ6S3LnVeOuswGdYfboWFve2rJB9Vn3N+N5L9rDT6al3cyKBiHxZfa3v0CUAfx68h
QCuK6PvnkD54x4bBAS5xZt+rRmZyvYK4WReoI0PPAbSDxVoLuV/ZSZMjN3s0Ejiavt0loccmOe5J
uRgZWHOxgjt4n2Y++wayM/MlyZcN8G5L++nidah2ou2lDCfQcIQSwH3p+J+Y4i7S5h5irwvurlh5
1L3wSp/Fn4pjqeISe0uPEdQwm9gWbUV+cyCiXpkBUw9CiiOnTf3zc08XmH4FF9Ht6VFU5JvdZtGW
FDbW/+Q6Pc0yt6yvWYGNYEWOwQ4iFqvdmAhBffiFS+t9L53aT5/bKsYkvycJrHZm8FHEdloKDi/I
WI1KCzAV6LYhKGRbAEP9DEu8tl3Bnfm1f1B/oOXGSdqIBe/TyEQUiTvr19CH4phg3wWyD0LOR5gq
WncjIrH0a4J+6IR7g84eBy8D8x2WBhAZxukjH2BNjQpP3Vf5FiLIXlPEJc8sPyoR7iKTBAEh/8Ex
wSKoiJx4beSEcy1TlroD0klbxre/dgpS8QgvxafxcCnp2DOKDnXxRtZ5T4pz8rV/DJiVtJoDgmLD
Tt5als2nJuCNiq45MaUOP5M6sv1wrcGMisnXJP3UpqiKEzcibxNMCwmLQs3dCJdjyzn5si1QJQy4
Bosad3MEMvCDx5zXamErscRUZSioFF6JdcIOLEu6ZwXPGZ/cIy6HisligJznuOA5/Y6BOpGR9mSf
tuETnUnCxv0itWLM+yA4ABW63MtBqyzKN/NE+XELA7LluDhO36vTBb7qvOct0xTMofr5CIyrguZu
XxiuuiAkS0Z7wYDOkJaigZ6yfLYkmSiyBefdGGZ2dnU6T823id9frweb2PXlNfzponWbLJIDniMY
xGxOO7K7kZzjASkWsLyd9rIcIP0We+JFp87mrPYVGW1ZSDnJLrs7nohOEoMxyG13k5SjESgpaaRQ
nIcRMlKmBKZddSr16Hkj2+CHKYFnKVMkxx6AVP+SzXJoXil8/L5yQP+mnxwYf6T24WzWJYMIRzO9
S2H/rXqzgYEIUVS09BRzGggYg3yPlF57hAEZuAmymn45YlOU8P4KUi3cxo7SSxrVv5yy+6w33nj5
YHGIMbLYI0Ed4Y0/U/LlxPIfXVWlR087ZCsdc5U8N8P0xNl/7T/Ofdo1OToE28kg0cbsBG7J3AUe
Kyl9wqKQTGyQhZcuo70GYQASW+JwjgbbGE4ePNSRugHP/2FpSbsJ12wBL5Ip/pprfSNcYs1AuYFc
Pee5lICaF1kSNNzK/wjGVnBh7dI2KKf81oFFXaRUlcLQwqnyEs+bGjlEZiXfWM5an3vKML483IYW
wlT6Jj/F+s+ztu9a4YzhaJKaZMfD9y+gn2aV502FKv9y4OqH1ZKb2CIQhODtu3wQWnABdQwGE9od
TdasJH5ko3xtFsb/X8QbUolzD7eRLG3A9cLMUVj6MyMwXoU/eYuQzG2A5GGlc4eTJM5mfhjPLi2b
szOKkW15Gm3LH7mTcO8xT90SkmzAvJtjl9TMLEtcW8lFD/eL8nNZepbnrasZSesil8PRRnvCu/Iz
KW+RLBB1ShCC1lYiCP5Jebs8uva26Vckea3LNLcE33ztyBX+4QEE2KSD/7yivlYIdsEjTKFGth0L
f5snSxbbT2brqbZBNUyC55u8BEe2Zh/0KQrX4C3G2rMs+aRXaXfp+td/lB/RoSPYo0jAWJncadbI
f2zPvune8wrJGWeJanacadqohEqsApkk/4WofRRw6GLxTh1Klr2BgNyl3/n5iIqhiQjbcsSxo0Ik
RanrfzteawV2XsOCp0BqBp3olouBw8FXzfvoZBNfAzCksp3TgGbELD+XvJvWvpetzljhw53BLaul
1TH4fF0Q42XtXC+2ZU0N6T2WCptmyCrD+KcPlX7kexbt5D+g502tBmPM0B0fZdqBbrtDjK9jMLZd
b2Kj/h0z50Dun391rLHVX6HM0KHu3ktuA7yJG5zGrg1v3Q1WXLeltYCZtwomeZCFgS/vdNpzZ7tu
tOmhDOR75brhtcPcPdGI7+3nXiv1wlAl2JNtpy1vVTpFBgpdewkHw0P9X05uRRsxBRkDnP40aqRB
ye1rD9GRAjZHeEXfz2x+RFJBkCCTXW58IdPKfEGI8nOam0kI6k7rAdX4NnYkfSEpwS1BvZ23eDNm
WioIltNXNF7R+TH4vU0uYnljhi5dM1OOiPdFaKdkxK7RHEbQXV8+H2wMkovh8n+IvrPwkxlawiQA
9LmVosab74Ch9pxmenFkJCphN9lYvkuVDi2K7ziCaTPUXYccUFXtmZ20bFI7CO/gDRwZuKfhihGV
3BlBs4LrQmuZGqZiB399X/8RW/2K1boZFS8qnHJOspk98ZTzsf9Wj6/RzhoyY94gKHXWXIpT7UBP
odr9sa1nibD9KDtYPd6MOMlHnPGj6L5PGi+/64MOd4GuhBRpmZPTeU/LF7jymW3yvVpisyqoi+L2
IcBQ8oS1hHODiW9ukTzDiU/bQqs3jswypM+aBshSMmD2MQkt8hQbVfg3sFSRLz/xmqQtgrzlqdwU
O9w+lQuVTVSxskx+e6FpVS902qTBQQholP+HYBt+yfXblurYLgcpM1iD2065ZhzMHwte0PFPQPL9
Bu3HY9RfQoFAIt4L5o3abX3zzkhA4/sy8WTv61NjxFdcyRfwjGSvMWzYJr8/sfHdcwa4YhidPJAk
S4IVj7nTAKiLL/vjLx6pF5Riv7UFOzqc9BoOnIXBzK2K5putGR3Tm5eWmKJVEihg522AFYmni2E6
Cu4rHg925EYyWyeQ735zkBqitT5Frw5zJwceeMpPBzrkUFxiCoJcXZnfIyiZ2CH077m8RMbSInJG
FVe8d+G2CscLSL32lnhTSEM796a9Zzbp4e06jwFD8FdME0N4LdOKMtoqXs+70GkmH9xvgve4GfJm
A4a2sBYlmWyROXer1S6wYf0YiwnhvsFp/1Kg87HKwZnJnpA2CZZvB6GlBc9YFUuDTuqwOYPQUr2L
P9ORrD0/uNvW8BqOm7wAld3yJiPm91dyfrCMM9h3OLiTaNtXab1QhjhNeh/m/Nfh+56pZpgpZyqp
1ltqZii8uxu62yj5qg4gUNE3kDmR3pYLV1l7HwwNhIODdVJ49q4XYKPgRPwsghvlLlEXnP9G6LzA
8aTuwCdQMZebvc91tqx+qu5X4pDm0RZzNNlAnpOkF5YxF1xWC/3KVV89+iW6Nmn9bozCChk/JYUU
yMkqkPcODDjd/z+1W0yxW92zPaMIU/D4BGg6GYo74IFS+5dQ7goJWKQzjo1/TwmtY/eLJOgqYqgr
4P6Zg0/zNwwrPId2Y3OVm0XsmFejukUgwl/nSd6FtYA1tnOxo0WaBCtqehMFqG68gHPCNtiHXU9s
r+R2qBfGQLJmI9NTHAA2nTKCjcP0tSvcOj3l6Y+tkd2ftv6C8pzwCVatUMCBuSI10am+QQ45s38Y
OAKmCaIxG3S8BQvfede2jwQ4jydbjORfRiBI/pF/E11QpKckli4BalSswC+KpA2E8frfm7hV2tGk
nLYiajj0AoRsZyaqbb1IW8Abk1YFYLGZBbsFQ2XBjU3k29rkxQ9dhNeC4kC3idq8BoNbjtSLkjua
9Xj15fAhUcNX5glfE1RqL/NLDlSH3cKAEBcCh8AGDOzH4dDAYtyXEVknKj2Ufe+pUbOCtW4d4Vgp
ZEzuBvChQIw1nOSYRrPvIlr1CFfoyedF5D75Gytm24NJxKZt0eaDF6Y+YFFDyYUjRU8qIDBUjpGM
UgCoR9McmkDhwvKKXEMf/W+20tiN5A53BbJwVATXjeYC2bJ+SfZCNbquvRXwIQVZeXLt0LgRrnKk
DVZexE/Pve0P+G318YmwanflMYjBMs0C8DMktGMKsylUzq4q7fyN0vi61EbB/LYIjmgRD+TOf4H2
lqTqECfbAdGc089zKEzHD4HvKAZbk/zlz5fMCkWFWQRCewDbq7MAOm2HgRyHJAH4r8d8Fcqia68q
M+MJroqRN6JN7yymSrFQEhjB6+Bk1MopvAWm9By3y/u3cEzhpjM5Ef/aXB2CZ8RdfreJJYzkzt5e
UTHYTbFel4voXMbLmBoFcsEuSR7RdiNGDjKzNXmfOHdoHlMg3O0sAJqvvETaQ/sSyrTJyIQ8qOaP
ZgTnrliqe45ZvGpSSEZb+dlID6/e+S0HKV+agPYhDWCNAFgodf8oE3xrTfL1cDn/y1+MB6hvNDxw
C4Shdk/bdl4zNEnMV24suXQwnYa4WjgFMWl+bGiHXTnzGmLGOdKmW7lVMUDBAsEUmxTVDZAdHmAX
Q9sKe8aRyH7i0qnthIPr36bsxIlNetq4x3aueHPL8UcWBM+U0a1JQBy+oP/uxPX390BOgQyjguI6
OdmktxdDe9xDVhzwYNo8lK98cetLeNSkSZhThtZNlUeKjxAT2BHyUjexRWYN9lqKfAppuPXfxlB3
n4NFN1IllYdE3n+2fp8VV5uz9gQC7zVzGsIdkKMNfj7/wq4o69M8HMKc9DKsLmjRwoyRhA0CFfPX
e1vFHfGMXpUL3R0b83tACQHOrmNAJRVUR39S3nYTKyAMQlMQaBUZ7O9SIh9Q04tvN1hDuuzghPpr
GImkOrVM2611D61JKgzjhYheld5VJDUd6yw/JLuUdHjFg7jDkC6mgUcixWzdnNYQGGbG4dVm3znT
SBo5uy4vh2JUouo6saMjdymTRTVsMXT5LKrRU3/KQ02FlXE/oBUAFabITMG3lzb1eDoui1680dRy
9mz3kPrA0rPoRos5BDA64oneDnGeiM0zBHOGNE+68NAjzNRDUoakGw/SP5PeLKKMWIqK+SZKm66/
Ltr4S0sjk3H7SAEqPBRuVrylZReJLVe0bUHnlWcoZncOlQak24vOz5YX7apwX5pgH5c3d4aOzA9n
UC4T0thYutUzNgeyBa5DaI6IwxrmhnMXRZnYDmuKv6uLIsPNmqUi9Et9QWbKcKC1hI+3UTDQqaMt
Y7pyGbNAVm/5XcCaTTyHUfbvd4eMJvLz57AAMBwWsFUZk9WE5UH1RrIMfv4P4x2PHdIjj76eyGtV
Ray4z+XSYnMbvolCypGoF94H+N+sjfzwZ8K4+UCQEO/ewmcP3tXlVMzB9GNcf6SvJGe5N+ZQLDPh
UB2vRHHOci10955rbQ0Rm+YBsN7m18XfhvkEaHzqP+HvjoEiqIW6qITtAzXx1p9PiFv8thkX0vKN
x8QWqCS1dxHvh2Tdkujmm+gRWvzPKz0PRqR41dZdDcNI5RWJZJxDrzTDgqldxW7/UKcmk4zsnk6A
KWnxS+L8vfIrtczAn5M41+OjqgTtLjRK5eGkJL1WKnmvreby7L7I+ze6VNxrfTuNgLordD/4Xdjv
MaV4ZfyB2Fy1RJgl2+ibqFpeDGNOFZ6iqYxSAsDxsbi1jZ/2MtKSja15kbyU+wILggwh/HhwRe3v
+WRMe5gKCTNW5Dmrp5oMS5Zfsg9guTvG6YQzCEV5rqZyZLiqK+w318CV87VdOqUC9iW9/9VThR4B
va1S/Qa0M02nainQTPxaZXR/ghCOGiNyiusKGWtHGZ07qyl6cy9bA9c7DEwySnXvrM83nNJAyIfs
o6EenBawQIx/xp0sDAoPHsQZVYB4gJB7Sh+sLgVUYLcZeIyiaDm979US6AlMIlJfZ/mgIwd+07Bg
Il/t/Fj7hVpKV4JHr0ux2ivy9vWJ9PrKaPxH7R7JwVLdeTVyBluP7MUoFwZY3oehxQIpWcEPoW++
ACwmrlsrCQ4JT6L9JnqphCqP+mtLo2AY5gHs25VaU+IfdoYWCxftiWPeiYOxW4pjlvG9Zx982CLZ
A7tODgtVKkTeoyYyyJBLA8bX9fxA4jOiEhiefAQ1Ts2aWQaLuXA1lpG7nl/2lH9+lEoDtCib/oiZ
Moj8ZCScZosIqW13kWM0XiPPsDvDcxVcn8ihU03QlZXnsf4ef521ji1PE8NNaCPWTHhMswn3dtQE
YFSgsX44D4PQKM/aewvMGqPHPpr6CuPwVjw5twfjR0l7wHWcduWse6oyc662dUvXislJ0qMl63hA
XS1wBi5CPEXrDHsXM3rrDg2tv4uhXJt653wR8/9lB0BcSPmlWlFe82uBy4GZlgOIWQObfkiFsR9Y
TkJ8g58LqGayoeeUj6gf1QGHmkQsx2yqyS+PnxmhZktJUL4MpGRuQKcWXduli6EmPFJe3aZ+2kjG
9E43YC61fbGE1N5pw3qS41+x0a6HqC3EaUzPKSth1QYYiT9sdQwjOUCvnhJNZof+0O0ZJbBMK1gL
Arnbc1dq7BYAYDGfUAraO7y0ajxt17gXspPDvFGZYCCkMZXcWR4EGOlKq8zBqmsuN8UjQjIuBqfL
RJzEolMqz5TfnbLYRUbVV+RVUtUN3LqqfOr/ermdlPAisA0SankBAetpxoeFEXGDFNHr5Hc1hjFp
evhmyGwI2yfrjbSBG2ppQcBmYEjUtBKiivKtF41v59sUp0oQVncLHQnNmbu7lTKS3KP+aZrSpgZ5
sTVZs8vSq23XV5sO398FNZBtwVGR2MasSZfW3iZKPduWLh6fTz6M1iMhnIO/F03/H6E2qo040tkY
SRQA0szren6ycLqIm8/yg6JuSnUtfdrNCpvZe9odrisVzlV6oZUa8VNZ6YWvoIxST0Gm9Jow0E1p
TF313aMtGLojfHfZr5Icn0DX7BYRzLsru4mORlfzgBSQVpaUmiGFwyjd++9EyTiKlntBCZUOPdj9
YMcRVk4TwnZxMD0yc+0UHQByPxYCdEA3/jbKPh6qblfmmV3dTorvsfScA621rSA/HOWhkQdZpapH
GhE8DuQpdElAgtY+HmZgDMVrDUen/CHaB5VbUTPL4mnqFABGCmhok3sGZmakNlawHsvYJLwzSHzA
naO8d30UasMbNJbKwKsTr9Schppfwoq3/lWQHYxcu/TsW73jGTT89rgkcQT78jN2+VI0xnckKwn+
thLWcnRov2qv4unB5etpGGfzZJkQFYJcX5QchBAj9wUYhsz5jvgjgewDUHa7Yh+HwpcrguHG5r9L
8EgMMvTLHlkYMpID4iILtBoa9gAFcb6zNAzEDmE+RWY6u4MsAvUtJK5IrniSjfCPMZKrmDD66KUY
gnPKe4slpkadwbeNvRfEwPnaDrwFnKMYzQagzj+iHTasGfz+oMMGQpTDP0GeXPqk1k0uhVoyOjVP
/rUPdxdhyf8XF952Z+kDtFyoWtgjikw4lvvqruiwYs+zTBwxEtGaYS0+oT5dg+ZCuvJ3YxQIt+xX
cbxpsyfTvlXBn3eAiCoZVY9QRv2BxXeDwJwbW4Dvbuu4jw7u2TMtNl+e3r3BSm9opWDluX3Lah9s
MvrxgXr0funk3RnoizGO9yb3VLUxgH3nHWTY2JwsqKBzPerHE8q39kuGR/vqQWomoFaNHloOJmtk
HsXTAxRYU8rSU3hpiaZJkmvubOLjIIwS6KUtXW76ec0WEHkF1ESaizby9HPG50JLdB70RkfSzEqJ
EJHm5zjtERAHHGNkLWragncC6IUh8Nh+D7Us4ipBuh4a4wHFfS8aWktDnqMRq+tHaeihPtnPJ27W
FmpMHXg9/tvRa0MIXFcW1YmJNTCIDqze/s0AySNoVZx0zySlS49uwMicUSzHFPaifwiWkRy5rpfZ
lS5lgCVi45VSgl5CcjlQoiRdZuCEqxIl/ofC0YLk9bn3AgqJ0LJjH6jfwaDzgaaL4P9K083n9MHa
VzqOMmkwgY95ZfwA6Zdk3T6ycq6N4+fM55bodQtW3YS1ciHf3Bax4TzvMWxWY03T2x8gr+OaOGz7
2fz9N277BDW4BruDeS0bojocJqCjLXGze1lB7QIt/XxzFL42umUSwt8GG6AMt9seHd0LtnFEZ51q
Vz57rwhlYDUtBa32WZGLGzd/VTWdinS9YxqNzWQP2J3/LRdXhTr1c/OC09SUKaPvjGz+rQF/fb3q
wfJdp5JUJadd80SX/XuVgcrl9zM03p7Lq7RJRBns2y8uEQo4BDjW+SIh9lpUwfnB5WKFcoxVpmlO
JP6IyB5yClTpboQ2NHbtwa7WbGzNRlP55XAoOj1FRdHidSJTx4O4TK8jCJXaT8+tqBXGPOmvMv1n
KrecEF+QEroMewej+U202o2NWGa8wDbBXsWJaLW83EYO1al6B68ID/piXEemxRrCbhQYwciyjcdZ
Xe61pylHU9JBWx2fKJ9qG7af8YCdhhH4xAekaCLosse+AjiAe83lgKVMQgi9I9h8O9fcN0T38Zla
I8MDSRfAdsGhoCFbpKKBcxEIR3T+1rjRkzTXCXcKFwT3wf/qgSfZRR8oZdpvROgNvfBtknzfx50X
IrCD2W4hG08D4uiV7QggsZbGQlgSFv+77ARvVJ3mux+Jng43V+bLIagcEKReNs4q2m/NYEyD0JMV
fP7ukBd3mKq4jDVrW4SWWpLZ59aQYUj0/gJiqK0vGyjVPtO8rUjbScTS13CrKPi0tBdANyZjDoQZ
ck97/9zk6izXO9ruY2bH1KZIOYp64Wr8esofEgTIHxaXO09CtHfh7aGLPnGpP9GPCl9lJStrQsT8
gOq5l7GmKQTpR8XuOGbPDuT5LWqJMEZkKMH8kzKdi53rcKbPD0Q1KbYf1VkYFp/WlH8Rpefpxymq
+D/aUq786WyKPX8qsCXKGKed5/GvLowLcKksXxQCscs0UeCuXY4HIQgIypcIupXVeeoz0bGXqmaW
Kd7Br6Nk763vgUQMjeWxTxjTrfPyQ/BgtvhNJEYHt1XuvvQCCpnZhzg9sSl+utmYAmHPn5I1vksc
FXLMUujh45TWvsf5GdPLVfzL0Cb49Itqy7NV0qGQK2Ps1rmBgjTBdVC44wfhtFqMHvSEl8DqGXq+
n7vQNrFzJONmLJ4JhQNxqBIs2TV5inwTJ8qLfz/lkDahj3cjlFYZdue/71/4fgJHRX9lz1AocWDW
J7sA8PLPvo0AJek2MYXVqfrplng6yYtrBk5ZBzKkIcauBr80KxtMRYEymTFp8ofCsYAtThELAxam
7hTz72r4Ehjy3BBD1QZShl9XZIJxxN+561trxKS+SwLeZJPHSPN6TJf7nAxK7n1QOgsa+j3h+gdk
319zbetnRRsDX+h7SBI4i7YqJJACkAa53sj/zC1hRYcW7Y+RmOFAUzPm4KS31f6acWA2sWfl3fCG
rXad2CMrB3zFYbZoU4XqOXU+brctzXFZCEhUUXv21VucIbk0uNQs+pNPmNjK47NbU3rLNwT8H5ZF
zJAD/NwD1S56WfIV3/BaUFFpKAPVTmZ6iZnH3IvaWqi/Druf5hB4kL/eqkDNXSAiJKNoVPfOYUYV
eFz8zrwTqrhKHBa9aJu0pGVzSZCiElQEKLGh2abl1w03N0Lkilm96oSW/X31is04pHUQYFUWraqg
XD6LGSSkkG6Ca1WLf7DUvf6dPw3pJbX/9lAmlTRvCfTEWh2kYorrdqGpul43fp0rtjKnVN3L9hFt
db6KeHQ2WvQfTa/G+lDw3mk4VoOL0Ii450n3C5GC6Y7ufWkyFnA45Q1B4gvZH7SI/ByFRdneEWrr
PmCOxdwtUAllfRUSoKXqKg/m5vfJRCDVBKBQQgAbna3EKpXOy8ouZuUPbztkjXN2HJ4uGxtzDn9q
uJChOpD2QmNTbyYKF4cvlnjzyrreeJbb/5YqBz0FgU+kdtCmEAyrk1Aw1Z7hSvWG0MiZScrot6xl
s4GajZHTdfr0nuO5gy7BBw/DSsex9e6Lm2qGODJPI3IHiiZVJarwAlBZl9aUSttlB8hbIGPG7+/D
utnvcK65D7G/SsRx7ULjyiFraMNsWCxBTo9VFlrZtlgRgRJeORzweltUs0qlj6Z2JIbUy8tA7GSZ
cDehR0pBBc9HgWnyN8T0sz+g2HiMtLaWq8K+LHAlZrB0uENi8FjbHS/yEucgzIisAIrHZw28gReP
aJMhBfF/ObHgAPII1P4yhR4Qait7b87N5KqKzRmOqeCueRa578s2bPljmamkOs86slZPx7L56PRL
5MrTbywbsYF0+vaYJoapxJM9QxdpSxpbxJs900rprAD5dDCKCG6/3iTvhyJi8mlF6qjusyCpqEba
SafXGPpQWCSOBIK0BsbGHfcCpeOnMHzBOEGwHW/RMycXAbtFbKdHs81i3w7huyucbdm7m08QjZwj
DSIegZomRClt18MJGhKUPo8u7VEQicjsR47hUM6IYeXZii6tBrEjc/JcQkcbLLV4sy6+p3n26zoK
YPPD7NT6+Nd63jbSx+TVnOINnkJvQsSuucR0PIwxJVwu2Z0VQQe2/8frIq7uRKNGpVNP/3KiUA8l
WmLzHchQfBwEpW/mwCtnepfzOhZRpKcb5XYc4aQOwZXh0xL1a5/3mLgU7UpnMFpD95HrVBfmfGLI
eH8ED0BlIeLZMdbWZWfnvTz6MvjLPI4c9wqTllK583G1/nbrdqwtIlA8B5bO4GTg+p8ANQdYp+lG
H4udWUFsFMOG9kUtDhF+64zH1BJdcFTBWTcqeWQeEnZ7+xwjguucxKSRRQgAO+PS9/eE+JnfHr3N
iVv6c8B2lONdOJCharKmW9y4obE7fQYgHmmE1R2jY3xOjV8y8b5Rhwrq35YjoKUI7ryZuL90aA5D
bdSwgeBy2jsyup7/YHEc7wjFRwshiQpjG3AaC5wonwNAWK4Xt4Opd0pAghamqxHseC/QcE1D+Mxb
6xdqdfDh1syM6HWoqkAMzP4/sHlyXYfUyTOWP9x0OdThcfHReseY4TzaN3srmOF/WMZqF7CWaNzw
yXHldEuRu+OZep83u2ryuFWZwrxQSPMBbIND7y5MHV3imxWmXigK+hgScxoNZ+2dLir8qmGAxlgn
lD40Spaamp1r3GBLde5/H8Jehkxg41eUXXAL9i1muXK85wKN3QFJ3h6TG0XTDSuFDcRBbpMio6aq
uhC5h2KIQAqRTov1jXnpG3AgkU+km3mA1bHe07FClrH8QrNQ0/KQ81lTexu3mSyht0j6FLc/6hF7
ut4DzFHxfX1WL+Mh9FaiQFncQOTeWEURzG3fzYrECZ4MWeTbmjcaa8zau68XziSbQ+tAKE3yoWF5
bcNtj7yGgCPFLSnMUIVv6MjSAxW5oRxq276skGtA0wTAz9dO1wq68pTGC1R1d0fJ7FarLXVEWC3K
JOcvReye624jcwSRZFF139yEkZwve8SpjC1WcCGjqwxeFAfzx+NdFBvdwYc/KmfC7iWHB4bxC6IY
AuIiDaGdNoHe//mW0BGcDBbvKeZvVO9thgAUB1g5Ye1fJyieM3yn/TMMNUMQtfsr/xj5WNe1oZhr
Fi9kqxxxg8Ux8VA8CDAP6XJOXy9rx1hASjgFIn5250AeEPXx36ybK0zf6345zHzlZ8Qv1Uolppq9
V3CqnzHCbvxf499gGnbc6UjBhjNByX5U9gcswtNAwjbH9QHnONnvuOouKp0blAUrQ0oxh83WfPXS
cC/nDWlTVWckYqyAe4c6Gi3uQuqvCYzjll9XnT1KoUnbq+Kw6d1Kcp226gS3aa4cQBPfuhVsMn3D
FoZYYQAfnVkyxrRzD1xYtmTCcOuIj3lmSHJYvfaz1OxWY4Qa83WYaQ3OFSnccka8+cNoXB8SrN41
aS2ii1JaqLOP/YboReH9hSWf/OLssDUzCdGrcs+7mqQrBIjtzw4vik+SxDYpiTgjlSrzGHOUvvxP
blmtID59BDNzXFl/W0jQnJjh6hswDUOhFkzwjzl/ks0VBdgR7n/xTU0peL5ilf21zKEv5aE2G37V
jKKSDnNfUP7FFoyb2hJNmY4cZT2NzRmhoELQ9ZVRnovn3OaVmm4GdsiOcDWR0SiDpTGNWXbFxPgm
xfvea8KHFStd1uaFgfyG8L18Hz6oI6OyjZZoyE+ERkTgG+0mIzVXWSyx+3Azno7UOQlgLqWNYhIV
BEnQ3w5lo9eTwQI3sPHykeQ4ukzNi53nSGZkc48ellwbMo+GkBrIIC0ppvSfhWF8zCZ++HWdad+g
qioiyPS0fZfOsGXCzNNfwYu+L8N3MZCrt18vaWloMGo7YRHr8tdNidXuO32klNLwmdXr/mGkSc97
/yCiuW85vQDzkXr2LFgLjRgwC7Ym1ahYadG26BewGn5zIboLARyxSMe2aVuN+KXFLs4/7RETaQWS
CV1DjNWGGoSIH0xdbzLvocViFx9Nws+sgnkJtuzCKIYALNgYEP2De2gWk+hlnPUpd5WvPmA2X5nB
1tSDpDDh4ntXzJhHkEXbpmgdyW/Sg923526a4XqLrArPJLrtr8Pcbqnoyhrcu5B7osCxNyKuUKv6
zAnj1OHjFlmSIdacLMxHw16EWer+c4b/a4WhZ6xSR33cEaQCPZo12pHUpN21zdZg+sGLS6JkwlKk
qbPyiCoGzMuwIYDqqdVRSlujAEbxWknbq1M9WM48sKIqjwDI15EYpql6qTOaN2Uy5rON8PEYnoZ3
Ksvk+vQtefpsvrEr0iC9OkcD6OSCoV3/DH/AYoCsUfcEpu3Gi6Jv1Ae6GitY4AELhT4Gn+Lnp41m
Bxq0u/KuXjT9vGNfJCtGNDqXZAYr5qZzdwxQyeL5MJ3DlXntpBdeSEycz3g9Eq1ZBp9BgYqkjpfe
zXsA1TdAGHZeB1DDhLZ77KCaGn7tvcpExkdNt8j+dyoTphkQPwwnmzAQqApmbB7ub+NOUwswIXDD
ParihZ1sxSOznrubMGKobc7/e80yGWhpYcmpu5Hk+tHU+uUILAt/FDDmfpchI50uW0Ff5S70S2sy
h8ZhqGVvjNQQuxQF9H0ryMIEt35SGHgwZszrtxLNCAP/zUAhR4HP3MFbwE+sOVlGAvmP3MKx8BSP
voU06u6b6r9REyUNSPdOl4gGOoIWKZJFTiSqkyWbfHtk4y2zWnodSQqV2JNw2ZctbYVLgNY0mg07
5Bwima6ZGDiIIlUvNKbwB5NM5HHOgSGrm/WQJ26YvINIV7xNpGswNskoO8zyBb4Y0+CWqZDPgQ+A
xcJL2qMHZg/Tl/zMd0xNSZ0ZW2vJBGrIKuIi1W0v/Sv8rdmP4QRrlynZHYmDyLpxD/5bFoQp7ItM
It+YdUrNiDuyo3IGW/nUmwzaQM7hugArvjvKB+m58mgI21ynY/tqV2e7D3AbY9ftHKjjHBm1Uviu
RMbhtEepXlNQou7szhu1N85coDvNrKsW+gFEOtoFkFXZbO+PqkZj/2bQFUMHk405/KBx9bHtZEgs
t6KjfpAik+T4OoSPRizWPOsbc6KBTmiQJJYUeXM3mVJNxpfgc0GQsYlIQIYCZhewiYLYWVozWcB/
aedqTsmZBNjnxAEOtCmL7+9wrFdjObonztKb80ELajH6hheek0OiCVM5IbJM8oILI4gzjAYyyv6e
yqCJby5t4ceNr0ykT10P0r6Mu0W07e/lEk/dXnHmtAr5CCtrcA6PfatQjurUBGnwT0Y9dQ9+03PA
PqDO50qla8jRIWirs8BamAg4U/IOtRkKhsRz8k8o5TSnU4dZsQ6Usgezn4Zaior0txkBEBYA6A7g
wsslp/m4hynHD227W4qvo+546DIVh1zH+isn3omW+OwZKlmvnCmOnCFn0quPHyaLWJxvL2fIuF+T
xC/nNb8YCsXd/Ba6VlOgiHKVIMalZ2gzkUpVKRRj9qO9xXbb1w6Blwk0PVZ1cIQCp27PxnvvtYLq
IHLpstqeGCRDHruiv6upDykyD+/tQEOiMvsa8RdxYqv+lNOeyPkubofjVdK3xxJx28YtSoRA14oh
uf3yyqPzX/rHcNPTDwEXwSLkQ9Kj5wG7XdT28oZnBeGCTZBv0fDCqGuA2omgNNtLAZhUp4/5YkPR
qBjA06yn5g9gvAbok3mx0gzaUYN44PjxVGEX1l+YZOg/nLHzlHo8X8l1tGCtqpqjQeMJ7iQKSrFW
vGW7ye7PgW9pkzfWYPrxESapnJT+mHHToqIRNZhCXiZJVFOyVfBZZffDFRxUmSpkhq4GjQ/Xsb9c
Jnmw0myLEMxe5GRbsjtFLKEoXRK3q6SfUMt0AJ3l4LBgPa0tfEQiozRSQ56DF8FZR34lOgPmJQVh
eT2v0nt1KGBoO+asWPzfPYy7brtoO/lpQvZ96MV2fTv5Oh5MAfIwz9wqp7REtWPtFj7SFjnU+fH5
nmH30iOcwk4dIJAtawUjeLi4RhTreHfyFs3hU/+Gzh61fgg5Loe78OGuIs1AM7Sm5d5EgtNRf6DA
syN0WOYQrADusBl7KDzGXdhtD7ZBy5JH/99u0hHD4+IO1gAbJLRC5jtKNngqktWLapOT7aSvGMFi
Q+iZcTRtccUKUrE89JjHTw8qVf52YGaBuJvvqlDh1IxrPrsQIVW4QbWLBO+3G39SF28eniWLhaHi
2fvQm+607PM+iFMd7rF9UFcQ/FTZJswCggXmDBr/vnHGoxkZBdV0aKsSV+4N1r+/1ayRMApZ92fI
0VHNJ9LC1XzMRhU/Hm7+ChE+D5CR2qgpnRwPSjxN5xFNr7EEIZwTN2Uhd1ut6JgGrFCHQdTIDl7u
jAv7ZjOs/EycYjRpKz+1RbjkH6qRkAiQCos+AvWq9T8umbkrEPM6PLAJIIk8kKQLGghxL/HMDOUd
cT3l1Hxr+x+RQMuKbI4q/1MMrUH6o0WIZBbJVMA5aBvTk23ZRarTwbuQpnkRTep5tLMGXeMiTJVZ
BaCSJ3TbqrDRI8FISsW0IVNw4oRbWwpYuBfEgPivbl7Wx7YmcpfLsR+Cto4pXsjXxcuVw08ETYFa
bsT6GbtdOxjkgPwpJOK5xqVcx5wku97yN+sZ/yb8jXCETpkaUfQZyD5iH7rpLV56YcJ3K/A6h5ki
1mIQc16+03uKNC8J/qkmv4fTBktauUYqrZUGAg0M+BVG/ZGjlUGxyn22WiZUFnsgqym314mpUs4v
ALc1TRloAzQ/JO4IiZjpH/UUnN8TQixX49+RAu5lA3MZOZDk/puyB9a4iSdhiq0WzQrQYo1+dX5r
uuv3daxUeiry7kRXeisX/jPtA/LjqcO93YGeRZknGTQA/rj3yH5kfdqZwO7DdmMeL+96KSZijhS6
ATDjtBptDvv89F8K1J+2YaJBaQtym7R5WKuMcmsM1eT+gcj5agI0hd1kikFtP+PJL4tIhY0Fz9g4
8Mur1E8qW9+pAd86DpEGO6PN4WGIF+jK5Y4n/eSH5jZT9g1lmzbtfPSI5nVKgYXpB3Rlbzcvz9IA
HXU0WsvBWO893FU8NTblNCmZduAPw7l2BhACUJ6k3UfzBhAwAjItdikqs/Xr8pDWwIPQbcEDINS0
m/HGdgAdNjqhf73OfOzZKHrLVrfySlnNszRHLIMQe3qSkdPbh0t5pGp8Z2uve5XhFPCTsv10ms/G
kDciXF93Fbq0gpBCTK3iBOzbHkPYEqTiIzVrUsJTGekj19ADnCh20PhnzMnYlliaAV+4riTGeR8w
6Io30KoebwcLodMV4PN0cn1fSVsR16jP0d1LbuIpQjWKDkQpS0WiGqkUONJWn88coCN1UMyhYnd0
typRFMpCq/kJ/GcJb/XZgsQW41LjHNjPBi40fo5hhaKeJ+dEK02ECu1sCqAL3cVoocH6iz0liFK0
0ybF/Jz3yk8PpESSg0YIJZOexTYHPNZljQKu2+NpHnDmiJbNzf5RdkGxJ0nflW2sjSPSO2RKQT69
Z+D2HzFMefX7EqxNu4tv/RTPtKdGb5Su+aPCB1haGYpb8VwaPq7WR4yitTPA7uAXvHuxDmbPax73
1yDnpS27xS9cnpsfc7JeuqdEKA0fcDzqVuajqrWynTE+02yp1YEpVb2xFD9mJZwlAZX6CQj0nZgj
7Esj7EQY4KqB5X20nw+dzI1T0rWRSFxMC4m8WbmSNAVRORZiWySGPMrGFGrBdxIw4EGaibmO0VcZ
CPPcOVkEOvqW1Orszi26gc05ELyDOEzwtzY5bvqLuJErxOeQ2oy/Ky2kozTnhluvpQmON8aid2TS
c4YxvZBFDNembSGFh1wMorc9QFSvHaANNwjYpdcv4N6RfeAwOnRaHQhgRSYKBpbgbVZ3w0dxuIhR
UpjuGp88gOzXAAqG4/p/7L2FmWqECV3prJ1PM1tb3cPQNTR0V9Ev9Bo0vrOzbGevyajwKCC1GIXL
KIadwv5URmerRKGDtsBkO3PfWjgeiaiAcFpQlUJ3McKhMk2yBSKnMzyym+nKRXr5eDGF6Iq/1UvB
EkeBTqKUji1l+DazU/Ja2f6O3i3UZpFhE/QpPLh/LtDlDd2UR7Rb8yoUtk4D9sUOyWnXnuNp276T
N3Kqe/rMLaj9DcoJ2UHHK6a3Ifmy1qiU26n3OC5qqtb1+VyTsVcqLJfv343hlpwZsnsFZCN7b6LY
78fEJ7unUxUvTiI+pIWuqcrTCS7lmFDU5hFtGwFd9RMjB4KNlns7PNucLQcSmaG+iY9xUtk3GsKp
XBAm7IZ5b0rO02WolsdBt77ysjNT8K8HMCPgPlZGvavQPeH1TDiqPyu/xuSvrc1ra+tOtknYVJsS
hNe6kneTuRRZBg/6CByfb9p+6+/dNLvB7b2cVZwiKB6XzA8IgFFL2DnjGtL2EcZShEacwHwxkSDT
0BUACoek/VDIB4548NcQMCUtWMqKot1OsFgxPvyI2QxzqbJj3sxcchBbnVB+fQ0MCiXrnpVtEYGh
khXlx6SAavDfl2F1IiVjsY44Svx2cwSlopufH50urEQjC2WMA5xdmYl0rnSRSn8l2RtR8vvTg4+s
wE/BFZDFdd3Xwojoy7w0HJD9N72GksqgUMzhgclV/NJORyBBHfUnW8AqhXn1+Pr5L3D0dAMIEbIv
ShJvIHEqubwU90k1vOykex0jEnhvd1On3PW1OMvCkPWf9tT/AhXjgHbhHMrLeJds611H/UmOSfSk
gMSznuPEQiracsOhisZg/OdylwGTwr9GH0WlCh4NZaLfRYFEpM5L04MxAcZlNSmNrGUBCy0mW5N7
e5ax1Z3/zr6nX/Bzn5eUw2nmqP7FNP+H2nhckJkaqLZciNcVSPFAPtUnLy2f/FjE+op/zZPGRrOm
4eDX/87S8+HeKw3xaJTMTGNqzZwPygyG5d4cGydAEt88G4Dpc1YpP3ChQAmHPNkJ+GVoCgyHQdNW
60EICes9QdAtcJwiQcBBTFHQHiIme/8EH8EwPZANSmBSU7SMMUpL/w6tcFwtOxyRN/O9M5D2hAMC
ctVyWjEGbrnjYhV4PKj4gOGWJkz6VSpWJ7PyXowyy9Ic5Eag7vN6ny93+GkYEk7Qz93ubLSjJTOm
nW4CF0Q21iGKjoVzPvKL3ID69l518AtqusV8n3uKPwaPyUnqGA2/qmo7z1yJ6b+aGs3O9gr1SP9k
75Ucf0iCqxw0YFSRtbniYv+jNZvi9xjh+Nk00307jRhcpdYxCOXclkr2RZjpDBHq0fZD5K7ttxfj
uuVZd4OcSwfGh7r939DEQbL/Vrp7KXFT1ekI5tWqjNzrBVk3cGYRFEe1r2dzJquYWHGpSgLDp+KC
hMx5Qr0yInCP9LB0O0dt6eKQ9njaPFeJ/YDVsEaTzaQNGFcX0j0nzxCuar3PiiLPey7ON/f1nrmL
E8CU3Pc1vcQv3SaTcOwYzSpMUKn3A0yo2TzTJ1wcb/EE4NThHWC98UbNR9t66wh2NTx2Z0NJ24tX
PaoI8DEXWvVFplLVwNahExT2iWeQMdnIA9MSIIP745I6uT+GDPSIas+8qBntRCRyjw96j2jt6zvn
cbeM/DMYRlMetnYhEAmeatNN2tISBHZowS5NElMWAhDHFZFdjFfxxyh+vpa+Wg9qqXGe2yB0F1nj
bPLmspFc92IizX7U+gnF1PjJA+GTHmOiDd8ufa0V9CvteundqdC1i/aamnY0VawUN3GoBpch+txn
z+tw4mli6fMOTL5amLiQMkdUNBvGYTLwNb0dUGheJOnK7HvTuuzoov8+T68Xyw2LARhlYYzIzJzc
k5W3vLPrbhVYloI9dM56LJrPzxKw4yQk4SrnRFg5Jt9AeWH34l35SFYMRDwefX4zk6GMeDXbSGKQ
82UHOyC5A6d7uYOba42MTd4q+fJtutxPcyfOwPfc3R2sGgA+/B06g19LEQ2L5mQIzUJBgdTZEmwU
rX58tHMSuk5kZVcMYXg7IXTb6CywbS7smymXhIZWTO1QnWUWfqhvhgxjZj1Zo+ghLGdeqCWOcWzp
oQNB3pjJ8LYYes5vj4x+pDyiddcRq7chT9K1xnGZVYUU4jIcpZFy9LXj0eQVFVaBtonXkwXZVUsA
nHadW9MYLXbkoQyezwB7M6vFjCWjd2EyYNA70IDGRnUPjI6+nYTSoV54tpctB1CkVE1RDTlD4J+M
7X1GgR+IqgRC5n4k7SL76/X+v+hvrYurDFNOqk7kKU4Pm2KeOqukzMAN5wh7y7/x5xe83fEqkx+5
chtepkoETb+agZhbTst4v0FEIPdK3J2sGxrG/gh/l1yC9UN1e4ntoIhkzLP0rr0TQAaAMSom/w4+
0aTyc1hNIf4VWN0qyfvXTg7p1pH1YtNNL7tOq65569YSt5xXuUXntpOR7RPDyCnGW0YqSla3qhLw
DiP6QBIyahTVSx+cVGg+gORn0ho3JxrAklkvC6veIYtesNhN9cDgVC60wIRI/jjQE6UCEMoF2ubl
wjCb03GL68d9knGn2fnG4JUBziXWKA71QXTkYXi40JJbJXwyqW6vyIAizDrq4bpuD8/z/+tQinDv
lnJUCPxsDHj7Pp7fKugckxgqr0dYKtq2ub71AztEyBErcGAoyeQB1VjPnI7ftzH5yZ9PWgIWdT0R
3OawWXNyPfh3OcD/vpPDaapn4EElQdrltlcw/vNQseZviXu2D99oai+zU9H8Kzjhh9d74x6irBR8
nYAq+OjPVmQHqAfPKS4lTYah4xaQC9We1HJFdxLKdAdgnELYd3cwU5ex26OFJ0v6VSXs1fi0QMhX
s70wjypwdcW6JUPrjm1uDTXAN3anwD9UhMuAcQlk69qZGd9R+jQyljYny3gVjgFHeoWFF0wdxxBe
Ep/jRp5PwrOzoJPZfuoat/5rpIyYpBJbd4Qwdb3rXNsFBJZU+NGXtuJ+Byr6ioFDZb3uHB3tk5my
w+JoSZxviF4xoZyj2lk717J+IJljfvXlzpQsL/EeKk0i7UPZMyuDs7hwdO5hQ6H9+psUodGCItUF
aezLJBnW0i1vrpiowJFOvgNaErN5J3J7l/gOsC5kV7f1gFcdkLPvp67GSgY7FHXywBTrZ9YjcJew
EG5Eg62vAD28umb63PBpF+O3nvyHT+ZneR+GJ6scyjGsrT9CAI4eVQd4T1WRQxIuY21lfzKTGnrF
HeFDB1MzmEKKEqjoB4FkqJ5GadDUFiU6lUKvJLPryjtEGaLFMAyhTYFHnJKiAbsxuzPiukhJcEK3
sh1ktPnyRc19bedt3zNpVqzotseAuTu86RmvS4iQl+qaMdKHyjHC+kmr0aM/o6gLIZA+N+RPKGzB
vpDVovewa4r1ALGKa0qjRV2xTP9yMmK4zWKGwFA9HalbZXRyBzRi+IlDHCQhCuu8AXd7pWLY9a96
I0SsFMyWHr4XexaQgJUJK5CALcv7EbQx5jbsSMQcecx4nEi8ZDnSleN0tDccX+A7YZlMom+LSmSW
Hbbaui3fWOq08RqrkbjqY5DJ7kX9iPNu9Vq+TURdLGpQ+UTb9TAvf1+uBR+qiVMN0qO4ZzSdT1Pp
BefTMUw0G8pq76hyC8MmTsHOXr5LgowEkgqMDoODDQ24bL7p6w5MPM2jpmbl8tL5IvHryJM96lXb
whzUCuU+edAMp0HmHLRXnTPIckzyWiBnmIRAL7L/Jy2fO74Q8x46SSGhGX+564smkNM0yJ66Gpwt
FqT6mkLtuBXsPHcdblVOinwMtm79QySYwa4EOyC0TujLLF1JCe7BvlIp3CI/+gK9QIS2RnaykUui
Jj+jVr1LCVrFvV8U8/wEL9VU4eIiQY5eBQQ1E2vMd3vevHEl/X73J1F4mA4HfyARz/blHhbYoy92
fisrrNxa2KfQ9LUl+op9iQvsC9De4LgZv8WTFA5hVUyqWZMIfVtO12GL1D5rADzgI8LC7VkZZB9x
KbHUyQxGizNUaoS6AK4bBB5CPJ+UyrunuLmHI7s71WLAE/cscPwiy6woemDiJmDEyzBUSFHN/Z9E
hscTpx3lwq/qep98vYRkgDdAW3g0jdE+Y9j/HdLupNGWiJ8ZGsPorE37/Y4fvSj2GfSfXUscXFBD
FkHkr7r9WN+Zw9TLnHXzBwWZYqmeVRz9V05L5/3KdtqRdRfgu4ZUim3JAD0TJNs2FWw4/OBSRtIY
9QD2EpRbTaP7BK4j9ivIWdKbe/amYcP5PAPRoDrfsrkBwhkYEIrD64TmDb+408bVR8hccR2HVKTD
tO4SZvlgks6fxqEnzu51pqCFLv4HFzmdhG5QCjR4ggZU3+WJRafjLyrW9PCaLFSsWdH6Wozqm6OR
+LPf6wkJLAg+bP18sWUZcEWODviH9kutmV2kUKN1DrFezQqaVt+wjrohnN4uRh7KDcuEX9Lr+xsP
4xkDPoG07St6quYD7m64XwaPdNhO3m/6dyvc9ZAGkwK6OqVQOba1bB9+pnVtkhOocvFsV/OlBU/m
xfnHznvgE9dOUQxoP0v0tZuMtv3wSJ1HNmq4HubhteBMflWWWL+tCqPVFpIlP2IwcuFTk5CYdoaS
y97QSRfed1tSsmHPeTdFycCQvby6pMUa1gkSds94MEY8WnMm56PXSZtHj+PMS4FgbVoOp/0M39L+
eWZuj7lz+yqgTSzKTYmwfEeQG4TGSAeo/TJggXxiUbH0t9eMEwXJ/0IKH8nujo7id2cn7y4yXWV6
Wn5MdW+VlbVHqpDSMINhSjCoKS0IsntjQty92zpMr/ZoyJWvjNggQKXKZvxQ489eN8Uwsjdua9ns
YxC+HZCvSPj9UR/ImsAmT4bhmPw3aQL7+W3VKw9xfuHQ6msv4x/UNrY7npewgrTNjPDXJOYtznbf
biGm9bxmke1G2DR7AKM26SbRjtVgzRDDJDP1gWlC1ZlW4OBcVcQHM72VDF+62Y/jFbjuYYjhQ0jO
sBn+8ePooBsJAT46ExkW8Zv5UUjulqDAyP+P82YDFgRmL3Sgru/urFPeU/ps68HjqMKhiGq6jXb+
BLMC5RExwq1xzHAk88iebK0pLWj+qK6dn5pnILbxcxc83rqI83fgGztaWrmEWnBLMwtXvFshqUcO
FBLQ83iIKPDN7Z9B3t3HsnqRjq0wm0+5MWGEo4IXKN0UJd4UGgNrzE1+8Shzct5RSo6CHGbP7Vrj
xSBQRdkRfgB1jcT900I5ZoSV/yy1RcDWKKAWPaiCthfb60mFfVEXQtTqZYizWSeg7uVXMuXZOO4Q
uOQ+eCQdY/QgaVmFAqDtq1Wrt21W4tVOtGcGCgEKnPwrCyUq0BW2M5UhP7LNdXRa8rPGj6YvKZcf
gFCI/HNBry7ci1cp6JOilxV0NSvA5uLT115sc+cOJ4LCMKXNR+ptI/eGXpWb/hCKhNEBuTbqy/Aw
EcSVohNZVrQ5tKoUEpICe2o0Uv+ViV5gxdTOqZ/KdsHxoZGkixLnpMTdKERCGZiZQricc5wZjSi8
toAy7+NzQB1dUJGtYPGdRgq3akGNZI6EUMmZ1XGhNz58euc4oVjgmv1xBxyMvL8GjY38twUKCHn3
uFlDaa7wXBdm3z7N5eCrKYlOtJnSP1GRoyQ8sSl+IQMo6Qj9n3Ay/ZsgcRnE2MNuxWV1uk9URM+W
dMjDKZHyrXZXcUVSWw0e9hKwLYwQk2YTO7Dto+HEwlLM+4MhVH0nV4UJRZm0GFyZnFr4MnZ67l0U
1LyLxAky2fvSSZ4QNVZcOKD9pwqXygUnwK1s08HE68Ir0GUGY538I9gWuL7kKAI3Eq+WOLP8hNvl
Tpbu9F8qzB9RifFS0cCqrwGDQKCLZO8aXqNUmVeiMFdoQ6ST8Vq7fDug6WOoz3L8EtyA7uvl3GXg
AE8jDUpHQ7ytv0do2pgK3fs731FWhajfaaFxABCthU3HCCnEhJN2mxTOdgMGOcsNW96Js/5GPF9O
1SalCct3e4uCR8jiVjmNgcGd5SUXwijYYBSe05/bK8+Ono3ze5U4et8Ps6lBzFA9X1WljWm2sYyx
mwNbaJXNjPb2BHczsFwdMeqAmEVMnQl31nuOJPs1+ZSr4NIWG7c4MQAahIEK/ZoxUHemL6nZZXEs
XziYUtPPXAi/OhK+tw5MPnKF7fjKpf7fzDkT8kneUwhmC3BxJ4PStYRHF4o7DNJtixHXrh2BUDT0
NkoV4uMie18+9Ob6QHuzEHXin8jOZu1eAHN/j/yOoIeFbhp3ykq8zIL2JmysEagQe2ENRu6k2dEL
zo+8FHlc9WGDFQdm2JhzvNaGyWjo7DneM9dfapNZhW21NJ2a0qe5lmtWqhGVbYdZlEF0aILsrmOu
vHr1fO74CHGAnCiO9/SjU4tm5jxrzgN3c6iMI2k7I4rrsK7bRBOsQM+zIos2oB8dF3KG0oEVB3/a
dRlYLm5Ss6CkBIv8W823wknapc4RHSNo9LcSTGQe6mbqbTf4L5Raj0RAkIPWbuhmKVKgnYUXeXi+
IlNBZ/OFhef0gCHfMP2uo/23dfaWnz4erS/5aHQezamuMzgkPQuYTMvvQS0Ao8XJmj9Q9bTf6jpm
FPzmbTERfYBZsPXBJjEUUEIWi9MPTbQZ4d7SH7R0iXv+FdeQQukAHSCGaOXeZ/fKaS8oLRtYZ+ut
kXviLGdZCfM2wuvKiOTLLirmkJ9I9kJfSG4cTvM8Bpnw8sxuJtyVkJHrx+pEkRIsBn5ju+1JXNRn
hAJU7IIJQzsywS/C2uLWuC0lHLdga+QEb67Wp2JfkkPOEEYHZHWfLzAg1BSwSATIlySanH0gopVW
w2SknMX/9EtbAP1O+g54t2YK2dlkZe55TKyrS1UoJATGW2oVxb3aG/Aq4KDlwhIrEeiJd9Z8hSeX
ty2hmbOVJwxrsdqUgoYAWe+i5+mmjhRY/xdiSs64IyZyWE+G31GXR/HaTq0NxwWTcjNz7Zba92sh
4Ct2ah5KwDpAfn7puBYEuLt3ukZ2KE8UceCHajN0OuuEZc+AIzAxjGoMArU8CxaBucDcw1wtIW2i
31kuRMLnaqE9/WMyALy0/wVA05NiUy61nyw8I2bROCVv8XwSRVOMrTUDafqnN4peza7WQFP7EcXk
pGrsqCxpBdmWCNzqBe01+c/KM3/kbOCKV/2kMtM9IVsoy7+vBc28pdxdQ+n62VU08dgOhJ4P4f5F
Xo7CFaHa0eMnDN9sgpP8tcOlg16TW0EFOgKyXOz9bfttiTXaE31MWcQQ7BdhFuwVXk4n81Ozu2ly
eKkNxRV5l8TH4mN3ySnU4rkHvaR9cihjJCjq/kow3U+CPQ6ZAfpOUz2jqPw04J6Ayu54+x8PiaQ8
WaySX/jKZPPRmHsGG7RWtq5jeFwzSmo53rB3JzGgbA//1QY8OlBpiJ6FmCG/bxWtRNZsZBrXeSIw
p2qEpwa6baYEEbnUWXM4bed1uPWNl7YyxKkFyfLRnZg3OU16VFEZgGWrwTjeZ5gBz6WFJhaTG3gj
ewT6gQReQqWCph7FP/cuqQxsjP2dfJYqCzTY1YOrk+yZgyo67X5v9hszDhWu/Vo+GH9KmBIt8lRB
w75hD2cMmrlstBnQk/baAwrGJSiQaZD9QbGDR490nD6qeHtPAvcqtKl5oCEkQDudoArWnirNvQ9E
hI06TG94NHI7PSNV16tMkgF+Iunw3NzvOhAXr2JrmRUntWdMdqkJKMYbnyNmBH90dHjmtP3FDHeX
98nAU1fXy5hgf4Go59NlLfD4K9i1PqDQIUlGILzUGqNtBr+x0wd3W4Ivs3WZvStMSp2+p92MMKOA
FuzxWKWQDf4lgu07oRNGaFOAm6uim3MamHL6e+VcRUB+nD0DZ8psFmObJEMIrMDAzhPni8RzZ3HD
yy49dQfJL3SzdL3AMUHFSyVNxe91YJWxLrbnW+SMH5XhCruCAz1RIHKFKycGhkAKKJTPrwDvTvC7
Gbdh4ixnm3XyK1nxytudY2YoT/gUoD+H2LNYnwMeSMmIwkSn8EX8PdUjn/lrmXmouqm3RGrH6owd
b6lHy/W1s6dAFjcqSUnTW2VKOKc0V0uly8Bhbfgb4RHQJvM3COiEBZGQmINmir0RPPSC0JOctyak
nO17S2C+IWMM39fWM+3LyQhJNo0vtqJJS/AaMa66o3YRnIDi173Q0pIfeKG2KtLYFgt/iOyWt9H+
N0fCG/LpT5MqarHmgY44SlEwfPKoqWmB9Rlmh2fugaWmgGLL080BEjuKEkgznnabync603haBfU6
qotTP5PSVX5WETHDx2zgT70zw//UqsU+RieMeg6C/rEBlzJKK0j/g2Vv1kImAGwzWM+MTvwIsfRZ
TOU261T3pJtjZe0BL38PxYiJS2p8Yv0IF7I23C4PopXBIIwCZNAtLaD12daX5T4HS5aYTmA/mYlz
WRicO3vpZVeIYXv5a13Gp91d+spF9uV4V2zO6FLblRI8C2IcdOiS94xuVlQCHjfc6sflA7ERGPkR
7cHjhQ+i5hugu+FlMhtbS9WfIRYm8J/+Nq5bS5/uCPrxYDv/HY+QOLv/Y9rTEjUGLCABl8ujIG8Z
82gaDay43EPSG1JULvNLxl2EIs2PobMmPyy6t+zAjh1e+Qz9YgG2Gt/GVRIFTILBgzTNzfzv9MxK
kEwL/xDGbS1qzSMjry8jaN8SYEJ99psUaHe1C156gXRa4Bsip/pxaq176Pzs7j8vrZeA+EQHvnhs
Y1VIFwDM6Gd18pnDBzRbExkxK261g9o3+5PH01bi4xAy4uAIFmfc0uvKj9eTTbOMUKZevKCuZMCD
8cds2LF1t0t1WX8DOApJnMVuzHutGF88ITby8Be0BeY2VVPBjpEOEh0OhwQ0NK+EKJYWW+Hly3Jl
xgnKGP/RFi2q7aXZeYAbO5XE57HJPShRuYjBwf5k5tPvee2x2wceWICoH8bXVAwB86Fk2dlsdyks
pTCXVj0m4MdDbZV9sg6rlEQT2Qc4Wvl/INbD7mRyqg7b20jDFlIgBf6Fsl4KmRmLVQNHQgQAEQas
bP7u5p8OK0FNQaoSnxv8KZ7h8B1LYyj5MhNgFihtCCpvVjtSsgVSIOl59mgpWpeBUQVO3TDX4qqx
T097JSbdyX1HRpUz4jqkn8C89rm0Z6c27mQZKAcooSuhJDqGVpxGoBgU9Gcz3xRvWSyjVdlrSc8L
SGWBeRfxtSyk0anN9uWPfDRJkEr9oEkFIO0R6KJHTSNS9Tt+bioqIcW4aiQjJZ5ppMgIydA3BcmF
waJ+zAznH56Wt9WiqD5B/NiyLw2OadbNehpMc8vbN6KRIVFAC5y0OF2YApHidik3AAqwRFDAF8c7
+7SutGE9I/HU1UvoOmKWaD+G2U6P/M1QYDtYNPwfwxWO994rfXrwQt0i4zOgAo3DlLGDTTdBWqPT
I/xY7isSC8XJQtRWEjMgF+IGm0iqRP0R7RKqHBGUDu1CVWp+P4I0JIz+txmnNFniix1xjqiKPKOd
I7BhCRIpDW0VrofJV23m7/o0jSCcPHohXpeUsH1J7bP2AutbbB+8ge0VCw6P8pOMnGtmhS3edQKR
yyy6Q/t95/I6IPAZXZ0vQhvRlX9sxifpohvho0jer+cHoWxfCVn8t8fpaFUQ0yztlNlmQHCjyzLb
IHP2CMFPTsHWYPsHLKOH9piXgxIepZe3EC4vrve+ffTJrhXbeYI0PnCbKJsN/HNat4jYDRDZmNlN
yfoFydnwsg9gPAsLExjl2NvGSK+N+RmMuf2bU61yKwSa9PHfiGt0Q7TIq2cN/7LMzUv80oxwolw6
aYpq0TwYmnb4ipZjtLOWk49IUaXbzVD/VeNJtwmB8XINn8auEAbi67nxiaxnUv0RGzo2oP3oCv7l
qtX7N5g2M+EUej+lECjhzhkLjFgvocGmmd/6B/MnLA4zyAtxVTSH72fudoS4Y2rVgF6PgpCbhMdV
ptouCep4Y1DtsGUPxrixFYHNFJIIxDDyGWDQDIKxfjALY/YsSpHcEOJq7NIkc63vNzYCyngeL06U
2Tp2IdnWXKBM1ELDIk4x91Ci+uCSHFaKh9G9hjtmzybfuzYS4KRt0GOHvtVf3Jm/g6o+EuYaApnd
FQkqW9wrw7ZlwdaGs1Zwh5MCES4qmY5dUCmcqk5s3sLBuCOx0Z3dtRKpZW1gjpDamtAZPzjhdEt3
koKESd7fE27kXStokHbyQKeAbj8gOga29JutjNKGDnl+cYGUaXaz/n/argI6yaR4KwRM8Jo8msCU
opLG8cqeTkeK0O9saJLLJSMpPTSxy5vlHU59m0W7Bc74sZbT8qIfHzKN++Hr/3R2+Gce4670rmU8
a8UEdmy4TcfKNeG1QAaWGMtwfFtAqTLsPmFVc29fdc4okn//v9qWAqw8DG7k81G1LtG+OCbTev5y
JaJ66vHbQkmX+vbj26vPyXiSoxr7aGf49gUx2h2C8KxOy2kmt4n2Os5xQduqmFMGKJ0vsBtWGyus
+4YRfRMac/SRNvLGwSf6i+4U4o570WzEkVE2FnK1cepjvO+Bh2392dx/0iYhWKT5WBUyAhiACxcw
Vcjj9sHJ1Wxz1UISKJy9YDXFVTO5jXbQ9srP99+t41FbuIUTpAxEzb89xjxbQmr6YY2xF5Dzxhqc
tsHj29/d1xFp8qW2mUEm3JGziIN2UW6gqK3+wO8vLqmiqgNdODtl4Y1SKDWbd+tNOfHU6qGVXM/a
5CfIM9e5BhCNr/iBkKY+g2rHIT2tCBu2f6dc8PpBnlby2afk8oVfNkD+uq+0bHEmRT6WRXsRF9tR
2UPpW2ApqpGqV74HEdJKO/Wro22t92g+jcyKn85SXhVxB8tBEvddRusrxuD1FRXigyauUhSVWq6i
mM8VueloBBBzwSpiicc0JWhVVeKUeAM+4Hyk586u632sEl2Ir2Q0DzGGHbRHY0RFFOKQMKU4aH6z
aYFu/+GSAoEk+YXIpkxRcNpNThlo7L2UJtd7Q2fj9qmlv7O466G2tUAKyO/BidE7ZmEdtyrctm2j
y81bltgNqCF/wwljfsQhVFvKKwNje6xiTit65DY7vLnkVCA47lIQi0XGWT1YNhWOZjg8c5UwhA7W
PE26wlv+XfCuKCRHIMxFeOe6uNnWw0mD4LIwvgl7VrDadEz8jVMK8w9SoONmIVc99EetRBCH+15T
BaLsoyrpHXPzSEfdLFCw56lTC/7qSTbuxLQHeFMhyUoEAz6kchAYJ1EOQR3lIYYHP6XdkMqmSoOw
BAjRVyNo5dNi4zgSXJsov67u+tmb8tnifvm0/cXMWDHJIMogYeU+qZbxr5KavjpusyUCwTEEp52c
aQjFAmnzKhEKPGkUiXbyQJhvbtYBq1fQd2tBPZWge8l85mC65NKup/vKM9wQRGV4PeWUYwrYde+F
+UqjUtNMqGb2PgoeuRrQ6DW/XLOl+WAZaYHkSNNeCRDOksm8RhoSJVJS1OkkgQZC/u04M33ZjV1z
BPg5SYfszbA5te6FxFfvHi2vVjCoJbG/1upi+aISrnIgBQ+6CzuCYc8aJcTzGdyW4p6C8N/ktKPn
jhsQzNrnR6sJCQ2ykKtjanDsoszNyl6wgZ3a7EI5nCyM+KAzOPq6N7B0eXf5wuaoqoPLQnOnjHNL
xYhYYx6Fc0exUPxjIyMvYaQEuCNW9p0ZUiiZBJijcJrhOqg5mGaQ7nV+V7U9SxvHxwN34vTr+6dr
VDXIHaEg/92kXU+CkbBKF0KDmUmsf/N5f4Jc+Y9XtAFI+S/IN9FeW/y6ZmCWgfq9BowMNyATalOB
Lp1SKeGXJPrFoD2g0U2q1iqrOXAaeu+1pB4BdD0Z0BNShJWjsHokvA/CMe8dX8cGwCaprZnofxDO
ZAl4cVcMvY/FzGxyQz+9ZS/98JvIgDD2jTMvEC1PNaqRe4DiQ8N7oa7WJJnclz3pvxelpMyvW8YD
CCVjpn6a9zh9MvHWs53bYMS2Q6Q5ZkzY29lOwdj8u8lyI/fpujyEPXgPRVVuZVomsgpwzGwHEL75
fBDJA/x3oSSSEb/YYdaQZFX3IOvJ7F1ApQS8eckBfa0OtdOqw4VB9Vypaz33ZHQM6PA7LW8W2lml
88SrDt1FkXMsHGTGosXDR48u/+/9R3rGBmDSDpAvJ4CJ1/qO5Xxlbhaas7I5Z3kHXVrqU+HuID+J
Co+eAlubuScSFwNq/hGPuGWX02OAZ+rwh05GR50CjbLRz61Ks0Pd4phSBCq2RL8OfKmiq6TW2ya2
2Fw4Z0T+BlSvE16MZMSbOCQPE4yQ6kELqaPkuvw7WK+oBOwwnzs285HArrt8aWFERCp6S/wgMYca
RIJmRFD7uZLpY8d06IL4ZsyJhrea5TKg6xqCzVGi+LK8yjczXW7pZoAeYAZJzzgM02eqgEt3hab5
+j+dtBgIc+nMf3247EvqnSQs5puXy2Ton56iMxqFgpKKH831RA4HNMCtOzp7mAkA56GG3NdYEP2j
Wh2SMW9zozkIgc7Gb1yuRiim1hZ8O/96wb68QMBbCui9+dTiK56NfxGZZuKiclE5JHENqBxGsCLt
LVOVp9cU7FScnbw47U4rnJYG7nKN/DcaFP02lZtJEtUeyAoGR3edT0uYzykkqxxp8b/U6dOcgQBL
xtyCTYbph3cUdnuxslSPVDEDEbTQRS4gl9OUUMhkmqitIRUGTPw3SkUlXEZi4hNgZa9rMl8+uJ8w
ZjsSUyA1xHyaYoJF1qIiW5NKnH7bxNxiHeAbrFMrBJcltzKJw/dsB88OsloPci7ygIoGfD++QDGd
jJ3qm2pyGOriHuIGQJwQep+ZElgUiGrWCsi7HBUPrq8Z+2en6UcJkZY4tfCkxjyQUIUxVpWlD9el
NU+AUmz39by33XYWGjefRDE+TX69WnUkVua1KALmMtD1m5525NwU+uTGzRSxkOYAW47e2PHIkdKA
hEmICabdmwmInjUcdjc8gnUFH7gFRDCYrkq4VXtLqfxAGcb6MtilGbGuZJQqTMAu9r5Aqs/X8vxC
QOuCwDYVNN7QtvyokCX9Q1UIRBLSgMkflgjBTmwW6I1sIGICDLh1vPCH5x5QARfULm8d8Ggskq/z
uABqzPuwdsuLx56izgE1EmPlOq51qFSb/AM/zWGYuzglyZL6J3IxWO87fsLcOjdblMMLkgzxKAMM
0k2V7zd6G9uHspSBGXhV1GAMwWW+p4hf8AQAfoSvbjd1p7yIJ5aJIdwpl1bLwxsdJf8P/k3PXk+7
wYLpeZ3hV9sgRy4SW4EMiVIJ5nYgpFOlyIzageaGmVzW9SMpnk/T4FDxo6XYbJRsv5Uwt87hZlYE
yMvWR0TospDRx6n+f1dDlxKWesX1PSnoQCjIJ8JxRtGwziCo5bQd4ZWM6UdkMXw4TGTWnZoVB0vL
0nqDpuW2XWBRCuSAygmrlQfmwPzToHFQ73ZM430Z0XTMlIvKxpLbuGT/CEoTVzWBRYtYa/D3u36C
ffJD8CKmm/axkSKXb0x/EHhMiS/MuT60mFhgXikzUWV3WJASbvNUEJit4v7+u4d48jqGYOAFP3tF
QSxf6ZegWvcfnw8auhVPkUMoGyp4/xIubfJeE4YEqkp5BdP7Ez5n5+zx+AbYT7Xcwg+oF/VkW8/D
IOMHF23XGS7so77qdprq7qh6dwEY5M9KXzs8RE5buxnYmzzOZFTxHpH8BlC7+nl6/2RzI0Gh4FJ4
t80KutVzKEAJ/FPwFpowQ5RBFR1hcfluMkSAGzzCLpz0sK+M71UJQiljnRXScqgDVV7saTT2K6NU
6KcQp+V8ZQmC9DrN67vveX6S3bzJv2a6UK03uHUYU705qXUVLS+BC+o8LSgetTe2H+NR7E5/8Q7h
yEcMKUJkQXl13uH7jLzzSIXh1UTMC99sGaaiaGC8QeR0RVvPbneXagY3zFG6DxIxSrVDTvwhjKgi
UGtL2IthUDTQc9zJGYnBs/H4rBkGc9svprZsWaRjhabZ4EO7EyA/YKu7pupSkzTvvwQ6F5uHlIJp
bCYHKWXQ+ArbNXDlQAoq3CcGIZH1n630ySBcW2aC5au3qksi7vSodTH9RiRCoMqCp2jy15H+PpIi
0bnlNAjpqS2rFe9TMHVCF40IRIMIrQe4txf7li7yqIUPIJ7KKQIRQ6WUH3UlKhg/OJQonM2h15V6
Bk5A1VuvYA87aL0GUk8uC+lTT/V4KwZU8MpQ//ZGLHTR9CG+mg83TQ0NWrWcgmYTnsAef1mTXmls
aTX7qBCUmYqeQaorAlfdDrB1Zq+7uZ1UpCawsgxd2xcC+N9H7wTq8xyj2IWINJFEtQt4iS/YXECr
tzvBSd5zaPnwxjqI5KaxhyVl21X+orgQbdn2A41vWcfUvXmBbSs07JWsKhvOehL8AoiFaN1JSGa6
FFMyskZ2f5zeytqaqc8rJN9kJ6LUTlT7ZWB5gTJuo7tnNaVRnb7MPrr5JRU5R/ZjSD09M+N6+Ix+
tbw/xgx1EOju1aV+cuVu+0yxhY1VxGdREqrAy8gmtVgS+1GHgIhXH09hJEJqG0PrSY+5VsiW89LD
ghtas3vq+clYujsyELbXr5Wv+cx/9zWOlee/VvrrychO8CudWZLuROsJsaRmZvz5F7uDBoAPiphO
suTmuvCJQTpMB9N3u8PIKEZiBnDzBZHHMa1GOzdPNjV+XKitD/6jwvc6zchoRzYK5h7PFjFzR8Wk
8yJdDUMEjvVwWbewjjpxI8qUfHYD/V+woNuX6dYT0pIPoQPHSN5os/aTtzzL5Fb9Z0mIqEHgJqgS
w2CzAwtg/ZNoQwICU2ItvZAUdsG0KDrSlp0zXwbMFmOaDwHYPz+pYJoEFTTiQ6gDvQDConmdczmv
gyN+OpaUbgZyqLXnwc/+hdVdUXhs6m2b65ExqtH13kBijY6J3y8eIwgskwXSlCb5sD+T5on7pZXv
9OIl4k1CDVd19OvIl75LiKU4vHUAX1ZtjvxICWmeztaSPyhsShXt4wUQVI0epM/GjC5vV779qgoQ
L8RIamzK2rKNRnCZJWJiymDYM5mX3L1+b67npoHJpnYywfYBIo2rKr0CLdAhDIgtnOehvlcxJpAE
UlDD4Q935snA3Wxfs/Nb2QoophpJr2qPWhRQlVrsQB0nv5wjXRe4BdTqqSAFqzQfHT37Z/CZSYRF
fIgt6txfO981mQyRzQdUfyGTIRk5dr1AluA6v/biQMvmVGKBWuba4SspDm8E7XFFHWkJA7syb6zg
rdoxUm1H4p2S4iWv8nNTPUx3LQRntoL7oIyKn2O4UJzPFFZyXtTbxTnxfn1WHqu4fcjMHh8CKRqz
OCJsx3z98oGU+LiFrHGETl4SvQpuS9+gN0uDTHsb3SIxDAfPbiotIN/44rZ3aVfYAoFV7E6ZsLeN
XuXhFKlfqxQ3W+1tiQ9+/k43e/NBU6B7z4K8IX31gJYg3lWzTmmQPCeBx7uA2DrBDnyc0AhmhYTF
KFEt5WUW5jvqiqUeYmkv50foiB697qwN1cuUjM02ZPcZU/chIKM6CafYXioSQzecnZhTWVQprQmG
5EY7pG6Dnv/awJoTXYYU6VgFKAXQkOAV6gTDyry3BZhtnjt9havvwncBJpXrD59ULXbtg7PYxety
pFHKfj2PiucQ40jwVvqcHFdFNXMkuSS7L6DUTqXgBXKtGdDTsNPEin+AIUvmIaz3ClQQ5eS/SUKy
KJEQrAFEYmBILoh1GbPnsUrmalok8Md5o+z8LWE6wuzWHYqpTu9HRIsh2syvy+2FddiWo0xfEBnN
+OhZFHrljR1mI13Vbwix+rb6wyDTBRLYtIaFUfXqLc5yfJzlVLsYnajnXenCHpysgCyIb4qhsgfz
h8ACi1lcZBwLnGZ9qsUeNBEFzCmzVVxLOAmXNH9hYrYCyNlFd+dlq7A9N9z1y34AbtLAN5NImagN
YtV4YpjZNM30tgdBOZ1HZdrgIAbUm8KbFUX+gMC8g78Sy45XSGIQBgN2/bKfadLa52osnmpdkFg/
IvjucNG7ekeFRAbnZaHXpK6099FKPWWjWNUBeVBldwIzJzm0akS7Ls0wgzvh2iYualnKsfoPPd1f
r5oLMQHcKfJK84yZIDkYEJyXvHWOdPtg/L2c+6WQm5T2Akq6i+wp39ZoihLctgzNSDMVbsxVpxx/
6DUYLW1gpl1a79i3XaEFhu2s8dFKK7MenqmgwsXk7MNFrezoPPic96OgCjr25us72Go8hLwX94sz
346rbYmzvai2IJ13fSFp4XNNFbYZOk2REFy37v8KrWponuhS5/3OkTz3hTw4X67vvRlkIF8d3AZa
xk8bZvJaEnBj4H1mxAnnTrpViOdjiCJDlOwXDemgmdtYwMzfRikK1fejl1WtOV6XNvfLGLktDT54
EY/It6Bip8q55aE5Xm/dp6zOQD5CAPIXFhTAjJ8g5g+OsHjXOSRcgVtnaNuacKOo2QShIqSMqQ+6
Pbb2UdyXgsxOXY7MUh+Q3lUXQrvcc0h1Zhr+A2qhu+Yvt6pGEqO777OQQyl/AWhZ1ik2WOdQpXE8
ukt+4pyFFzWd7O/Nlk2aDkYv/DXZuCRNavvK7Wpz4qR3sblaxAtGHCZ4tvZwzO9Bfngh4Fxa4ISU
GXHCrs1iZj6zEOGu8+XbhF678MjE3/BnJDPXxvhZr1C/TKTcLkq41gc3PKVQQReneJI6Da/zne+u
CVC3uShEAQmJpSw8Rz4fqgfz8/yfxj6OJ3vlqdNO+rCLLlh7oIjgdcC13M0GRGyOjAu8kMQXb6HM
sg6z9xBvEcOjPK7/Rs9g1vPvO2qJYiRLA5FKI8wBe6thuU7dcPdXi7OikGN3gRETqp5ZlM9m44Jd
R5DQB2sjLtuTQZJ4IFJ3mj6+F7eThpZ7J1tF2AROBVZjEg18ihDWu9wMyjiG8mB4TfnqfMyZ9mjJ
I1ap21E2HMokWzcjxwirXuzBvO69AHrEwU78IqVCeoNLcuR61SYp+8VIOOJpgQ3dQQ7dPYLyjWdl
Kvq0ruc5eWoylQCKBVKeFFG3+++Q/HTNBZjrhSXGxWv3z14s4y7Dtb7bY7pSHg0AA4DRiSbBVB30
UmLtf+DOmubG82oljAc53qwZ66KWr6hvFfgrrliGTK+Kg+0vyO5YcHGiMe4k45ucK2QXw91kIMhI
o6Zv2bIw4azGHT06NzIkwwLF8VETJA5PN+rAzJMCxu1d3qlurnWKV9v45oCigcEwq+DJCZ434hJ1
tv6J8ex0I/SLWugMcmpoQR7tU/a7ZVgtNbFPyPcTIkVmbXWJx6cfHRF1oImbzZ9jgGLZGHoKQxhm
BcRk65FJ2KiL/feMsDmnniBhLKKFS0vD8w/ls/9tL5BsUncnyZwSHSMeSGa5kVfophdqLRroelkW
4f6RSeSx8piuP/T66HwJC4Uz3BZNgzKTgdvseGNASBAYqadpNV++L0w/tbUfuXj+NuQiSvwCDS2+
F6I/tdrALtl+pocJTUdUEMgNfSI8LL3BoTxSRZgw8zp4Hm1UYXYo0184z263FRZPlNoYbddapO9h
MKE5K64XuJleki4SXMvwtG+ab31ou94PUA2oYP33Pooi2Nl57zG7+/CXg5fSz2sA7qCKeDDbecGx
WjjQwCGi2lXEJpv0SPWFJwHfsYHr7D1c2/g8yf92Gi1rt+ejV833uFPpf4crXVogItYlujzQqCsA
uavFt2X9mLABB479yYYAvgL0I2G2FtjchKP0Uh01WTSuvSZN5kfJ6sFW1TMAR0bw5KuCI6g+W2WD
Os9+RuPNT54kCKRPbtXD4LRjo7pfMQg3FTT/lbTPZk4v4aGtH6TH9ERtRLm6BDUwULw0W+zl5Fty
l8H/mRn5g9Z7tP56QMdSsxa/1XKrH4G7hum3p+WnV5CyUJZcDOZw1gu2hCmrZ+IOp9c5Xy91VJTg
gXbN0QbEv+Vxjj0BGhosP2fMKCl3dQxurdX3/vNOcXMAzN3NrTfigE6tlkxrHjarnURbP6cNDrsu
F4OZCpHxgai0JKz5KrdL6AwkVq0JGJDD7xS2CvIuZjeSvIvGbdYgu3KfpkEuT6H6+3mqMSN+MNDD
5CzGqBJNyOvFFlaD6owvx6HozJd/+FcOA5MziO/NeIEUO+3C57qvTCJvwPZUMh8Jlc9mvjA2GH3I
47rlZ26xEB7DtHv4HoU6zBI5cqgCyBqJXAxqCA4s58DSsdQ5+Vo15vlYjR656uzFeqWD7UXo2tBG
mWJj9Pa9bBI4ARbsnDE5MgxiN5upuQ2cI5cekG972la+dAACjg+islsafITcdSpW7ENHPFcT3HDz
srEo4Tf5ENDvmztEOeNilCxep2KmlxTtPXeOrN6LXD1YqNLGPfftGV8Fi+YUM/HlwP9xF37Y8rTP
Oc+dyc/Qu+Uom4ad29ZJmpliGCaeyX1feyHwsQfl0+cPlZMFQafYEknmx8A5eS0nfoHVdvID3xTl
nJ71mJooH08TE4BARpD5OS6V5fHGB7zFdjDvOEt86E14Ay93Hymi5Fgo6Hdg6Dt1LCji6gikXdNR
Uok1BbCNTAq0O4ORWfau4q0Z6+8Xvv2mvQDbiExNzR4jn2rdtBROaetCwX900qBDQtI4ari/8syz
qx/+PMXa3PvQirVsNkGoDJJ3IIp2IorOUlAWWq2EuVYYcsDUMBus8D1ntYu3GlQQJSUac5s5zKu7
SNrkrBo5Ijv87pa4UhtaWdc9mAJeTX7GLcAAN33iYQ1FZ0mn4BbZcLyOQ8P5/QtXf49uFuzJ3xS+
24UGde54NWWRwy83yE34ejg1R72VX2lTLl04xdk5bu76ARCLWAiqrYP8BmgjLP64ZMhrIHQpKR0n
maOs0iMWkJO9EuHEFkxLLshK/nQGWkIQqAsiUdwOtFlJGI+e1x+jPSNXVqaPzfYXNbBWyueV1+zy
ak/5oYcEzGoE4LGXIf8gESVqHXfMIA5Duz9aS8TI8vKprbHOLm3DUv53rXnz2HLTbWqvjYk1vCwz
fRr/UTZWBT4joM9Cj4LS8imM1cZ3upUPJHziFccI+j0cimS+m7IB3ej58rESSySa2yVlCIscLLoZ
KZdFym/Beo43paUE9FZGYACKNQo8sUSE7Ye6oLxWFv7SRDn/zba27k0pF+DKgnapizlUkVBN6sob
ptxCBijpzGWGIOeGrYLRwI8RrjAEg5H2YoVmd78JbRL4uaSWd6/pXoUIV5JzY6RLjKHmwDRemqC9
u+ujJq5+2x0ko1hCmlUvNGvp7G7w9kbDsICKI25GydLwIAQr778qam2m16VnjNnavLnMvA3pQeID
my79CjVzRjgWVdK3CTTj9YIANoZtUPqX26uIp1evSgMHAiE1TS4VV66Cf8vErw+JPfeczLpFV9rB
+XFMC20oS2Mvh9bEVsGmCsIZ8Sp7z0j2SEjVtjH1MSHV7y8Zw2PjGvSo1dLYnjZ7KyIra6KqtgO6
ByZja33IPS+l7JCak9RXYzJmaBlc3d2d1WZrRBIM09SHd/0PeJ3vW3tEfLYOSU6Uj7CWOKUr8PZ/
q70sZbg/oGw2S1vpxU3ClrIhV5xf36P7ygeduAArpJX/tzrfK/2RqbwYXImkGxF5WDUMSp5YlOlv
WTi+f/AV/5uFTTYTBJwFl/98WhuZKbMAb/9Tjq/hNhuGUttGBHkxCkJ2c48iZ1H6/GOBQYoOJ88c
cr289vJuRM2z2ekTxK+gikMh0cfI9aUfEkWcnPXeyQcppVNcHXmb3gKgAQQuxuVto4rb1mD9QTRp
nrGWJU/UtyvH5PcQNeUutbAhKXKlBdjVu9XhgX3PPGq+54jJfm3w5eEicBULPgdK5qrzE8XFBMUN
NpoRTvbiXfaXPeyX/UQSPZK0CG+5NdPI5PqoFas6ZPzR92SQPBj1iDBMDR40rR99736KqVl2faf3
+j+xTBS9GM67x/jQ+stVRRIuIyWVb0J8jLE7YG39P3x8OB13sWYPTAgdLW22pc2hfhPLUJUJXBf8
4vXaMWvpruTOPmvv+nS8MuzV5amqHPPxU32e4l9YZpMZN1QtiVtQnDkVuSWzGIXezLEuRLMRB92/
jVXc4gtC2PJxiIzaRjp1D2+bAK40Q+/aKvfaR/MjgyPKqZ7eJldFyI3RNxgcUXe3qMD0yrytWb14
qAJKP9X3t55RaUPbz/pHKIEVgCKS3ZgRtexN/94oc7D6tSHwX5hCv5VjOh9ymLu6dcuItUTiHMjm
DNk59dRJFiUTVLiFy2/Wwez//EqdZNNhVFfWuvEmXPSxJx3iZKqpeoj3hwCX84bh7cAJHnt07mKJ
Ti+Di0iiDwIE6xw86L2PSXySSpx1rljTfkR/kEUp8IT3cigLvoH4Eijg/ElV6uCv1Greo1k9UX7c
YsGhVvMoi0ca6yr38Ux/HeSW0Bk7xT5HsTWdxdozqEi8rOzU+6KQdTcSXqwIj+hgzhLcALuObkjE
omuuYWkFxMYRMm/ESgtGGOCh4QLZvs0LuusHQ7zTm2QIZ23tn5oXmFMPTxb6gf0/YZ7FfjVJ6AQU
NbnhLQk89p/2GJyN3LYUjKkoHHcoEJqlMICJg+PZCboYfcNmYw1qsnwpLwanpdl59624cQTB8ZgJ
HH0QYjYMiJR0h1EtXY7XG5Xg0yNwUxm0Tj3udg+oaUS3BiOl8wcheP3naI3QjhFQ1XrWzwkDly7K
UHpTauRLrqM9MiWCdPpCkINquZTJ5tvgFmL/Y5vvQGlGbpjB0Ou4A5iTAXvLEgfyXoUS90akpIjN
FSYYYWsHwnXp+r2UK5qIscg3VX+4+zqG1x+bsvhu99TXDPnu3VpGAw37kpyFCBNLgMR3AuBRS6gv
9PbRW71hpjbrvMSTNrCSvozt3Lg5Mt8aZTd3vPyUU31/AzSxC7us/PMl+7wcDUMD5bA94i3PhMV2
y563P47qgR+RfKWTzkBlZ5ZYvXHnPso1+RnWzuidTanjA88mKaT+D75GHSWTPiKxdBPu1r/h/myO
i4hCeatwdjRKE8IbTZFomttyuSiJawGeyqTNPO0ZnpH+lt1jqvvl8qXXnbM05x8PD2Wd9yrUqRGJ
mtauAqkQ4h/OesR63ZXmuFxE8VMtmNeBByRV95wxaJvX05dOcskgdRpzp0WXKrO4VQX5wpgNRBwc
K0Opb8eXMNf8GtgBjd5+stPcPCvXFt5ldB7wt60LxkebqZx/HS3afXkFa69LzhHIv5vCEOnFgm+1
F1D15jOsW5ZvDjFuVezJ5FCuD0xJEWpcQXB7DTgKhTDIeJQ7DoyA6Mh4W+WE3x5O3zC4tMNfprM/
n4OlpmDUUIn1A6Dhnr7czQ8YnXpqHU7q+/rra7yAgge8waISB6iiPOvah9pRFYvzi38+V2kNYXWA
+Dz0BW7cCT28Xqq9aUycBfFsxm+Oe3sQ1jEZYs63Xv09Yvdc0XwHAFgqPmXERsjgd3A21wQCv9HD
NI3tBInsNuZ33vWey9qqFaJaBi3lSsQ1YLleatx+LE55PIpmgP0WGDZH0ERrxFb4ZRetiTB9rGx+
frIdY8+2x7Hx4vij544HrguhIu/Vbyz5JSuIK0LZGYbMytOus8cupOa9vlzhFC16HtOGmqFUdBv3
nTrkJhnjaWQIVU3zysrX4NFto84AIT0PGAN/X6Kvh5lY0YAwJ9PAZabtxc9nAOoYtX1zGNJcaspN
Y/jUNlXyPIPjwKpE2RXOhCojyHm/oaq09iD/DzSL9MQt9qmDhkaePVmTBLSnBLh1rxCezKNfYtg2
YDMNUGuQQRtTBeAiHBA6DZGp+X3n5JGFXFh0CAX8YpVBW5dRUVqv1+pbfBtEGmVUVwO3TiVpC/Lc
6yWkL3r0UW7V3yZdPUmazlqdrmZsaNxT3IIKzixcSjJEJPcP8XyMuFE4NigqSY3kY2PacvKFLQ7g
VU14Ak5LPRHl4ary1C+Wl/ST0/vysFykTv0Ario/ixhTeBKQomipnPeF85FgZcZhmwJvFQP0gJe2
ARsBiUy9LMck3rsIBv0MD4l0etpK+oSPkdicUOp4qx7f8au5UYL5ahifyWbz9Yy74uzSu+WpwY1g
W2wz5i/EOhHK28W2FFhvB6nvWEdYjAp13POySfleED28EzUomCvXSVPSw1H57krIkEWPapuCOMCv
mJKZq8b0x6adnl2cZLHV0Wk7NiRZNytmBBEUy3SAkxtLv6pCnvHrGp1XYMJQgpTdapQaY75gZoAG
uNJbFnEh9NW/2Px5T0uvC7rwBAkoJDEr3+KWGTO4Ygb3G2i3GyIwo8kHKe2U86Ceva1U8ITEhYtW
0bFWXdew6OaitCe1in9yHwdvu2y+nYxMq0roLaC1bxoHAq7SvlGM5l86mP9txj8ap8unHh1kR6l0
KDGjsJDsoUEmQ6jwJUGcMIyNp9W4JzPEDwhlaT+tWRUsdwGgkmgOtJkA4X+RW/UpgrQG6BgOSrOT
ExHH0JADQFhjoMOZEVGSQs8QD8QPm+8l0SwI7gpZgZGB0HagH/56my0lLP53shE8Y0fqXLersBby
UCXw53V92BQiVrrfmGOwDRtmaqYLX8rMRfBirR4SF0FwgoH67iE0ejwL40E7AGnMeRACIwnATTXT
9SvwZ4euiV2gA01WsRDfiA96AedGdcGjbcKgi2YQLl3Puga689+d2iNgJVCDVmmAoejqt45wkD4w
fgDWadCwUAXJfgGpvjRTDeb0Fo5+irKxR68biDMo0ePJ7xv+iSZskziFtBhiOmPgy92EF/awIXx4
K3iWMo/SV7o54oo/CMJ0//dYIu6MFLk5SSJ2gGGJgvMABQ9gXmtW5HcUuGGFLzsAeyLkXI/1KwtK
ZrZ/r1813JNQumbzJi2aPbYxRU1WeB9jm8weySEM65KKGAek9qjNvNqXLUixROudymtcnUTYsxlS
px8QQPEMd8pvlXm/Fc1M5pu0y158IZ1tOgsKc8FsX+Jeb6PEO/d38kpPn19abG8+2C5q3JyYUd5c
wchGO6jWK3N5qneRDNEULx/v0V951R8qEfNUDzGX0F5+fKBqoiTzvrGq2vt3UFtIZGFMjSaqpXFc
aSS7cIhf+jNyFUiVeFvKTn6g+i5PM7ZprhPjZgsDMNpwnvoXJes5HJa6M0QUEEmXR9AiusvLn3Wv
4PDh6FjOGZY2+aFFA6kplKKRZNlA/I4SmwU76n9PXe8HzLyOvHDwUVUgiYxQetA+SbJcgUROkDvf
ofRSyk/hqVTiuSVfO6CRdeuva/6q2w7gzgkzjz1pC/psHuVUUOszHVLoNNOCL5U1ZKZdPUCa5bPF
60WqgHrq5VSujWhAksu2J2EHxm4zVOcK8JqzQ2d1ZwJ9UdkcgUzEBI++fs5O47xahJLB0GXIh4h2
ekJ4i1niIjeGivMVk5UOfTgkezeYAndNO+jiD+7OXzyxR6mXFXOrehCGkW58GyTfCJhfhBu88iik
/ie3cG5geqtwIQbHMJHKJ/MbA7wO272P4+6uPVg20ucNmQPwd+dzrEAWazQy6kTuJFGGNUTuJ47H
ErWRpgC1UmeQrefM4CiPE7uCltb0pPA3lcmB2H75LkNShjmOVLF7IWXlURShvzVXkbJQUerHj9n7
Zh6DCV+g6226SMll/7ZA+6MqMOuFTXQBSIt8ZuCbsJRKrPoiL5FvDBL4syY0iMdRKB4CPAAJ24cG
rnZpYVCwF2VFcATt4TpVnWehzxeWU+ZFUQJlPfNRkxBvfdmkVtcLLmsrhqpWYMo/MuXFnI3zFaKo
GFmDXjoBKndpK/fsMtuJNo408J5ZJaMX8BzRdpoNN1d29S8+tNlIAxOU6hbI+UG2Ij58B6Z6OPW6
DcTL8xPne/+d733GDBtGTquN+hOlNAfIx4PevK4PCETvcmNAObTm655X8v7KgILmriephuRc5J4r
QNLAygSVlnmH8SGRxKv7Pz33FzeaqnPiJTBY7qFnIGlX2qy43IXxB0XRb7Z+c2MP6bFwTV30UxLd
OoDryyvDkBFS5bIe7/HZHOLblxHftO4yJf96XP2mVun5F33nzHP8YPNcm5XiRF3iiDfquH/WJbIZ
f4tXtmHAMcdEhB8+bf3Wl6UZlZwgl/cyOvrBCQaF1QeXhAfaBMQnKvDHNlH3q2MUg5FNfC7pTBFM
3YaoPq4EK2Lponlx2cUnZvBt8LsfJtmK4q93HKTcEAVWRhUViIkge08qHrLNzvmW96Qk2HtsR4hJ
pFTH/K2yByHoNTIGRJLG0flRR3UMqzZRf2ed2KFGpVgEk0xAal/QqsyIlhpyxmlXgeJ6yBMPjALK
ZzBq0caJBcq8BHp2a7q+d36JsQuDorCvqz3fSVuHlQn1LnEDvThwTC1jSek58vlUPeFRKSLWn9jo
8iudnQO6PmOArIe9PaWLvRdv8SfXPo4+idRj+X9/e+X0cQaX4dYaIQniWGJaAI97lQNlbDiJJbhr
EVWWaSDtRNsSFBtbxhJXpjeKXwsmfvxFig/LEBqTZEKyPElisAvRgAn8TJZi46bZpo/v6ufbggX0
A59U4DQ3zY0Y0Sa9YeL4Q+FAUbqCZY/7HYvOiPLZzdXBl/K7a0Nf+elRoc1gk+ekB5GSIoImn5Ho
CnsJjbkSADPYYZF9dJM38FkdHJruvQZSp/eRPRleHYdL2McOenG4HFkNunSbyAcsZuXVHneHTjGu
pCw3ZIAKrZRQQyPOEhsutfZlBukRRChjnAlvKHMOredkWVyoCIW6ZwV6+ZQUBLH2lRkcAvFYzTFm
4InRdduCKMmkTR+BpXCdS0A9/okBtpFzIOOf8Y/TIE9FJm18fn0e2MfjUUQiEApoc/yTrAJw5TCy
PE+7D2mk+x3OBirsHLol3c+9hW+bp+GycwOgzIR1SO1UDjCCOl3O0vDKwTpiawQC94V+y2qsssV4
oBanJbc08EaWX21UGC4XcllngDTXNzY4vxvyK20t/qa5v1QO7yKMrsm0U8O5vJ2nUmZv/ss7dmyO
7iSdQ1hKiKPWTq4otFlswnhFl1Qfdh+bDk4g91B8U0E3E37DxpR8TVElIIVASEVwYH4otSsW1QWh
J8IEe3hSPp4KYZNUeQZKK4s1ffEuqFW7jHCMOi7lDLUENM8+j5RSEYHT9A8BDCWG/bwKGzwMzQDh
LjBVQMb3w6ofRv7VyPQQiNOxJq+YmZJerHMwOwfUhKN/X5LP0MUX4ECsg1Uh27fTjzQFs5dVeQBw
Rg6S6SYOZahTkaaKSCTsLFs6RiA+/PGPSXRJSsno6VkvxOEwNy+BmkqinBDlb31UfzGQySiTK/9Y
HRlo7HLceCvINZAzJlS8dfByzucdUg2D0ljEjeokTQx6NiMZtQpaKfsnrLzroQQ/l+rZOggpPktC
feR7foV4B+wmzG4fcKoH9Row2yZlpJ9ZyO6CVjo1OHj4qZwZigp/U2w104D5JijJm2UkVKblCN9Y
BL0RhVFb9NJWnwoU0HTS68K9k7V8gqhXCOeQdK+wZ1y5t2GKAWQPltjASVimHPnawgdsEcoVl+jP
8Mgmx/4PNao0sK1ulGiyq0zsLN0XfDhPSFiFCwdzWEmvbJdxm8vWLvgXTzQShwsPggUxfcpPxVnj
XWTgMsvRZX/9S6cgN3OCR4mmp6Jpyzzx9JDlKXQq1hGb+2iJlSrZxRidXjRP3run+t6TBn73r7BW
qeQ3Tx+naUDDXAseS2h14k53elna6J3/uqDFZQUrZs2Wia/AcPa4jowKjKMPqaMzWlbRdNL2T/7M
eQiTt2+HZPZckkK7WaBa38s3aJgYfUi4OVWjNh6BQs5qLuPh9z1P+gxbT5hV1ohiPF12wkBqSl6o
3lcxxa+Qogz/GHdSZKD3pnA/k4BRwcESmZUvbkBaUpgJN3Ze4Gt0qlEkJjBwbIyqMeNKF3JMUXc6
skvemWxBCe8bwAxizfar9RbsBCtEl5nTBfqfurWyDpI1JSRkeCfmO74m7CFybJ8K+CqBHXZAjhsP
4viC0OrfPMNf1LbPv9U1f+tEhuRbJopSu27IkVfYyJHEIvbCUB/RrbhYmOk+fg0vrrJUcdofI/J7
9SaSHpxuL9/AUOlRYy/vQU796TwUf/cxrU24MNjfZUGuRWTbAIPSVCeM750LPEjpQ9G4UAsQejJM
q5DGne6+vARnD5h6zcoaRJZxm97u0OsW8pGCwtdizpDY57qMBHsfA2n7KmH0cSt2T37lB1h/pO1+
fIwiutLtUqksPsan8z/XjvfKos6/tgobY1otDPr95w7UkjpG5yzPSKC6FRlpsHdstq20RQEPQ0CP
fdpE7AiC8DuzROMrySO58Ymk8JrRqDSzaekYY7f74jRRAkHdYZNUHDUKcvXG4VgqW1IDH7n1B6+5
PpIdMYKtf0/TEkUes1zWB+/5H/5nQMj39N07K9BGbRqoPQ149c6Y/0oEAeb0FV6dr+IKetNd103W
j55/LrQuXPD6AsjuDljT3u/BlPA+Rvq1SOxAsyl2HUFjExxlqa0dM6A/tzbWIsUoleicB8wZzq21
rMAoc8JzJ5SmStUYq5l984djhRdv+q2oOGTqaOgMXku9KiphiZNNAZXO/NAjcU7hgo9m1mQq547S
tH3oCbZcKh3z4DdB7MblYyKmgl3HIgEviQEKpKq5j3TMT0qGtXvX6eW7smfQBCCN9G4HL3e+Chgm
yZ+PRup5TKcgedYqWzKPCskBtJwCU5tF/9pFqgdsSHrnYbytHwJ82qSxcYMl4PhX2QHPKNIa/wPx
2lTOS+Qy68CiehFYde9rx/yAcACqY6g5eLVNKTwBG4CA6g/MIY8ARqpyCqhqiJ0MWwdUSWu8z80N
mlwSH8sxccSs7XAkCQeXCrWuT538vQJbyOkePbXqUcx2YIpEfs1UvOiwhy6PWP/oDr0CmREnx5W5
ombve66jVKPSITQhZ8oxaLm+eUBU6yokQebrI/O4nlppExeH+mTaGAuE6rZxDWgf9Y40iiwf8kDz
aSJTJChWKhzPG72aAfdP8xarlHm3TfW2+gAwkZalLmB3HRh7rMFRKkqs7hLlqJJ8HMxIXAkQS1QH
3LuFHVV2w9BUQ7Nf5xbZFwXDQh6QfNzDpAyWd8O5A7oyOqhb/tFYZmfA9yGB0IaLLmztEMLTpLTQ
oGgqshS6VHM+xsDGaODQX6I7Vm8r/RGS0Tog7rCiDiTlbKBEq4FEuttpgQvhJ0kSpbAPtVMPrO9U
gcue89sQrl/7idUfuGElCYaiyucaHLdRit2X3JVedId6d7mJ9S7qizKAszKUPPq5HZcjL9sk4zM3
z5Wdfh/ugebTyH20Xu6lQHqJprWhwyIsgem8N8K16xBUn2ekSRnekNPVzoaH/e0A5w/uAGKdIzdk
QDJmVjzkE0MLmIgH5EqlYgGSbsfkzYiZclplQGvZP5qrufYkXxE2rP7IzbOp5q0YRoPKdDZCbTGr
B53Qc5rkFvaCDTeF79UD6o7O6rYt7W1F9gPFp6eGcJIMoHpdxdDGlLVb3UI8S3KfMlerOxYqhVgg
t8t6xCvMFXRQm+G7H4bzROikfEACA2CxQroicYU/tNSAKVoqTfG2Xuji8IZ0FQd//Por7VHrqfpW
GkCm1mCdfAfMHYDcb20Ze+Hxusm03z2Aol+9Vt1oRL3Qi+UyBEnTOxxlq+WO0v5wllYeMaDvKCJt
sG0rgnWGzX4BVeGRvt0e83NjgdTdl0qfkw5h6C0+1cFJojYi0leDgNp7setMVAWOP/4Ue9Ig3Ggb
Ltr9tQkD+A0Twb3fsU09Q/VzD2cGcVrISi+YV37Wkik1hbn6vsO3wjTEFyJRULGzA3AiwNOwS2/5
Gbh8Rl8p61/N5z1pj4uXicHde+g/NlHRN248Won+sgpxztVNuPAyMqT5gqwx/yNVO9/LLfq4ZfLX
jdLXFRtM+wLHi6vavbkylyHMl/r941rjwR6HtFJJ0PygclEd1PO+vzwAMzji1fp9wQATZie4M8Ol
ZlFgCd7o2tZvjM1T5VejtBtyj483xeHQM8SJbkAbtD2IQvrfgSTonN49rzAAyuofJpz8mdEKJWJB
3VAZLq4xUtXT6+5216pDlYAulmSn84zgxh7L2D6dYKqO+zV4XOhjLc/q6SDgVmQJBTfzEmY4kiuI
mxtaNQUQyaX1xo5R0UCWOH0LY8bispbtCp+cNg7rlJUHUPpm25SACo117XO9sdtVOWcZyli17GCY
o1z4Iw/pMgAyAcGl3WRlVpm2fLnM5aQsJdsO3pQ7xEroKwlhX45hr55A4uXUmj7+NfGD/zXV6MSB
+T+IPT3cxLzH7BY1nwE/vWjCyQQmGgM0cPmujO0OPtU70z2zdOFOepQc0taNOV8VaO0cqCCQp8tx
BIMWLXzN57H+De8a6I0lvIwsKnZCiCp7BCQED86m1W3vLvbShJsAREkW52zcVhFbHuI3ThB6luy3
aK/Bhrg2w26h2gFNK7b+3bMUB4Wc6Sx/mnEt/MF1hjb7KarI8DxrhSC2+7iO+l3eAgadatyDMOXF
XCvmfM9lK40/nlH8Ev+Y+fvWn/1VGnbV3bhO7b9jM+nmPUhBUeCrpiUETfih09Ym5fkeKjrsxeWT
SEfXdDP9NtFCuNN1HJvD+zJoMPp00sEZJtfu8hI26RYkoq/rANqiS/gs4KuajbcTH+8iQHIc0TqH
4wukCvrj7SUyKneaDLArXIf+8p99Gkuqjz9IfVHF23QLRJHWYav73RLYce2DMu81umbwCZi/+t2Z
mayEaiyMx6y4hzXLhbhDihUHwQy9cNGmJfCk1AQUpylY5GV/NUNhCTmWuIrSWnYxQJzfPHzbISIh
JFrQPVubpAE0jvS0ojn5/j8YaCYiDr6RQzMObS1meYRQvJADRPZ5LScG8nsnFfwVNnxbC8T+E2fH
FSWemklmXM4rq450o+cVXCp6cjoUVhFB0ehIifbPd561sDKIBkS/1vn9IcTMywYBEpuFIBnhdBY6
oc/oKXmEoMteYu8p6XK12BIhn3p8emJMIv1q2BeAgfm5jgl2hAcWIToicHeYq7TMexOJYH6MvW8G
I3vYCkBKEzL0DdwmpgNxjAt/0QP+p7NL7kAFzQ5xbnfko/QghmOo/OgTGi9x5AD76z/qCnkD8m1i
oxZw1tDgyGNx9ZggXBL97D1Mn6W7eoN57K89SRh7gD4jrRtZee9O0Mfboj7gwqMIVZzyuz1ljwcS
nI+p2WG7GUplPFbuDUmQN+R3rXLKhaxqQegYYW7HKoSkp1kTJdaxRL4/3rwOhjHtFaDy07JhscM/
Bkc98kje47EW1h7Q6M/JFG8aYFBdaeCEulMslEtyd4DXekuC8X+MuqnmQMqIcG6nYSjzhw4eQjyw
nl/xnYOZAwSxOHsZJxw9y1sHEMRnypCMh7ZRar/G7Hr5kQMSbV73FWXB1RZG+FGCDaWbj2Nx2adQ
CPUrraW/7od2iOR4B1s2dZUv2pEwX7RW48zRm0bULEW2jL1lMqUfHMxjDpjCDPwPillbCsShKsfu
hTroYsm2h6HrDgSH3JcfJ/XnS05MdNTCyHrUDVI3k7VQxt+P7Nr+2YKv7NG2e+M2U8tm2M3qvi1n
GvtCrpJX4Z9NFDO8y7a9eZ6rj4A0+fUUiEoG1CLeTyYrCTRwrGRGk/s3bDBA2Ojjwg1pKLU+D2W5
bKaQWM1fwnbi/33eePt0if7thxNLH3QfHHwLJuh+6DSi8GKZl4sEI+96zPvc7iOyUAqEH8Zg67k4
ebnD4GcfTv5/GTIG+59Img4qKw1czXWiFgdtQMhMDKhBAS3ofzUO61cA63FImOUEoAiOM+0d0oFR
prpq9LjK3NacgSE9JGyM7xfazvdXTgwP1xAswyyksUyq1w+47CD4q3Uhrs3p+19f5tBwVFcA2oFH
3xw9gcRkqKqciJCLqtJYUYvi20zBuDnGSnwPMuq6f59Z5mPDjmvLvJHq505+GqGDHrh2L1MZnp3N
knOyHrld7KSBIC7cUsqmZcOtzytH+9MJqjwKfZ7so5R4gGi/HiIvcv/pKIAJAQcCwhjlOXYUICsL
KkEZlIaMkYdEqh7apSS3NXZ6c1GFLLhwf/Bw9BvwHOb1hhzPGRsSr+9azrt7ZONA2QP/+ETPB5vD
Dp00qelNM0BQaUDEIHahE6p5XBI4gHokSvtbOnHCnDuXrqxyQhjpWoHUDG05YCY7uo7ReAKDH7Vy
Hsi3YChl4GwV66127cbZxnfseDfXc9qiifkTIJdyLNEryyHiVrCaV/3yBnah8vawnJx+qFTsfCNG
cgsehcnq8Lk6xhJqKx+D3HJknLzA01xLxViCeh8GssusvDEaOOueCRC3PTwy00V2pkGZPwybfJby
vonL3eak3PJ0Utyzt9cpkSvXSgrFzxIs9OI+RduJyNR1N5a2oNUJTLsnueLvLCIHNgy/L2rtC6p7
mYjpJx5c/bGrkCWNMmmCl09oNCUscRt5pLeEObLw5kEfZ2qFLiMwvHRqBjP/Oza6UI/sMFRhpmAS
LAkJAB3E1uJ2gFoUXP1mb0LYngxqV1ktwFhINiuU+gvlSa92t4//+nZrLEuRbeUPff+q9tDaILzq
g/S4no6g1FJnqI828QA3axr+HfVWL4JpnoQu3TQHqYy8LaKxc4JlB1r5LnY3zfSogj7fo4o71U7w
qJak1QjCqo3AQqjKTigChVDGHImX3WRyk2RRTDkeDrbx/kMQv/gM3vk1rMXV1ZSZnefrexygAnGi
Ip6OmLX+nHny21tOPZbW5U5vgJMpcb1KYu4RRlUwMrznV3YnSipB2QoDfLf+yqolcqiGfSH+BnC3
VWNf8SCCU+y4O84hznubr1V+MPikAcJM20kgZ6xZHeMOwHS3bmRLbTTVGLeIjsSUQNU5cNn+COGt
y+u1aySYkFdtyA7NuuwBeZ1gvSBQBMYGeFj7+hy/+k1Gh6uHhDXmi7oerN9xR+KU6EnRpAQExMKt
JFOm8P5BQpzlgLuy3BJvhzcYJwgBEXgACFTS5ENPUaeJ41tsAJdwL+zJnJym2FFj06zMOIGPZhWS
vbOTIeenZhCIpoF+nH51VqK8MKFeaoYrel+hUH2Kwd/SvnvhoJ21Ls/cLtCI5TcCUSHusuUqTaaY
HCu/Q9OADzEfVs/1pwHhE5c2Kl/PaVMB1WmVRcJn5pbb0JbfxJ1srr09I91ESFOUvy9EteZFNVGJ
zriummqwFqudVPUH7LjDD5i0T1wwH/1Yxk1BdbR3BQs0MS20DKnq3okBTAl3mhs+mrIH6EHs8kvW
jOqatBSukXmmLdoSanJaWqWOIayb4qy7Gti1cyi0MpQLBm9TZXBHusQXIsevzRKuXRMAeIC5Ax+M
4K4dJP2SlnKhp1OcA/ONko4rA0WprO+OZS5rI1A4IuSPOOJH5XuO/IwQJRqNtudCtDa85teBYEr4
5U1J2wF396erjTPQaU6kgO4vsVGXXO/Q913J1h101X3k0DkIefD3a15myaAwPcT+lGi8MMi4ZXWY
+ef7Sz+uqf0qMoun82COt9xWf/1a5Q9BEzWDs23HszV2T7N9mVHgnaBZ2dEMAeALYbUas4PklTyc
mxm+ebpXOKAhXevld0iuThh4p3E4AcVxS7Az3n4SO6iYq8P8VWLQFDH0Q+vcakJQIki1HjNd7WRS
giC8BbokHw5QYTCfV9LEuk7Klituf8HPPVrO/Mr8zuKNqmh++EqOKQls3vxfNxcgB9m5Jn1pzqQf
ifYwAtkdIRjEdWgqp0mC9MlZ3qG1cLrCRrOMoZwSNpNQktOLkK8dALKxYwqCSEzJH9m9bKqmh97a
h+39otbKu5jUSJErCuKGZg7dAQWV8oElZs2Z9t14DigrUeUS0R28nDZMofpDfBbDlMWPtvIrBQKr
nPwpmLvyuamTETTC13kkZXIuUV0TwS71vXy/tRo73ZFvK/IBi+jCVlkWA9mcme4a5P8CerQwhPCU
Y2AVAx+orLDNPb2+M9UYD+wZJ41EciZumx91D45/YnT/0wzIeV2JnU30dbZA5HL56synbBCgGrWF
QV6DOMyXB+CyfotQl0TIFT09y94iRA/pfSC1LFPUzchDCwsuZuRRNHFznQfCK+R3Hrq9GFHQKHW+
mwGd9eGH1N7IIxh4jBjotnGZtCFvmjWYp9nTnn/wjx/6TlYcl1EfR07jppfhvugnQ0AfrHbXNxU3
jGU24gCvaBg+nMptbDr1wOr9AvM7GSl81ybYPJsNA/cqJTSxrI+R6WKNgKBrLaUlVRN5YHs11hWu
Z4KeEhzgDhDHsCohWZsiR/q3Oe4KmGK7zf9d9qfXEzKvnRE+mOk1tIUDM8Bzs+GwwTeHhnB7dju+
iF/bSZTACJ+rwf5tAZ4pVTjWyWHUNRrjLnY2zOXwbz+P9S3ioQWdC13pLRXumse3pRB4bYdSIzWB
jcc3LwtMVSOYlwkgpQHQNsNQN6s/g64xeV5/ioOWClAGYl6J4yu6TR7L38sUUrHbvg8cBFJRa8W7
DZNy7XoPoB0219QzcGrS/dYjSSxwUhNyY5n17i9pZXMMCUARauG+tDZnJsATC3AwNQMDnhKULyIo
KzvQObRLPrzOYV3okUMtSBj2LWtNeysPKRK+ZNhkL2JIeGcUpW4RtyLYQwxWC/vsEGAcQ8RVD+jH
CTirWL4HrxkAxTvJHoRzuRT2K4qjB9zemE+ZWjhJ8xaUzBkQ4JR6VbUQywzwrQuzpfuDOc4ijSuf
0gAaPsTO9v25p0fcSXdVPAwpJhCY9Ns2oyRLvb71SglhbVg/9nFL8JV0dt/eDu5dl3gYRb3sBvnq
bChLpJVy0rXPJHATmhg27fBiBopTOWBkwZiL/nPwSDONw00UiHiaonUC6j5zwmchwoniDEvFIflp
wG8drgZqkQivM1yT6j1PXHurkRYS2rxCq8mRK11KOk+/iO0dF5Wh29qVA90TwFaXGoD/hTZ1BlyJ
W1xLIdqJQH+OeyqfzV7Fjes7E3gLklJql6aefaE6kCoBaJ2akZGX9R1XYl0BDl/uFU3GGnjH8xDy
0YJAlHI3ilq8rJwcqjFaApRDhUmMzCdbWz7Pfo+J6PNfvBmLFapqHq5YOJyPCWWyEhjo0pe7HKFq
YHcx/npHaVvH5vYby+71FH/TrYGDDDVsMSCtY5+vne0SAgSvwiHBzeqMA6fiasJWfas5PXYX7GdK
7ChlWebl4HdLrIBFTevnmRFk3o1hGcR2RsaQqROeXQMbzlZ8va9FPu2ImR/IoJvhyZrFUzuNeYCr
0S4gZNbo52ZZjp7kSrH0+rXvNmnytZhLjELu8I1dSRQ9TU+PtYR5kJOPPr9fuX95ABOpxpdOqjOg
digs572lH4yMNNjW/8CeQvBphcaPOlp0cRbEq7ikWVJCgcg75ZHFHzF21BK5+xOKJxL8e7CItzRb
NlY0aEhoDMRvcO5H4v3o0BS298Kka8zEBCupwUhNp6HNpY41B6SAvTnO7xnbSqMOXsQPsrHwXSlE
zb6szBoR8uU7QMFZSjp0CyyTIz2Sm96xDlJaE0ceRnkH+cj1zPYWTsVVdH5B+qdHYIdfbPQ29P2/
RfNpdfkhjDq1DcNjJXOopvp/6dDvT98faZTFGEAQCStq59xb8nmfFnhqA8V1EKjcaUxhbzSb8r2I
Dl/fXoAU6HcV/hznLDMzgH+LLNcVnoDMJrNfrUgj2xVptDsSXjcLYbMk2dInDvGmbIRJ2ObSZYCP
QY2SRPPrNw8SvABIg8WNIu7VYfhbPXzhR5uvVWsLDp8VjCU+AFvLKkIHQOdjsCjdF7V31PMMEcyf
uGVkjOdysOd0077Ov4RTtcPIoPXEXpa/Nu31MEng2TY7zjZKrKht6n98JRgmxMEUh4vePaF88XxR
71NyEEkYBcK+d/sbASIgYTCjV1XaN5Xet/Z2dHGYQLb2jUyxKv//cl4ECvCEamO/8UTsSl3KzXgL
sOT+j8skAqto9qG+sfXfrSeEayYr20LyY9YN/RaunqDMBO9ztkhhZlQ0BkRe3FPtNK7ubMiNPUPY
WKkx6UBohuAEtqlIzZapBJFrchJ+cE3gLfqdmbK+zc6cMhvbTvpA39dYShoVptEEarxaR97sbL4A
kN9XT4OYEyX2wlHQYSm9QWGkcFBZYrzJeQ3g2Q1bRp4ZD7ui/GHub3DulrVvTbD4jzpE02QFMyXk
G1LUGc1KkwjYZlp9dBphT6LuBvHUW8KD6F3TXT4tFqreldIEnHT/SfjfKGcBqhY0Jdjfut7aGwhm
SBAerWPuo5800X261JWJXKnw9dU3X3mhcaHfIy/jitRdoVy/8YZkAE6+viBji2wQIwGx5q6tarEz
1J6xmOfUD69B/aBwnKDWOpAGPdpbhejRJlBPj/C2H2SfqLhWkBVAVFtVpWnD8icDutcusjsKw0t7
ZdmwdihyEBJwAUKUxyl623OqY5S6pXM7X59y/C1gWr7KiVqar/uSuy3atVPPRbo66JhT8h3Ky6/K
HEOQDel6IlnI/l2eo/4ZE3N/gbmc2z0WbRFDkX/NQ4i/BkG7ym1F+W/U2WLGHrhzSYc+xJhkkA/D
eHbF8r917vDwP6C0R7zyHydgIkmALzy5/69oo9GpmnrRPwp3ZYBsfv5W8bALyA+LWA6oCBXV+vRk
MVdz3Qx3zoQ5Lpuw1RavS6FFvkItP05eUt+RvHcZkYfZhhcmOJDURFl/arnt6X/dHvBPhbPL/iet
4N8A4YrQszTLOVyJey5+UcSlp8Z/sQFFjLlF4uBo0jSNsELgEJa8/nIsIjkty+Dv3qIvqVtY0BwE
+j0U+GKuVKa5jAaqj8WTneCDWZlwVhydb7hIyJ+JM/QaTH9oT+Tbu2BjgqU2DNCzWKpsiLlfzqdj
8JO0S7CHQVnu+j9qLuF0XUSgXusEq8N7wHm/LyQdXNsJ+jJcrGXybPa/bOo9M6j8X5A/ePZRj4Uq
9WL9wk4mbPVnEehrn6vJwjotfTrhZTOWIfovZPeXlvPGIK3+3xRlKLz9Itmc3zsg8G3I2mO05Hze
q87AfNCNi6oGHGkHtIQH6EpKRy3i2Aj7Aadk0jIh680SjSc4HcnKle6J1Ill1aVlLrH8w9WOlqgH
wv6lV5WuamBPv5xPQeId5W86P4OTgfAZsuomiMgXR1aFxw8waYO3PeLlelcNMBTn+dxqTNZfUzqk
hLZhNtmHW5mLivEeLPrZdWC1bdQpiq3R68Yw6fFxcUcH59wSSfyjf0VhEnwAzD4b0kQMdP3AWKDt
/KZzXvQ89f6euNy0jHwSSIfIXpHXP8iZQEk+baJTb1fRiqKpdpLWZ1UHhw53C6y0FOSQCWfslM7+
z82lvc66ZMVtPUtRUQdppw1nK2FXr2ulu+WfYMU+MlA6vBOg7wJcP/SEr6qP75oic2stxkqKTv1a
p501gFOledJ6tKv4nmPh4WwrtU3iMwgvXJs+S2hiv/a/LDrdmjSCRQqKRs5OIlelGUSleguOfhzL
D5CGSptMG2z3UkMaMHzX9aa2iWOLeNqqv26MUUb8yXWPr0JnLHL4HoanXsa34iG0hrROkjh1kEEB
X+FJQTeSS4ODU4jOv6FQiu8TI2MOSSz/PsLd7So26RfMsVgp7hcxG7gQ/9K1fdcFMUKfyQWbDSgY
gk0z4Jp2cFHxcWgeGm8UngryYBythAjJKiS/WzLpx3x0EQi+orGYI4E7JXefodxiU1ANcTNpF9oq
FdmimCbX86npN1al+3S+tQXL505G64LN6rcLu0bWHPd8LcYg42x2S6gSow0BVyTGJPtzcaH7FQL6
cNkjAkjXSeR+nZinBdsQoITzboszN+0rlJUWSFrQa+vDF9NCkVSt4EM4z4kt1yDTcr36oUk1ldSZ
aw9Zf5M+1NWMeY2FjsL14OgYHOcDfiIaPigUJoPNIcg0NaJm0z7rjc332grc1lRtds/4run6M4GA
cvCR1nWJ7wlXBZVT127oq2MmzvMYP2Pp7kn5wp02QGvxECt7iJfNR6XZA/0RuvlwKmCKgvAjf9nT
UL99z1AC1KYPTYzxtFy6hDmjXw5nHWu0TfKNydxNIZyifQF8ywrk5RsYSWMmyr1yYvncSpn9hi1K
Ty+VO3FDCIR3+3TqceoD1/xRLyn/5+c7ZdtNTgEuoPayQJq7CqBr8suUmqZUgSZ2LB2AjDZ6s3sa
xeDg3RJsNov9zuXRn4LQJHaf2uSctJZNkv5wbIQu+kv6mBtBhglhexZgS796HrFeo+PCpvdJDVp+
xITkk0EQFY6PExjhEmQm+xPt/F+qsMJUUjlTbIzcp9fqK87g/3zTXsYGIHOgZcQv9naiTr9n2UMh
biXj6AcWC6jDN5o7ju8a1EJFgUjib1HcHyx5OaBpgHXj3mRzkcpwVGMskKrwUqvlG3AcsaFScyJt
ieQ0LgiEZvxztp11tsIclG3k0q2JXA+2YcmiDTbRvnZbWOk44huaTomdyVX9bvqmujihg2nj88Xw
ISe+42L61KaeLXsvw2rO0Zs/KeyXj5N9kd7Bzd9gDZxQ3nIz1UiN7DDWfKvtxAes1tWN+ZZZMYxx
SYrjDyZzZQfC4ThvBjR1a7Er+cnajjNu2jOC8GHBoeiTKAWV5KQDO64Lq7nX1cyFhYTftssvRk0V
maa/ev3Re25ogsC07Vs3KM8EB07UVaolta7k9Zpgn4sVufzPiOKHJfpoIUB/9Sv3jt87P4E15QpU
5vQRm5bgUlSDbPHFfQrNWOpHc7qJsJhli90EEhVZLpbQYmrHVYfVbnYbMh4q7DG7ji9e7EnFw9GM
6cN0/3w2JghlVqvteyDXbMTpcO5bY1VMhPEFX2kqD/HZBg5CtCwm6gPNmjaesw/akctPy8HVdiBD
9cGtAJusUD+WkBCgYRfh36Krn4FSRU0DEgbipDJ/ZIvmTnLOXSgoVAORvazLmdL2afBRxkGprpAt
Qp0ed3uP+u+NIlu9KJsrFYxpiBgQtdnArCiB+u9NbmlhY5SL1FVuCpfA1QejYDCo2aK65gCVs0U/
saxxk632R+W09K6I7GSMpMwS+EBYp/7U+CqOkwVWjs0C03p2iCsP377TDduDpdNShlchBBx4bfNQ
5pqCi+8XJzXYeWzEmcTeWYAsrb0kjp0r5qZEkqIL/vXzgKN5gXQDmm57G0KUXaxYavMDkDBpx+QO
9nDYXr0yLcgQ80G+mSrpgRSQfCTBAxc6zVoHz1RneHxatnN6qO855hkeIi1I2CgG8HrRHnf0vyym
B2hesOTTFfkZlwFzCNHOkjQMKw/vRXDw1AeFW7xyoq17CNmDfYGVgZlC3sZbpxCSI6Q4KvbBNwQX
bBewF2iw/xKh077zghwr+nZdU5G9KiM9+5NGLYKA4We6AOVplgxz9fd7vxivklQzEUZISf/FYWSm
fOS4gcXA+6BawOm67uUtdxTJYcpG8PTouiC4UsGETi9k1sQUzuWjr8/JaHLhXz3DLxuxhfATaQRc
fvqYoAp+B4Xl3MdWZRHgE7/02tqpH8zzy1YPP1nF3N5ljSe+EXCy69k0hE8VJuyP7RIbZjpqA0ph
rT23V6mlquYnzjn70EI+OJekGQ069jhqyFqNwTaQKYt/3qMSd9baLmLo/VjduOUHF2fXUt3eZCaC
mZglGzfoMzqq6u+otDEckJ18ytUWo2aKmB4mRsX7x9OQ2Z1/g9S/Xthf4wZjfM6IM0BGBZDa1jif
zKhOQZLFBuNi+eifbZhrWMr0ZCoWTw3dVHmIMr3iF98JgTJDj35fI5d4YODbaSTw4FHdCUVHxnw1
fSywd605n6zXnpzjSbqTDf2UfGVhOy/i+9pRlLGcjvXmCp/X65wuMkSkxW8RbatH0bPMI0xlwWvF
7dbN66PT7l+TfxEiBPD1FesWYDr3Br+IPBL5/rAn4vujWgJx5NOCJlQyQriZpRd7ZFAEUy/an9yH
Jdr9nTGD+jEJcXuWOiYb2qqkdGNQEJla+v0vb9qkDzAN8zvdHxk/hYb42rj6yOo2sf/rTZA1XuCT
ZXUvyHxhjuDSsdG/WRyS9INUIWPYjXOuhlYuxdsA8U943nACAc+HWasE9QqSeOESkHKCg6m6Dsrl
jNcBjR0RYmqJiCWlAihUUglxAkbuE9fhEb2TYtc8Y5WBbc/ObmeQdWGATo4VnU2APpNCQgHuSy21
sEDBJmUQ/0sU7BK+svyNLRbxjBcGaGlquq3fdrfhIJj6/3K/g1ZWac0m1ZeyUkWmDLlZ8HQRh++h
MQ1w95IruOaGQ4UJXBM9YXVqDrzt67DZ7hMFG7FPsekzjpN5RsyUDGwCj7aC41HluxGA7qtZ8/xJ
IjQdyGmuKrMcHrowucWG5dCgcUVTt8sK7pkC1DU0Dvjif3jsbfmyC/cpwMUNRyU5MIe4ysLMcDlH
QsDsIguTpdsKaGDl0E4w+cH6vOecO0TjmNBvW+LF5as0wwb84mcRtio0LFHxYFJqt8pIHKod3p88
AmeFnWS55vj7Pj6YClSjydUqBJftfvNS5r/ynLZTC+PAXg4LtM6iUCrGgVfREzRd1micOa1HYxzk
Nxu6ys96UFKVbsqDMQD4P9fFIU22c4EnLYx5HSOQjFoJzIy7UiHm4VUQfeOZQlzQpJOoxrDE2J1p
Fhp5PJGnmFdCasHvojrxNfz1cWetCbBHwngN/e3JmawWVfc0y5LdYswKSZAYDBLrk2y1IgMYe5wR
tAZN5sBHHfTCgsZXlEFjiBLGwEJgg4DOMxBHjhj6RKKI1EQ1UVRCqoYOHDhF/UvfPOm9AtU///qT
n2ASek+Fsg6/URlJ8/ZarHAprr3Ax8QTL9pBRa16JhAPqhK83m2NsiQM6+lUV5Xwoem3kuNR3URr
TG6U0WPcAcco3u+6SKCbnbuHQpGm1tsaUsJfc4B3OIfk/rF7IQK+XGCRispj00kICY0PjpTZi+w5
5ScvzyXMf1rLKdpqGjgzbCndCXj74zzJyST7BPxz5kCaizMazQtHaUuhiqw9yAK9oZMlM1cemLHO
IQr1DlZ5vd8Rj/HSQ/I+IFjenpfM1g2o5oP0uLgYFMtME0ZjNEvitQi4HQeUJIFsuhnhMfzOWFFq
ZFlKv4StbLZIyU55KKYx6q7M0EhNNTaqVlh0rucPJrq6mJvTF+BgZbKYtu+USA2xFW7ragx6CG5k
RNtiDJYJ9GVGWUPyBgR2ehEV4CwcxrlatPYqyfR2NcIP2vwVcY7X0D/hwiTrUCCWw7Qt+U75sCnu
1wUTAtWJgmrUQ7nLmxBee+sIoQcaoDCoRrkFZkL90mK2qMHn0kffnLEWh7IST10QYn04qJtQRUN/
ZL3t6xbk6KLfl5i1Fcn10MUcntJYef0UJfkUG+pTX4i1tZlKQs8rOdFvCk/Bszu5PQscsIHrzkgL
NN6mYkX/Rf6bNmaqPErR1265/TThEtJihuOmOdZ4thShkKAnYKYsz4TL46muXglaLHEXjmqzF9um
ORVRw/84XzOWyk2WRV/a/3j7C9aYKiQvRJFtZ0q2xKP/FJv14IosoqGV9/6i6fy/u3SECgnGVWs9
0fPVFpSftWLHM2IeAZgSMoID6jp0A+STH5v/Qnibce8YBUolp8cci6C8IPvUGvDumN4TtsaevrcU
1RFSnhb2dVECcARhFeU3KWuxUuiBneQXyK5rOdFJfqtiDbqNIaDpn8fday6ktTOYLnxrvuoFay1V
nC79DQhODO5vgp4tEsQP8x5udbnwGIae3oD79QIMQEKhDg4RWF35Wp5yI1zhkKZMEykW2i9Q1NMX
yG4Ji49Zj2C1rARbUXYMgH9zbIBfQ6vtb1fVEQj8IU8JuYWG+k2C7UOYq84eXoRTv7n5PGEf1jma
M2ybNl4isGtY2KmY2XpfU1gHEkhIsJYNfsX6F510rD89ESLTn08mUebLmSC+RBRg3tdyzfsjxazr
EfmG7sXdN6OqKA9/SOuCU15PqaPbSxlLVqduA0PzbKkukJ78oMJxvTAJ2Y3LbN0HZRmS7zQ0wOW7
/Y6cYAf8tDIMjQKtCiAbWEu0kNQDnLFZ2AfGJdRLRRbb4mqqxOe8/pEF0XMZ0bgNu0wtClv4b0i1
4AVTrDOhAAz2W4Rr6bFXOyg/JxdsVFnPCmU4zjOqnKsBEcqeEghtId7B6bqEWE8m6XNKUTU3sbsV
RxRCnXAw2qYmGMzrxawj8S9GAXCpL8z/XU7uk6ytTIfvwc52Y0I2QUFGQZQjHsAxi26LRH08+VZv
ClvkajXDjsuPm+OTwLv00jkGkPMLbXbrDIw39tNwiKz65+m3JGq3nH9bxhEF8oGLZBUWtKk7uR8f
XG6g3mBevGidNG4C0e0eTqrSsbhd+Lm6Oja0Y2jBWI61H/CSvmdlcI3j/umh15tMoRte2V8MGc/x
IKm3jdBhG+qZtVIjpkDRiD4ELNOAfsvqGgUfj2eiVHnMtjq+pW93w18I5TOdQhL+UCJjJu1TTOM2
sEeu7fLL7b3OkidzRk/x45JKVSMKxl+2sV0NmL2FSMMtNdxxRAxL+wP90dY8lSuWHeOuVvEgnIaw
jjlyOnL5CbOwIinCTZhoaN4GEM8ll/qqFa+uX11HilKXV/m9gjfTMyOrIUbtUR417QLIeNx8oaGC
TYQWnB7UQTZiGmhljtZV3Nrr2d9Zq3LD9mNL+kRgjxGNLT8gDv1uDbDdshQTtgj7mC8t0cCe1CgB
Gl01aJwfQILewKcew8THS8cbcPnPxUAGYuSmagi4o9vo9rcuVne+6l/8bzGG71EyLlcFASjr7V7K
2uWpZBKmQfJvL5vPaa3AaADKe8dmG47RpSsFZ4rxieduml2x529IT5djCln2fC97Y2xbnCBFrEDY
txgvPA2J3bdaQKAna9Bg3b7No7mUbC6UcnNq42bU29YkDkJKD++ZyJgJCl/VTlG/NQgS0Y0w3nPp
k4x593QPfxO2IMC8S80U/8qErrPXk6odwyNMXDurQc1ffesYLHmLwm4FQcqUWI3K4aCJMRKHOMC9
cb3DmPvlOLSXuAs852YsL5woE/XhPXFZRZ3cjYGy5+EKjOK/P0dUXt+/QaaUnBUjv5bwzW7B+as0
VWtQoFgRWk/pNJ7/5D75NAAUDlaTca3P7pWYdBv9sJpxSbLGuMFQOrW+FcafWxyUY493aTFWbL8X
UKtYY/IE0kJS1zb+0y8FM2plwFlpBktp6uffT/y93BwRJgv0ILXfw48oPVBik1tPipMLpuvLbABi
uQTF7Qw5crgYFAwNGN7HdlW3VGczJD6DGxTYbZmuqdSnhszLMze1uWIClN46c3B6VDy4vKlSa3Wb
Q03vrCY8rBUtRGEAh+gb65gj+Swj1tJOd6pMOI05eeQUXoTYjh5BZ8rMnIIJBOWL10rG50x9N1aw
+K6ayWxJbyXFthAZd+6U24esFCmH1Q4uHI6tqNIacCPVNMomVQzNMfdVYfoggYXwktiIEXFLr5D1
cZs31VIFXOtYQDyL13AS8ZCrdyUQRrXIYbDh8hpcF6N07ncdDrRaxKSGVXyjxFM0ZOiNg/ktJDIp
25Xfl2vt2D8jVCOwrQPhux/ZNezT22wAchfsYpejdPhxZm5llLouBaGjO42o6c8lrCGIxMkprEqL
xwEuzOvwhS7cnOXj1MzFGQT4BbVH0ZzrRgNTUHvrEdKXJXUprNTSiynATgUsPsPsV+VJzRUldiQW
ryKQEufn/QLB38gJLgDpk+HBVknNNF6y/PHo8SNgTsneKCJsn3WCBn567Fc6uxg6kPhYvxEGBDwr
EPiNoRh45cvTkXPTSthtJiEQAlpOlGkKFQYwVoh5CHaSvmI9Dr8vyVCQnjWCIpRv8DMxtXCb+Cqc
E4SMs6qf4qr2A6YBD6jtlj0NWWyj4I7xtmD4ZsjmKAAl28o7PYjBnRYyi1e7Wvf3vkQcdTqYNa9T
w3CnBsL9qJSE/kX++DyjBgInVcFYqG/yEYkUMwBxTJC8Xyl8zdVPSnpvFpm41fde4hEta63+wS7N
ZgHw8aj9r66AmWVzMX03Y12ZhpB7rvZzzq5+pbx5Urq36XJWXjavrCKjj73us9GZarUIlPEKn8u3
IjkjLIBYp9UnSxH/JA0Z1sll/MgRqeDsVRnxY0Q5wZQFUDWTN23H9j+eXgWxMD1T6+zP/ZIWiQ6G
SmOavvG3HDdGiHfBzi9Kz0bE2pQRZgNk7sTriKTEg1jHF5hLMDUfAHmw45fKAgNvpi7tCqcSju4O
e1pAvcbiA1Bpl9G4jN/Xi36J5+rVJlwTtJW+WY5zm3pct9v0A4McCNyKv+wp1tjPlykj6WxkE5lL
cypGI3idlfF4m+zpe5f4qDXvVH9FuhjdWX3e+tYvKUT/XbrMQ3/pwnbAx+5NAKl/5bmviW4JuszF
SZTXq/JKm6fTTBQlv5wiZ4BOVCWVqEzwMu58sEOyGWtG83an6Yl7NK7cF16thElUte5vJvLAC71x
1cLI8vFtJCD9SrTWcwnvSKMTl6GgYAlW8J4SQQx5+YKmpnQGfDnrutBPoflk50k+9Trpl5Oe+n9O
ZLpjCoZjupgQ73IOrdbCBtAGJJQ1DvdkNW4pbyVBST3QiE+sVx05sSRq0FQ3GZ3FXg35Hn6wy2+L
O7GClEbPLuO0Q2tY2UQ0RcEaeLSXe79lpFlJTUYxgp78gjx4VdX24Vp7bft0dBJCezhGoej7RfwW
7BYctjdHQePB2jqA2UM7JpJYWDzDP067wttlVpK01r46P+Y8YRtAcVPvtdyVY4+WY5HKOROqkjoH
VGKjEHt7KA9BOh3lZOVZUF0lKt1CCCQ/+dqO6vZBIdssxdY3gMe3T5ZfTAbKeN6wTY8hbP1SD/8i
fD467/K1if5/vn8ear1C7+IjCPgy+/rHyGvfabEfbeBtZysyx+8apfKxI/ZLt05HCgGZx1XQuQ6X
qdG0xl/N57GB532a0ds0UDCQX69cTGGFpvmlwQJIPAqQn9+q6eaXevEUwSLwiIt9U09KKDOL9Hku
W/EZi5ExkPeHFmAvMTlphTfokr3gL/xFUxD5Jaw1oDTPNh39xsycpdzukMhKiDSEavnuQJtwb39O
e4JouinFEksgu3dOnTjncLW7KX0lUjPy/bElXG0QEfOuFoJqndZeSnGxXWLra0uhREjm2P5kQIVS
zG4BI2drlP7y6xlYt+iA4tSPTBn3RNBRXG1T4wzZodMQmjWJ0dUshOUetcpXWUzMn47VksRVVQQV
8We1+ppRqeEA/m/LlbKPDPhDT6uSkGuVbYC8Pbw0DJexUNpoLdKIxX+d6SiAwX3ykNGbmhynSAY4
K5e+8oPgVrFOShlv0dK6HvMAzGWxCKMfRzN76JCs/TlwCR1+HyKg9Fau6ezAwBPV+qZ1aa2DlGfs
BvkzScWQqBktyCQQMfAgkYPIlEsRySnZRbHwZ1PGhGDnv23tD+iFFbGSZvCNdJ5NHm6TDMz0uY/E
G2KknFEKETlHGIQT9usmidnENwNnlhpv2X53VA0InIbOj6UZPzx+1iSlA3IElHSxke1vrcGKvnuo
eDQNcoigRXfF86huFOpnGMe9t8avuOmPDmdWvuwtrqmUj0zZrNl7yNaqbjzbfXMNvgaT4cpZ2ZDx
NSgf5HHEyuYR7bqS3nb5lG+bwnnDpQbxOzCCc7xP1phpYTwN5osGuduApq/7lyUGdjlg7o8KCs4W
VmJPUwErnbC0eGSwKZLOb0x13ZC/woYGpW2GKi5+twdz0vMoAqx3jt08o1OglCpVoo6LRBJdEFJK
LT9c5womKHitHGl6bLYaKtnMrKk/dzGU1+9ElEMliH9AdCsxzaqOqwRSuxgKd+jtWUb5Lc4TtAbB
UOJ7uI8GYateFglRIZ5OEZYqJf9qbAFmHag2Am1GA65BOhcW5N3Jo3Sz2qHwTLsmrGena4EgzpSp
K4twzOYmkhH5TWmTeQUk441RR8BNnK88GU91ihoc5QRlvyRig+qv4/k/U/lCtBFdHpQlEgl87UwB
1j8Lp1gsX+nzQ3E37tACSMN37KcNV6APjsSPzj1zERBqgCkDpvGzh5fUyPKVafyIxdo/b/yWqDvM
eGnObn2bxHHqaNCi/uHM+BbEYoN0XSRlgBsOfN1rpgWR3Qhi1ikWMgEUTFb1edIj7c2em3nUJ1/G
7Lvx7oG7VoEJSszSTCpSs3hbKEanTdKhnTUInqPDXSQ3thPasVaoXPE5vXz1DjxcLB7+a+kSQ6Rk
HKL93TK0K4I0zS+TfePwz2g9VwTv6pJTrUpdsPzYI15wSH708RgN+vSUGrzicdcyHv2QEbNbdNTU
w6FoMbmE4LeRe3XHtDvCUTUYioaMI0dnyoraaNYFIXrGL5xMcsUXYVm0RFdHOYoGCdn3qM+jwk0D
+7LuJEaLO4kwzxTtPmMGUL7UQNkJIY4HHYX8Lj7lJH5rpirhz2oHdM6DGBDGEb49Y+BqIRpchCmt
9oQGGG/8RMYkOG0vLL4F2Yp6Y7NbJpXITeE5HgKR3AXeI5kZaNmAn8mtSM0fJNwxmkuug2LBURhc
FzIy8A9DT21dVjsL6Idro4Ic217DfZtF+8xmGVvu3gYf42AhLrdK0VGK8n26z0suLN46TFdr42/w
sGWHv9QmsthbdYBchw2pREODuV6e+QvMycMIcxl07EVF76bF1nvTZHgtKhyJeiC2C7M/MXNrhcSY
cT5mju9MiI7G1mZnl5lD5oAJabWwak7VrDuVad5nBoHuqHmuYNzWkViGa7YWZyzRvoK9TEBMbGjL
xQzbCEu0wE9btjZT9cb2nnXnb2b7e95dsh54saZH9hvLDIzuD9V8R+EuqYDjT+kA/Pxh3RdbXytn
PU6DTqlWRifPka8DwoeY250MG4rRKCaY8Mg7IeSrLPinFfeOcDACxTCAx1TVeTxlf9iw+2U1TVJ9
Ta+Q9Xac6qI/P3QRCI7JSKTiRc9jAjNlsCG+az4gzvp1Rg8lMiE6PPpZzwa7bWv00cqITU2lIggM
ADVWeXyIZB9JVf51bv/B/h9N/kM66KMOgz7hSmhTQd6y2Kn4bYZiUGfZvOPHJrWQ0jcexh3jh0LC
dnVLgbnfxbGyK0OiU0Rp99ZVR+V4Ie/CRyKr0WIhPmPTaUGfo9L7WLEhdiCqv5alM5xlD5Gk+djW
9sOzYUWD/Vs1WYqaEPFE+AEDXtQFStILT3e/uanDQkj92bMi+8eCjRh8nDAlK1sop/SpmM4M9HtG
2pwgGjGRVcMZYUDxg6XkQdfsE8Itr/0WP4EoHkxenaIrEMgKDsooZUSkW9/YRHc8y5159/4HV9nB
NdBKD8NSP9T9vQwkGVIZ9aTi64mhOTSg4VjiOplxtAXVXfZTLy7Qkjnj1OZva4n0DRW1EMIujgJh
6JIgqVsqdYScvp+FQ516wxKJfnc1CpsCPBC4+uIFC6nv5Yfta5aoRtdoknosA6IwT3KB73v5yJV3
HxY9gh0Oy201CIz3B1dqmNyJW24TGC6t7f+hzHl5jPTQl0+Wul5aaocE9segkec8acnOj0Ot1AAx
K326DRoFISKMoMgWULCnuKRmSiVD6UryynDCZIkPtI86qY/aDCAjdMSgZAz3jlEkNw+2L5oG0jyN
XZXNoc320IbnJwqm1/mKpmxZab8Htkob37kjL3p67K+9pAkUMVL770Z90rLnbLu/csV8ATCmYMDA
PvGadxCX8iLtL1tgtezCff/iK+RZkcZWS4uBsVCwCEAtqiST88kIXC0TWCmCCLXxBEutEH/YMEZr
pcBQYDZ7vKnV/Kdure6FVKvPstx0UBLCadshfT/OwqD6Bj8xPmOMYYd+WPH1Q6FBaHuPTwu/+Vs5
jus6BDrN9Ty1XBxf0KAhSCMKFRrk6YnvWdM+T06amZWQTJItxNLxRpLlw77bxc7F8PCUBkiVoTTg
Pc9XbnDxdYIXvojKA9G71DDiYi3QUFu4weigWpKMZ8DYRWXB++qK7DU0QpnoBJgqvNDJ+D+5AK+c
X224EONJSKCnHxM5W5zJV11mgGz0WUHthr8B9JvXvDrp85SuXk6+eN8+yh0HT+Ib5Y/sfXGnRHoD
BsCC9+n80UJejtEQ3pltbX2XqUXEWbrqUdWpwpdijUGGn8cPdhCvawpf86eCcEcHjtH3uar1ECal
c3Qau9U+D9nN8Q6KTZJnEm4aFX1NwyszEqyXosaq+AIex7NpxtzuHCbI9q+r3nL5v/mUZ0/ub4r5
tivDRJWGrYd7Bps5hAVm8bJGijNabETq+S39Zl1JRzF3FRCg+35SseeLhSQ4mJoaFU9dEa/zl2w1
Agj+mckMzzVH4kvhchLAuqg9d/4KHExNiAFeAQ2DeIN6xOTmG0RndkokM9UGIb4LBXUbJpOO8vCY
1Waixscuwz5TsOqwSRNre0+8uEwSeLHnlBM5yWYu3ETFTw4VHj0p2G6AFjPtyt17w6Hh0Cmj+RD7
d4Sg2svioKYJYDXBEnfx/SSvOtbBSSYX+5zhTTbz5wdWBvP7V3JVC1TgbLNrngkKXObC7aRrYzyU
SxlrdVuE34RSXISP88J91rPdCF3fivUxKuxHJJA/dEV/LwDftvE8mv+c1cJ9mV0IsOFEBY6SQrNY
CEtZktWnxZpQaSJJjFVsTmeMYhZFqkNMgzlvBrpmsmz5GAhBrVfDhXjgk+xhSC+M+Y7ZlxKtS+bT
ejlHmMvMX5RZgy8aWXTDR/XI2WJa2/5WS3Y43jPnmF0oQYLxMWbpPsREssoAf0J4/YyhMW5cHuII
omTj4c3tOs7oSXrr3oBNRyx5PChBup1zZz10MT64U4mrLYp62muYeOqXqXTvasMwWPtiuQk1RBrV
Efg2abld5y0JJFpyac8NlxkfZ6nS/jpxBSnxYKWghxMYODcR3GEZyNGgaHdUlItGHs520mr0ZxNU
+ET0hkU2uSKd1pzA1tMHx87TsvZUvJHqJDppHXoO+KPwX3XZV67715DXAARYViU55l3O7jGcTZXi
IIh+at7Cjud+htuxSRBSx1jnlSyq+87z85y41xnAiiz7N9oqXQbIsh3Fdh31Z3xS+9r+2TnNUm4z
QaX9fLuHgKpv9TYq9WypRKqKsAnHCK27I4w2Hox+iyRpf4widIcMq0u86UBfcLrARq0HYWSIIjJB
gFFmO3J6tU/hUzxUpYbTtSiK5E1J3fxKQrLjl+qBgqomLyuLtSF60kKW81n9oKYHZuyIYRgozdTJ
SecSft2uU899Hiz9o8uUEq6r6IOZWGICZBo5DSKZxj5367A6F/r4puvm6aeEwfYF6rUS9t2U2sAi
t1Wd3vIuKTA9kR7TACTtZoTw7l3OCl5dDXiBPT54qY7q2d7kpYpUL0MDWNHqueIGCojQogedLx83
1nNx2Srz2XMEb68fR+aN3fkNd0llU2qfwjfzvmJ4jK4URiOgYnswdjZfNlB2v1SbJeStPLZO45Cg
JYaWPBwwhLqzorX/MP5wsLf7zvbQrp6D5LtpnvA2eY3pLbHF6xq+5EHWvadZCBUN2MT61Apfu+xo
dRn1WX2q5/PIpEPNJafprVOUGoqXl7C2T4ge8oHoWF1DfwqjNA/iOIDCIXeTygg4HxffIdwRpyKE
qlh65hksXP9qeEoz+EPj9b3My4wp22fXavpuQETaxWI7wLmHdfrwEkSoQg9w+/7UentFzQrCKr4k
NmBKPH0pnHoky3EmCvtjAD7eHycSs6ETaBPdX4hZTxHzCNM0gFdHTYiHmCQIjrtWeHtjzd7wEBz+
h3h//WY2ohNs4LDpLBoTSwg44NUXxUWlsRg6vF7NRkD8VbH5BKp+0NpmnUOl4yhGnlkoS6UgMlqP
ru0fEh3QGjmAOGYxaV8bH9pRmBxGhsnqxB4grcXMOp1BAD749YGU/1eQOfmRZ3Xs7SiYAo8ND1Kj
htxl3VOf/XPpwGbwQPSqTjA0ZJURIXG5S8ddfkHFIGI8rmw/xqo3lkExJp3xtHnxfXIlyD1QeK+C
fFukBrchRFrAXIUW1/ry5sWX2YNok8ScG+8aFNsOATRX5XIU3NMxrO2tpTUnVEh0GtmaJUobFI5M
ZAoZUAr1uzmKvoaNb+s1GQ8jfGsxeikkyX+GmpLIslBsvtzThcT7cSVZx4qoJGOIYaaoBsbp3k0m
chDYLs6RNBioCT3F5KiNOkQVqx2/nSujTxvQ1OkgINz9UiJ68AABvnBJqdpp5mRAyfBVV/zxXz3n
JSfhYIxRk/xB8oY4bx/xTPrfS1+Z8hVGjYgmjOIHp3KiNkiD/w7o71hQ2BZ54aegwjl745vW6ny4
A5uL9Lm2/aBlnQwjYsDMijDx9uaQx7ffFiqyCMeQ3MONgCm/4zIjDkUkXsLWiEZnbUXKrju+2Ugr
nu7pEYu0A7L4Ike5ovV+1/K+P8EDS/e3SxxlAiY+Y+3JzAYSdtfm3t+wVAO89m7IvxEcusF5gexU
IECiNForyRbFrSs5Vv5h4jE4/Kh2L5XpddDwXYwH9LYxAVFyLAYui5xwHKl26nUi7O4sjY+pp/IL
dxM6ig1BWFDcHsewSZi5MkTVsA2jSTK5lQ6NtcM/5MvkYSFNijzdRdsg6r3vMXeLpUFDSaQLASxc
k0T2525Fq4mENhXxTeSPLRZsZD5IsAAFvDLw7SOUdO+qTvDCHljjtDje4rrXr1/tyUf0DLIQufK4
ddkqmQCzhX3+S5xB8qm5hXFCbVkbYi6eSR/WswXEfz5zrY7c1g1hM1CGaEvsuLxz7rS2vIW5PPPZ
tMIs1kq6gZFNFhzL5B9Z5bMtqKDXR/hLsubXha0I9OeG/0ItDAR1OVTVhmITuqMfX4ImF1RKsMjW
UDmCnaOVtq+wq2GW5K+v/GbydPem/dm8nys8yDE1LrUMdZJDjLQXug1BEUrWadqEKqX/dO2yReKv
41mneEY0oKXg64fMzoZ9y2pkrH05QsB+zLRbfxgREtNtqkZvhf1H1tPNsv4Wyit9oGckKkD1nj2e
d7TX8IcM5frbhoGp4wyR67bjjwUsYzCuGZXd3cN4T+EXN8q+xNioopZXuDfUDV6Dtw8NRbTl5EQk
ojHeKc4Dsyi5P5amv6q4wGPy0d4brj8LK6V6X/ZDMSszMtoatHqYAypbHxOzkSMosMi1gWs2O1T0
WURvZi4zaMrw6CkWxSYCGshPOtWNgu19TIFmBiO630vXmK3X3r5WkvEhzII/sIJBrN9Eu7KYroIp
bqlm4CyKKEWGWFHJu0PPiQu1MUk8qSv7VlQkbwOtBIhqLxRkLFt7uK1zzRu5iXudsmG35fVTUihG
cN9RxI6PA+VfOtR1fOPa/f4VaEqvq2uxeahfXZ3wqSyLOKrx+det23xrJL/NDHTSoxiKYwPkhg6M
nLOJDFWKv4530jE8CM7Cz2iaIjtJYPgQO7w8ABjxlfVRKbjGESjAauKJR5+GTI7CCFMnuId4/2kJ
3hN0FyNDS8exUQZqclyeIOVPSW9ZRP7lwT+Ig7kiAUDv4FW21xGgVYSNXdiehRnyZwypXU/xj7Mj
Y+ht/csw7oHQZgEyG+wfZKlZ4TJneACkyNTFGEEnPiLgwyQFJBLVlJE/QCHJmn2kA6CKWHe7TX0R
KANW8ve7EeMAkMk1SE/5Ecdax6MyMAwIm5CWyglwEcnVYF2tG6GNnoz2vnLtY9ybKK1l2YPS22ut
awKxSsY68tv7UiJHy5tVXCHmjgohoQIqjYOjXZe1IVGiC45wTb4ief5r3YStevwpM/Psqc6y7Px+
6GOymk/5cj8Nr0Z+aKF53Sjf8M4B0yAYeCNCouTQaUArgP9NtoXAoGBQgeXZZ4OD4S/G8tOonEim
ebpGgf0RBg+qrPOrTTiw1A10JaHWEjoTnSg0XQ0hx/Q9YYGRGnotBJZ2odFzFFPQ+3b2M/AXWbcL
L/grgcjHLZ7iMmYEVJxgLVLJPg44Wd9ffcpJulLA+VXUepwO9FX86E5+BOgoo4shmr60KIl2wuWp
Fryd/LEdMWM8xnNolSSG16rkgIoHOOzS6RCuW/4XY8Z9QWBJ/HRXgKX3Zm0WnfcNt5xR/6KI/pQw
3TzTzIZ55D02ebMbbna2PRpmJiFPG4Q1BUZmK2SHSMSc9W4uexwa2hom+9lv4/YziiEOYG9rb/9Q
vdnPwbZcDSHK9NZadOMYe/q7JLyVZSgfj5gqr5lpMgVOvKvmcAytOK+7xG2NkZZdSk7eqLg8SXH/
Di45GtahCC2ydbwc4FnKKS+LcEpF1IlGPrGGt2ZalsxRK1igaBiLNFC48Ao4hpclFiNWU7bWxFIL
wli3IlzxtNy4Wh/pOm7nu0ENeldmsJE1wpOHjgMUo+9hQv89pN7TSQDI1hu/AOHlU5KzLNYWtZ6r
yhvQZfJaWydAlz0IhXX+576JS2qg1IXN46pZfECF/cskIzJNtwdK02sdBrJIBVl1C8nnH78WidwN
lZVmtcyPVplAw2FW1A6pR09ep0rlez9XcG6QWsXNbwEkicYRcsN9YyoMEftIchP2vp17oB6P1rq4
gYmsoCmH+OFtndESxE+ZLhS6Mzlq3KAy9wRZujvvIWaPhR9dLPi0k7yj4Y2lpHf+Zk+YODkoYsb/
QrcfeglbwriAF+e7vhL3k6gSfX2bhmMBjlJeWSkAnJcyu1Rh8XC7KkwPOczwghTcYNm2YckGKaNP
aJ3GrbUohjA6zZS0As5XL10Q+CiNloaKfrObz8CC5XBirRmosYibsTOxzD2gqzb9YM/3hImeJgdl
B8FIxw8nXQVQyFfbMMb9/YSKaCLqkbm9+FP7rloRH7Szq2dJuC3eXCEtaroRtsNwRpRSOIVd6Dr8
/QfJE70Dp4CnMx88wMPiSANCg0sFOL7oF2dOoFUxlYHYnoYzHitGWJUg016heFb/tvYg1NbYSscu
0gCljNUgPhGIU9lJNNy6N7figzVaD5KTK2PcwZuXDr2cOnqyYk9r4+RMhjQE9+KP8xrmK0T49vUL
4bHuHtG3bvrpEWypfQwRGA6r7efQW796E93EDKi3rXyA7uZl4IiAFWA5kb9hNy2D2PfXzb7NCDtD
4lpWzX78wDUYo3sQSZ6j1sInJn4ni2QOxgfPNO/VM9D6u/fPVaIqDUaiu/2Qc6L+8JPiN9NdEQU1
fS/IbRzPte8+8zGUtwFgXIRJxvBbbwVDw1v42AzIIrnhZITAxoLlce5U/qupq3+nUPrwZzYlSnRC
I3XL/iM4+V/JELA46J451meTCuzUHeKv/MwiZC65Oq3kM6mnPvH/TPUfcL4dNl80TFHWtAHmMOe5
SYIpzhxlX2iuwEYYOEX2bh7dXfsqeq3+VVR3FInn6h/2gc5k/gkRBl46qr/ioYAfZoM1os7BrzhR
/3wW01k+Ni6/os9ilybSBUXnJjVpNFDEP7PUtwk7UmUp8QpIvu4tGjpuYlnB8/8m7+eL6CbJRzO0
M+0pOhQUfdXrGEuiFHcXftBPjWCyhV7ipWvgjogXdcmKg6VmMay4jkCygHCFCyzQEU8IIllWoDQU
mxhg89W/lvlC0CPAZIB7P3DEUINs28QR9+aDOI+W6Hym8tYyPwdsSmCHJ6TDquKFqaFD0GnHhtuE
yL6CVh3d1Qo+fN5TxrwkiWtgpWcv20degHNjwMdrB19dEJKbvoQsh6bf0TV16spWek4AnJFqrwPo
AUJ1IpwzElBX6U2XXnQjpg9YZ/RZ22RajyzosS4R58srWokjAHSGdXX3s0gyanr12PHsZZNJo6Dh
ZKkfQZT3zFbHds9exWI4NhrVS3oe9GZAYR3SRtsAkCT+t3X2henFuwA0I+sVZtmQSc6UoGOMP714
lGVZULbb2nSlOOp4kieiItbCx9YLDwiLbKS73fTbgH15QZ6KkC7L2xmtX0tnD0/hW8+DtuRAz62j
pKi5XizNj3m7Nl/4iTlPr4d3vXQ60VHOB/unnQqf0YNWKUXJQhTD+c1mNQVum0cFciuBY8743z1d
THW5ZKMbUrKqOhXSfhcTSB3LYVM+72TrE9zY4p4O24V7avaAACMahG85IUnlF+bsR5BRISR5mLZF
5j5uUj4WG/bgE4rQMH5AglqFkWyX8q1Q7cGM+6oMgbo0rEDxCRhtfCRIPMT9IWAoSLSbH2rqRk1J
+EJH/EexyoFy2EnmLflgi9MVsjNohQw5CL0j2Dymi8Wp0jLHKRzChWE9qvyiQK/fMht2njmoCrbw
J6JyQeX7/Xv9KneaKTtyaRn215Pw1sZPjn0Rfm8RCBSOFIi1rRjTDS5PULL+xIhAFM1r4VPjKtkw
xs0g3R0F5lGwJNMWk2MN32GDNqUiQnxh6Avh7DvItaBl6OugFHFPDi17plmIzV99i7FVaq8qs4uB
bFEh1RzuKepoaP8rXgcP7cUPQe8xn/6FBgFF54EoDBCqyUIwXvlODAef5jRlz16Gc6vDgq3QlGiO
RDLqeBSjXWmDNLPaacqjSq7thkWUUzzrqXaK7Ku+mF+qsQ36OOJNzFOVIXcq17dLZRWKAV6pynIP
5VMBV1p44P21M4h7FYVanzXquv7UZa+VSZF0Asmx721TEMt7j/lk9JYMq/lMI+kMoM40h8W5tQHM
Rq/0grVlNFM4d4rggQDeW4p4KHMCmCnmzVIoS/EEOApmsRjCoU3zPg+hhdUetLbVkUqvpztTdT0i
X10CK6TbrTrYZ5YK3bjHxG6HgjXBPWc4zxw6gf3O/3Ez1a7zeNNCEpgl01QkP6QsHr7rdMWAsGs4
GiAfLszckTWiRD57XKrsK5xWFMqkxZ84/CXT/APwn4cKPZLxCmtqkF5iXqZM75h2/5meQKYRXT6J
7FY3EC3u18Gl/0W1uiIGIKvgOxW4i7G/QRAfDYaYmFchBhEE5OHt6YSir/20lJxdV9DPbZjPTHHP
wq2gNSUkMVI2XWZ2ANW9LlvxQxnxHNq4hmc0/A16c9WcR2FZlRSWaVKHj+qc2wSFS2kSuyNLhGOY
ee3zoG+5SfXD9WIiEZPT7EO91kVyVSaEIuH3bDDEJz6WP/eC2JSGQXrk7wzp4x7Ry1gjIk/lOAqR
P3DfjDQQArKhsd2lERXHyNj1KSrnxQbiGfDQykLaExh7PzV7peWCmOJaSS7ULjjLLlmpf3eNcrr4
CyLVU3DQO3Kn8whz/LtGBaBTaCTEOU3/yh+1AHOYnL/ErsIEzxcHXFXW/9omjtAqXTae9A3PYbU6
O6WXDL00Jqg5cIPOdyCxGVAvnazxXk4YR2oS34BORQm9a7CMf/SMdUBjH5johaoPlzhws7kqmtnW
ee+lUGmNaoxtOXlZ0Zb/zcnMR/hsc0gHI8zOR5fG37zTpNMWS43lEQi9J8xPNeVqwNpwItyeSsb9
/vPIXwIv/bO7jh+oG3yJL/4kuDBLcuPJAmp1MgU2cB/vSJnAVqP8B+9nLDly4V+yVoZrkDKxVo8U
p+MR6XBq4rhcFg0sDHVdXEHHkWeE3z2UgNuYzH8ODb2mWJbolp5HpIZQpc+20v186C5tZGTtJEQ4
4ZrGmo86T6bJ3bBMZzqrMaEEHsEwjwMmDGsJqgWuqXTK4eRWCM+wbQ7Ab9pYLMtf3I1J9R5c9UzL
hjuYXL78in9EwTG9JsYdEE6goUpo6YlkYE1hL3NTlvnq2aq9d0+mqzfJS+wu6c6YD4I9F96XJ9VO
4tloAZRRdHIA6Dww0LsJhK0qG7Ha2pWelu5jLr6Orn9u88HRoTil0iKMeATKBuRhgBtKngUehOzc
hTJNIZwmk5R6AIRlPrqgxPM/kIxKX6MllSd/i077t6sIgey3jhob+PZQj0MjgEwgzE6bNfvB2hY5
vwME39jrY9tnfyv8+xRQqVhSRq8m1xJ/ZuE37hFLo+lgFXRtnqfg/Pb3KVqzbK+TLQBpm+KLgqWf
v9SB8KK7jSawixsuCvepFqQAC8pqDPeuBto4zrtGqchkI9y8teUhZSoIcKMc8Xgey5WvLhFry4z6
st/JYA679Dk3hEuxgyXPYWBei7VA2DG0XQSETtSk8GZ76BUAvCSTlc3TA1f5cAxIJrsTp/PkbInJ
TE99dnepZckCvi7LRyTJY/ZkjDFju4SY+2dtdJYWtYjWq5uQCCGlzOdi2ebwcp2q0tU8M2WJpezx
UarKVTC6DA60Aima32B1su+zyNWERbOHBVUjSkP+UGtni+kwfJvXsH+6HiL7MCJrV7YAEGIT1dfI
KighlbwlaoDMH8e2ZQBnSotGc5736OgLyuFojcWWq31gjISpW04ryLQwdliYfqvtyGyL6Cv0dwUq
hMwsfIcSc8MVyCj3PLJpcnHA1dfw+j1s+Q6vl33NQPIe5k4MQ5SYLfpc4rNnHH6ajGSzyKY7p32D
pOgX+pFq595UNJmFwxx97/Ba8tJ0Mpln6jDNCV/L1wZPvI63eafXxBK9VWjnTXb4Eg7wUQ4x6kle
v/njhm3qFB7S/RZ1ku4sdYz8FWCm0xzn5R0TRGq6LZ2yZeQK9wqHoHl4DFG8UoP6OYB8ejJ/wXv3
bzkXSpG1/TpjoAi1f26VwEzjBxhXywRUOFlDc8Uq+PjIlPTXH6C+iXzevl61ysCqXyiL2GKSyWah
aufuSIiHxjsnCD/BmrwBXdRzrh5veEjP4vBdcF37Uo161MmEzbQMa6oCF2hHBrWT1wtS59oFjtaH
jd6D4NP4CyE4fxwN0ifMsEcS2ugHG1wjqQlfr/KXt3kA3vB07uWjLfyrb3i+GGwm6QlbZNYn6jP/
h4Qy7HIdAfzicDLKzA4nLHKsnXVtl/B2U//6DBjGhoCLrGIlUAZH7/D3OxQyz3XIIDtlzY69h9qC
RpLDzRoJXfHSd+76nr7ox0u5QWt8jfOLds8blVo4bzd8IPbMsXgJ6JaQkp83IssGEQCc+lnzPmj2
ENiPGkMG368HpgN+aor1ZbYDiCD/prXy4hHqAwdrd4fKco8/LMIQBZHJSbZ1sh+R/uMON3xsvOLj
mCPoSD0Ut+/8EXjjahSvBj/a6YRzfr6diGaFowtYlvgLja04fvUCe8+/m11TfiEkkVrHkg9YOqIm
WbamTJrjfPXcyVTLuMWpycc3MPijKmAHiQXdrU7iHxyQ/YAJ4WJSbtERd5sM9IR2FCONHpvm6+C6
UMLGg4PpAPby/1LC7fObKzniNYnKcS7x6jzxAtj/ONRda1KeP5IvTLCEueootlgKCtfiLsAuItH7
Wb4x8ePb5XWCG5ldg8qUchveM3ICIameBWxMHGpgvrnJ++at2wa7qOMhX8H6Hy/OFnTehkwufXnw
cUhtEB/nLpCZmseegybUvSDngRSLol7lVakrnFvKBaLYAfUyWQzjlzfp/7/rjTYk6ERVY8o5gGUt
VMrBLQNAdY7ZZj5GcIyzcob5uGvXix3N27Bqhj6gWZ6ZlCEo2/6mbnfzsL5p7aKiyPKNJOWwq27i
ykRRjL+THrv2b33zWAKh4kV4GztOhHrmRgihiWI2+K0P1CdcStTRu2of/7PLInBHRm1Rc1lQSF7c
1GvUFMeBsR1H9zcttFSTz0y/55l4v7wRzoraj6i1r+PPOlKOY0Ar+Mo+8beFvoYAj94zPe1iuPfh
F+uViADZa87+O+2JQOe4gii/cCIru3j4J+Ov1u/srN162S1mEIKLdvnao9HNTy5iQLNiqEHSWO6J
26fZXAs4rKlwuUJrrDiPaI28i+zreJ6NT4NNSjzeC3fkmFDtP4Chah1s3412EL/fIINsuC796FIi
VyDmFh/qbom5xophTvDGCAoauem5nx/0Z8vaJcBflUjKz5M6cwLB/GmdQ8rw4fnslg0TPcF8JbjQ
RFmL/pW/o/7apS8Zk4uIYUlrd175jYhAsFZoJ/OsTEm3mK2+mJuP7+/QhVD2tv4AzcQ13k3X/lTZ
4LWRORLtmgOanqWTl3kD1iKxOewu4L/bnt83PNFjEGldyuGgX45QWCBHj6QKcXmmTwtYCUYVaQcL
AQh32CQj6CN3bHPAdebupT9tJzOVQt6BwCwP87I0KgQxMC/+SMHkm+i/7sJUslvBq8mGab+hKbhT
4zLXcJOT8DqGL4EwdN+muwY09uyV+0fyT6YvHF5jiY3fn/HiO4PSKeVX2f9oDXZsUZrdj3ljZS66
4K488L/rWmpX1yDaIa+Hk4OAdu9267+QSU5e8NJpjv1VDKstsYWO/Gtx8wfSMmr4s4LKVBJiD9ha
Chb5az3JTxe3LUnIVD3t8ig0SN7T94jhPELA0v3fhU0cBdL38cdIo8IwPXIxpDooeQ06aXfq9433
lvQUl4fO5nP7GX+nuxzxN1WJSsqHnSP0w1s6U9Z+Zr6jZRaLM/CVjUKhqMRqy2FnU+4+NpBjK/iI
pGx14W5QVfFe46mC+5+9t+mDbpqBZGC+4v4dxkbFQbM1WNWx1jGcozYWeo84MaEa88arkfvE2gby
6bj5zKvNI4WxFt5ZxnxRPxvzrdgM4QdTFXo4ydN6us4AP1SJEvXemJP6+TeSoqqDhiYOJ/BctJM6
zG4JN9KGju3DbVphUXlPxoVdkvrCSWdH2KjAbGG2TFR1iRfKujzrAK0Ug49fUiNdCwzYlhgLxPoL
rjnaLuuIk1eWZ5kW9V61PKfsUwCO4gjUK5k8IMgorpgQR0hpCjBdY5evRoDSpLX6ZpBx77SjH+g+
ovGMfKf1Dtqk62v+3aUlEITnD4TXB3gbJEB+2Ts37yBAxebo4JL+P1TuWd4R75cXvrASD50kNpEc
URLf1ElSXK+pTxIUgoW+NI73KK0KwY7TEnijJqNXiPNmxdw502MynxKGPcb/xyZDXfL1wEScBkIJ
T7Hlq/mNYUgMgCFfWk367/axiwXsHY4u9pzYGrSHiH1V7/OfEE6pEyMj4oHG7nn+h9/bNXl00qvo
faryAg+h0t3xXqx8CnChfk58xbkQfADBqDByBn+kVCESf9y1gZOpA0diO6RBN5PwBafbLCQMNb4N
ON5GROlOVAKLANkJo/oj0S0+G2vVpIuQ4XT+/tCb/44fWVS56Q5cAAALOjqbRK3qzV/AsiF+zeVX
KxRRqk7YIB3hFb+FHomyK2HkHH/zG/W4Ruu0+aqG48py89jkCJ8szuscSAklhSlPjdkxArDb34PI
sf6PE+nplinKRgZnWvKAXZWdMclXea9IGjqyst7Kz+sTF3OwUKE/QTNbn7C8N1sc+OxKQRqdUhn3
9/RUmi7YaliWBKvDIIP0b6eDAKEENAhkEINgPD1jmm9KuSboYn3txI8nX3OhaamKR99l5/CLwqiY
Xz+rQRE2jrr3G3zQZktbIZO0iq5mUVG60S4q2o/yIFmKa2w6p1QPkY3EsvZuEg2MyQxld9Ez+Ots
YauotjCOfAWSErAh6My2b7SgzvdWgN7hVxsK6HRqZStoSkzyRSKNGmSTdCNg44hGYs4XMKLrBUMv
Sm03bVwaBTIyRfOoYvUaIoeQ/rIyCzit0DoWNbxp8LU8o3eCHONCkGGnXsIBJQaDidHP+VpROlFA
LshjAdiGwaoXxKdcvEVXparuxDq3Bkzo9sa55H8MlLYjXck1mh9ZABEHZHaoSKewdwHs13F7hu/4
vDbtNrZ13K7i3qqrYRgDY54pGWqUWFgijKfRlvQm/d6YuhkfEdYPL5qr+wwkgjuEIzfyjS226+cN
CUvgprKusdM+gPqy6OdQgnBA+3LCb7m+qOVD90baS5e2LQ17KFOQvCmEM+x/efYcr0zz9yQgc6T/
h/yPMZpj2gmx+FzTdcsYtyKxkZ1lsV65rUYQ2u6Nn0YzEAgKR77x8FvBuI0t+Hf46PZhLgNEG5oq
qXiXmFfAWXQ8aFprAj7AzcrflMbDT7VcJFfHios69RO5fvevCFh/r0Y5H1WACH6rG8WNHWhiXLWV
KUGOO0gepPvCYPxUxdLVnQgsId6Gd9z2ahYBw+mBx21GMHBm5OLv2fVJGtvJgrYqGDOz7Qnm0K1K
TN4hTosaOWIl4zDZ+5J7D1+ohNpm1mP0yn4yqrcey+K5QDKJ8a6JsZWPiMGGQdb5faUMg3Iot8rq
65jYpw/aDYXfpOIODRP5myPS3jgkm++t+dySRyWf8Fq23YAv2z93ayY1txUxb+84mnxMR9RQIyDp
E77IzcAiISc6Cq64k3cI3KDB8mS3y0r4Jxv1H25Fx6DfG76Bs+A+DtfNq0ukZClkWs4QHv8NVnSW
7re+k4U6kTaywFc40jjCUH6XqRjFr4pYedKVqL+sb37ATDP2inFz8nxY2GqLxhHAumunDYHhncRv
pim6+cE72Oz0VTY6OYLH/a3b3zuC3eGQDsATSu8Y9zFFz5uLsng5pigvCIItKkRvtOHqGHGK3J+3
kTo9aByJmLWytTWgRV1bpZccPlrZBJ2fEQoHZ81eyifhGDZ7sp0gLeKJd4Ez87P3TconSXTaNNeV
baiLNHfBt4d9ey/EawI5Hx/ZMolTls8r9xzEhY6uWkVrivlE5S1Zcl2x+8AbBW5QAD3BNmS/gN7w
JywssUai5SKdbspN+qRHdc6YfV0Jp23S8Y7IYBXzce6IsavIQA47RXZIraxrmISNjopr3qL0g+Z4
nzXR8X3PA09RS4aZAIY/mJVpoPSvUT7mIPL0qBeena4OmNfCH1v5Hkj+ebG5lV6peRepHzKaYLlt
Taz1j/VENh7F38cUoRUaWCcNYJbEaw5lCMPpjGDA/25Nnvi4dI0dtL6FAE+PUj1r7v4vSEgKR1gw
1vLTcB2sMV7C5w2kgZ0ht3CHsmm3fOsOYNuqJeX0DcxLVkxpItBvWxR71Vl0l+uscrwIUaBW2337
Od6IYEPAZJGca7LztJ9t6ErnbCpBQgWubmuSylpeNAxqsnJtUS9FLTg2Rpf158FlPLuIePac7i0F
bv63tzKRlrpSNQ6bVlNu0OxKa1L9TwNzMkEGjIsEfNjCTXtQggRNT9ugf93ltQ89HKs7mv+tkvU2
sIp8/7lDrrnjzeu4lpVkxCTjSUCTSvkMRXp215bwmP5wwt8cAXMlzbN1/Fs5pW6tmfm7THFMedv+
iaf4U8I30riIzJ0VD6cq9LISp0DoogFdOR4pESbJZ5TOZrc4JxV+pkLHIbevN9eG86aXT/bbrCEb
PLZoM8YxufA9pUvhHBL+g5cveDTI2d4TKogo5lUvcmSbzL9Pyl8ldGkcGibqeWlGSQoSB9v7T9ob
fKQhtU0MGirSMlcGbQg2hQaaVWNxD0wBeHrwaZy844566Tkgd29GEg7EzjfbquuzzbmWiZv04djW
lgKgJZfky3xUcPcWX1eyhw3r3PBnWShrKI+eWqgirdVc0VIDq24x+3cDak6tX4D03bhGbP6Qel98
qvOK8ZFRV/TU0jgKLkzjVDBGfS2WN8s1tUYgpqC3VT+sYs4HELpI5wepBHLLxpAk7AOrmhodkV0/
ZrDKJ2N7nvVy1i+cIXMqHhs/hATBG4DtkA/3tHEVLt6aoX06St88Jv6iCatrp88itzXj+7I500v4
oL5iZOTk3c43/+WiSUax4pRRk9pNWqV3JRww2wNJcAlx4K0dyPAhd4v6PX9zTwNLTKktakgQqkBG
pefIXcYJA0Uj4EtWQwl4kEwAB4RqNl/EESQap1Xkv8Eb2hGFGCUFBxeYKdpjKDv4SF8anLnyfnA6
OLAyrs8ACq8hqJx4Azn3F/pZA3cQPVeHpSJdfXYNHYH2Kzux3+qqU4VKTPjYynHZ5Jv+yw/6hku7
bcfzwTqaeR8fI8rg94hKYaAtPgFEblmzjv5/s7WzCqYl908MyxXc9VR7dtbDrLzDtMFeHDd6U5No
X0RCSn+ORSTcKXeDRFcHaBSURU5bEQw0/2pQ5B0ip2LZcCb47Ja30ftqA9g1zYlbyxTIlFMsMelj
e34RMSNeXIDuQ46H4+1NXmqfxgAK/bv2zjQN7Z5KLNlVLE4MbCBCGji8j/7+0uKdxcd3GkAhWRos
277S8K9h5N8OYUvEPGD4VOaXKCt5FyURUjiNur7kop2zERYyrFtPQCz9SOuYZk/83E/wfV9nG04e
LMvOicj9WHhLOa7WizQtL3ebCN99FQncT3fiH1TQq8gl4epaNA1hppd0A/RyyzD71KacCwnrSQW1
riw5fOhUT+kvvV9Rn0T9RJT8EbALNgPzItZ3aaFQEw+c8J8JvlhbEcar8CYkWqi5EDVtxWM3JS6r
CUNCTnV8GPTgPzoltzaYatgktQHya8Tjoqfu4vOz/BzdFWgvDyuRgXwGJHC5HXerif4KmSpKRJil
yY5ysMa0xnVM9P8ECscsxCWbb7o7WnxDLKuCMGSg9/yogRnT6WHHHxxXW8MVSkjv/ALdmkZhq/GN
Alva11KPrvg36UGGKgCt+KuIKXZId/XAqK1U6a07toVUUr7Afx8GFB9OYdUrEPi+FqJFo6dXLLYH
ZrYOuy4+JZdzDRAthdRp+a9JNEYOkSsaLUXfC15NZtl+YtGRcmOf7wbqNHfV+YM5i49Qssro/jII
ipT5IC9hOAfvSIhaocHu3BU7VjBqsJn2Kqm6dfBE2tnFHaWGxkRoGzXUXjaZEmwdjEY135vt22nT
UXyTrsrjjo8XDtHPQpSfjLxpd/azrRTuV5KAGdghr21W7N80bH8povaKZujsjSmPw1leLwHqYMYI
o52fscbggFKoj1lOhKhS6SGKFPUFUuKwsD3Y+zAT/aQjo56nvb9yGDx6UhvSyDEIPvpXy3Mvf1MJ
RqaDx0x1JDBZQf9g7h57wKeZY1IQGvzrbuq+RTXGWUaqLnYG1w0iBf39vpRHptBvJrOI2N/l/fV2
vqvzmV0ZtPVUN9uOGbc73H0+KQoat7BKaRxQPXCYPgI0Rro7CYlEbwq2MmXSClFdtLp0iEUNIsxU
sWvD1T47/eQziZnAfzJoMMcesbmtMH/ouKR+YBBB+eBo8JqRmp84vPyNvwfqbf6gmVuYngMD8Dnm
NI6x64M1u7fWGOt6uj1rn57wT5kYLzUQQVfWYV/Q8Zsb1I/GW0SypAOVDb73ZtrFL7EUrJO/9CGw
WzNCXcyZHYaK2MiJXjUbpB7PHzLHhbZ/lO2/s8DA1E+pkamz7hTBuczTY5m3gFtCqCPCWSo/J1Na
CnjOD7R+1d4+pbKiEcdT7y3kKiU9zFIi92lUk7IkUcJFEIFb2ssU+bkQNxVPNpSAfUK56rQvPPPa
oWIFCS27TirxefdsATEkMWlo0fC2ti7aDVdpomkH2GNXRKdgIwxXhVZSjovoHKnfX5CjjI2xMpi1
eL9e/uOaBu9PDfBPj4JmmZ/qwDcTgXLT7LCwGU4fuzuc3C7wxoj6jWbPDlDDTlTG1OAfNvGtPePB
kZM2Ta/s+INxLa3vgexhMJnd1FX6N5K6PvMkkUKKAWFAfrU9ugBcWyYYylFXsfqxU+FdqU7hSkE7
G0m/ZcU0XJTUsSnLKi8FP5qvDp0hdElyib9dTlPq7hAwso5sN9P7EPD2K/j7wAvZzPlMdGiGQIDW
siB4iYHgfaN3fcSfETyJw/iy02CmlIO/AJhYsPWRVTNYLbR8gxAwYpscHoF/m6pqxsoIKcH3Xknb
Ghs4nGVgcquiCn22RK/AJPs9OmCoMycQYzSeMNaoxdvGomS1YRZDPoBcfoJ9TS0LJkAes5l/sps7
dsf8PqkttZ0z5bFYbR0OokYOvnN6xXDuiTjxZ2q+JQ5mqGREGUMgxdO8GOmTvSFNTFzNK+JqaciN
79ZdthrH4XevkrOIT/li/hFjbp3OCLjZ2V4z17HSoaJNCH+EGRv8XdnAn1cTT0HZkrktQFtufi4/
gLZ7d3v/vgfgkNSSkZdP4tSb1qGxYTMnvtq/T+I+YUNs2HGwrtOpMKU+o50yVW6JGJmlWA6H0MO1
7NDUMcG0PaBB44gVD64bepjarSaFbWjOIpv9MbsX4LCerhog9fQAOJ32DulQiBpPWKJJchBNgRaZ
HuHWQWePhYJZxlrhGNVFExd/4+xOhBPtH8U2Sa4CqFOgc1BmET7jSdhgRntrl5rDaAxWn78sDUWi
2HXvXn3KUbXBknAc63OjCpMhWVdIQV8hTz/HksF5VLwkvvpmUQgYrCcwwhOVv9sXI6v/ELuYD7nP
5A+9DS34K617T09dfu5RLbfjqWNZ8+jiqwyVJwj/ueqTGRSaUOClmpk9PjtuP+l2xgr7UE9QYLMM
rbvBrETrqu2CMXoCjQ1GlGdc3gzC1wlx6nzibYNqG46DAK/lKX0nS/zMeKozJYmDcol2ST0aGS1Z
D+c0hbdR+m3OB+QJ3bnEU5+S5ZtVep/RnXtiItt8SbhYMAlB1iiP0QqO+/WvYRd9rUOGwNG3h7QY
oy6LkwUuRsj3LHEmwPLZ2u5MgmX7jh1Ivg4p0bCIU1DmZEBDoSfL+tGx8jvjObOq1UoTPnm9+Q6p
6dSvpc7rqqpSkGiXflUNwua/iSpthQfrZbUyGlEA1AVnQMxcf5+aqvfUouDyG834ooo8rwhGC62b
TqE+mvTBn0NO2AOemh9l0FM01LDfXv01LY4Hsd58vVgBQLUP32KKr+h5BTUp0841EyOqZC9MnM+g
rcdhytGiH0ZZ0Cm7pYIfb0uVoR8TrVLd76e4hWoVBqdgJhy6/G8wg8JlnJNtGXFDGlvgXKQfZtSi
RuSkSZOxiQQxCriJL/45t63bdMCBvNAgcTx+l5grB529uIc4NP950SLpC9lsgVjjgRBzswgdwHUD
AY0Oi3diV7nlsZWFWm/NB8CcN66II+Qk2SEgp25+Qdnen5J5NwM0UHNYlhuiCVnLb5soZaSYOz8V
Pq+VPXfvpu2bhvC2kxASe7pwC605wd2NnfCUrAQw/g2E0gYqsBwV6Hb7ZnZWE0wUkR1w3mqdkFnn
2JxKRSgcyPOsMEruYolfQmGhYppdtAWqZKG5nuEKp45qxbgWOIfitXe2WVJawlryx5VS9YNzArqE
z6zlvPn8uYPDAYfifKTRLg/kks6qx1lAYc29BdcpwbI6r9NZe9JYVJT2z7EfDj5Hts3p7d6VmQPK
FZe75HZm79vVhTptLOjFvQW3aU3zVQfAtReEmX3Fyfvf+yEgokJkfT9aMBoGnhFeM8JqZVG2RwAt
onoiM61PUW/FnHDu5BGY6JMqhWO9sH+vFhm5NDo9KUo3B716hc3zfqhHHfABownKTNJytf/0mGQE
okQVCqwg3a8RiOikyCFabQAfdeE30WCZoh5ICPzKu1cxnO5MBLoZtKoSZ2//UydPchsEKKzXUbls
oPbVVS2EZtd5+kLshyje2ah71ZRT+UCJQnTj4cW36mdWZG1DzGgFvWFPswo4DMiwY84H1CRMv0QU
c20VkIUi9vRaajNCVnwuO1cRLOZTDvASmsri9x7ruCs4A5TcbhPp3bUHh2r/mzmmExzKNj6zM0KX
bdKXJEJtjQiiK54R3I/6dsUYWTK1jpsLmCt1oySX4a5DRrhvhDoYG+O/kd3JiXsNDzZcnTKNv/UW
46LewNXzSmTGfctLqEvqBgwcF5+GQ0N0IeZmFfqA0A1woy8oGO1SU3yOoudvP6a2KDwELYhCAx55
qUiEv+KSYzEZzNlKHh9qUfm0gDewabEM5Tu3pm7KiN7BT094QrUv0HZ/o+6CGOgY6rSmP+XcYlxK
ViG5rtHC1khgXApPZvVTlXuQdFUAXpw2ctFxKtdNfyfsaCji0qibRjz0aqjH3qzNc+64wlxn7Mqt
ZfteuqN7EPDITQ6H0OYm1yDDeaeTFsrQ0EcIIVLeFtKHBJq+syipmDSbnZOkWQNJrbDh3Xy9Aq2v
jTCdKukSDpmJNKjgU6NBBffE/7W4mDhsnfYsv/yrwKLSDlTb6WjgOpx+s2PgzQnrZo1LZuvglOUF
P6MtUjzDLIUxnmq/P4jB3Po+0VOXDZ5KsstTK7IHDz/Wx+gL3sx6F9zpr6a0dDURmV/XpjMtKYAz
NnuxJ8cjINraNaQjGul/2UsH854M4S4r892zfiLEXEIIVUIsWyPt7/uJ9pX6ClglVi9jdmeAROwb
UYVOSGWdCyx4m3IrqSPmI/BBvRSmRXN8XbJ47T4LUPlwppZ7pRckNV9iXkk0SmuCGaw/4kGNzkvG
unW/b0n/LChuQYd/XgCber5tzQDr9CqfkGGHvCr8l7r+FSvGSFylnlyCvOoydtPE5AIiX94gvBlB
+sfE5IGH/azeUgKxQf6mmSLBItL1ZozC+S1g5qDjuuslgb2DbbfDjaqIFlgd66FpuhLbiryDc3OS
m/miJ+FoVxNmJRg4oZlrVMpL5KI3LjyaYCwzR8vxZ+/m5Jg9Nmxpy4sp5lo6DtWz2+dpnLSf7eBZ
sIH+F1AN1lazwsedxTY3FF31Mv261Ip2rlCdcnTWXKpct9L2h2kjEM+jjyMYilguAQgXOzeX3Ngq
g9RtUatQ1T4scBANH9OOpk117d+ur7xgF321cdIbU6LVJFpLRokn0DGkBENGge8gmpfC6lJxfjc7
LpI0cbqDqng+oF4Hq2asxwg72/oeF06pKRJixlaAAvI5f56Uq/kuiSj1GRRL3018ar1pYuvtmaqH
F/lgy1fespvdl/Og3z1vkixkXJMplgim04PI4oz04oCQS9YRfRCrkDUrAkchge60aGCD1V5dY1iB
c37sKjqIihgFaTidUEb2Y9OTG6TMpr6MxEr3eVnd7egXDY6+nY3pAz/Zt5IGGT9MBiOlfPJYhYP/
2p9LOO8kRSbddZApC9ZlDBZt4Tap3cH8A3EXu0Shp3O/+O8phSAgEYLpNDiwADEarx4a25tt/lX3
18YJRbsWTrm3GbbbQBv6K9HABImLlOKpq5fyt87Cgci76YDP/EAgz3fNX4q2RABmap/9R187hdO3
7Qz08qhmuMVkkP62pl311heZUDPiIaPX6/rCIcdL/CPdNZfBvm+M+59MdwNuixwzR/rkbLhYUXU6
Idp8L4GPE9ibLBbz/ntISGn2HncbRGiDcGJ4RbBVcLW+4n1f9sqdRZjo3l+AkPx6zG2CLKB9gABy
jNUq4xZI4KgXAjubeW9Wc/4Rc74Sqo/0b+MBGEjbNAprm3wL2FSFgakfQ8YhowDyiS5XhVQAXppS
tJ+pmO0jmrAgYh3GWK5Ct/yYXjNoex5iQfTMBidvVzp0LuezkOu7V2M0QOSNKrU7cYd8ZF4aA1t0
KhcHKves57it3Jq1SElT5kgANKBKVPUvw76aVJkwLbDLSCCnnD0mMu+rR4p96aYwhv/BKYLtZ0dL
ury1iF+rTKiRosJ2W/tSmYM8F3dYe/mMPJlIXZfnIn9bfLmou5QOz61g9cUcbbeMWaEPSNHUDTfx
Jlm2wrAyUXH1XIjMEiEiL9oodTqsaOowfNkFVWKRwdhq3CEMZUTIJ/j2EFV/jxJ71XsJ23tCXZqs
qj+puaBo8SOlz5tsIAFjTAWvNCe29uXHRfraIhogYWBRxBO67vdD/GYF/O0YLIBFeDUjTXnLMHWf
mVI6dkgrVnMocDY3kGVeVqwOcG/UBmLnXNXoBNynYiBZJ/8J8dk7OjomkMhSyUnq1vUL81EvKUcN
NcaJrRDy78d9dKNasPpk6LBSFhEckxFntjDQ0SlKD7hqnMweTxnqqE8g8a39zYLxpHnlKyIjvWe4
c4uDofMICz/ULKJKHEl93wNmD7K9RrjfR345QEiuIY11fyTFBqS4X6Q+Jb5WjjSD527VhlHGWiWs
Vpb8bdRTrJ20vUlr38UT05za9unjQPNpd+TXvzkV4NHrBII8n8tIujYf9fd6n2L3GyIIXQfsmZbO
LMMQtKxwj6ClQ866W39Yu4PB/vw2Qd2xgK86AK0GUQ5MPugsiuLEMy5AleNZIXCJPqC1WGjPu+AV
vf6KyRGxGCJ/FZmcfKTPsBPIDUjnRTDNpVSqmgjhbuNr6fBfZQVRMw/IFlbdcGpFKRz875gOgTJl
I07koJa3ctf2igfilu44/CZwQKLe9cWFI1zu8wNPR1ZxGOn4l9j8dBwhrIKUwxV0IoG0E5V54FLA
k5LcyBkUTo8P7XNJfNqQZdhLuPrPIBCZpMdDDyC9Y97wHbslyhBOxqZ0Sgzk37iAyyQuac/HwlWP
OyUzodsHrZ9AsYJNwVWswkVKu7BGtn95zdZ2CQlHB7+ze3yNS5qEDgRFqLhWV8PK9EI5VCvqH8v4
TJ3W0is+pww04GxZUsHc0TkzNANYxHhxen3l8NGJCv4IjV6VV5k1xjPkfwjOmPvd80pomJ0shsdJ
BwX7GAXkniKG1PYOKdoKyDQ6Qq2bEy9w9CCU1zglTC14YRwJ0C1jFo1PNcEXNzZM85hbBVkVckGV
YVEYW7AmeyQ5wyawLy1ouhISmARpKIEfWGnyhe9CCxYcC/3/0VKTxuPp76IrTbt4tWyf5riKOfZR
dKDwcHrLKCAe+QTwOZBDD/JPyI8VralUP2Hslp5fyRsDvS0e4qd/H98S1pAx5jtj+3WVbWxDnw6q
20GIZS8KAd5zy8roC3akJScAqSPufxJBcOMopfuWp8EQH34s5A4uit1GSZCu/Xl/mA7iWyq2h+Ao
bUw7JfznBxOmnjfphLjlaMSBr+4CSR50gYhknWwQP4btM58YEGkTPWncjYrJqzbnPl2GW4VEzB5I
3HDLOlJz8f9nHwAF3h4G7G/CfVeERESjAaatzGAY2Hd/XvDJLpwdr63pPkD7EjR7BjDX7L/6fbp/
qls2DGb52OOiC5+YUGB9DeJoYdcAb5vFfDseqlPExYbNGhh/7PTb9gkQbj5UIig+DCOR7at6smmf
8AwFUGGXZos5ByGI5AcMiodZIFyE02xIys8Cc/8EP64WPmHN/EVMttiGGrNDZUdrb9Bd+YvZkLGG
S+f4dDAAeJF1u5xOBibh90cGqwaQW24F1QeIbcbpHKqbZdbPHzoa92bl20gPer1RDwjGZZSo5CML
DxyABBYtjaJxPcMgjbnCv3Wz/JIkYSq5yauxfkd3fmKd68gZ+x+NpWL5lZD+/vOqPJ2mghB91V8J
DgclMHEJOZBzhVTOc205w/2+YuU1ObWmMzoWpYcDPwUgRNME2nl6B9Ip8onr0YjMgdDZFDMiURPj
seVg525neJabaEhJ1C95pti3solw8ZY6Jf2YXndOGltPYL/MyCibpsLPI084HuwKJsfoAm7aD5o+
+1P5JK/4rft/eQvU0t5t8qbyGjwjteSlZOLC0aI4ofwD6w5VLTKW4U2KlheJ+3SPjdAStFOcTsxA
KM5lZqmYMtbX27DU5EKEOa2J4PBvFUAIXB0zT4As0JC5a9UV2KADdGCPKnuNdkiHdprZnZwdlXfD
Ftn/MpXS0DcqVSwPm1ICuKCwfyoMhyzTTvD3/TsafX3QrRxvxePngYOhRETqJv3tUqyzhHN4ZDTL
trKZ0tBh54stch75h2KCXkEBBCzZOJcOuTmzMDvNLSkSKxWen9y3BEUcu27I2RnyvcOxjDIrDpR6
9gCL7bl6kZCLnynELiLQDm4CHHtW7k81scv9k2lnfb7DcG+Ac4bTZmnVySWEs7j1y3nc5//kPENr
t+AoUYKjnKWQzXdJPAxSMCdOKA4iaSd9IyViXvG30JmbrHYQvVtAy433XTG8ZA/mdPsSuaIOxJbz
Ac8JTOKT2FVenDqSb9Zm3Bj+kUjNvRs4K80AUywoSxCNMhwbTmb9L0vjF4mfHQ/IsKsBNSj8cNdF
mHtqrM/ciR1gWk9v+57xVXz6/YE67td+WGFMgqerwNK2GDPnDKjGHiplzpxzYu2Bo8M3D6mtkjLa
rdMkHFEBWwfP+0Dv9cd5+Gk2uZ4+u2qgJ1/0BQ0t3j/OM6kqsYVMWakgFpBxk12KpVzaqK61TLlB
VB/0JZRd4yypknpvv6Dawt1cY9DzsmC4WREiUWArW8bxxmMiIlbFOEv7GgS/vTnzreOzdmgZk0Th
Po1SdL8k4yUqqPJ7U1pZuh+hjMPSIFW/IEz2ipwuDRJqijd31WcZ56MPUrJdjwVynXkxm2flh0pd
jBvfN/0kongmUG1wNbFbf1MPS1d3Oq8A9xr+1TPU1dMwaxcYVzbB7pfZa/bUhN0FLDLfd9REk2aq
tFpwCn5ZjvLY7OEAKP6HA3GbwytAtZeT9/6V+IU/aPmyW7CZtz3UBlfELmf2nS3F0WFmCNwSqpt/
4XOzpYNn60tHeJ16V5Hd3iyRRGF9fspuQmovdJfeURJMJ/JxHf/R9gU0S6QcbZ7FSMwlIc+64OII
mzMuveVBfSQfTB0/EY1XBtyNsPZFkXHGIhiPfNhuojlVg0D5VwoIbCqo3zLgyBg/jWkhnc4guBBr
fx7gTgdPvu+I0ozEhIK3ZQ7DlGvwzwVxi6D+ZeblU3DnrRZ1h8HqTyUyGs/FtY/IrIq90TZeUzJL
TrVLlIOvrYUWf88cNpa8pApWNYmj9LK/15aexo1tX6l8XPEqG62t9hpExKM1e5qRCWCT7j5qbl0r
QIJBkqPalVcR+BfYB9bUsaFdiMG3GD0aH6s8LQXxaib8vh0rDOjbZGZ8hX9TWkqFk01QcdWopS+n
6kva0Qmv7EsR8txijh3FJ+6YzI5SqM9TAEV92DdZA50zXBRpUM2scz8Oz7ZENCt4MEGM7dWrtRiZ
/1WUp0qN5Rr6rD3tfHPd7PVX+CUodY72D4o+O6Z/5bzPj5eleQuGaVsDaxLxnQuEPU+XEevgfxvz
yP/iHSk8T8yBj6MlBioUOo+c5ADZDfZrghyQhcoBx9A1a6nW4VLT8AoX46qRwuSkSvE1NjFnXNyW
0odlI6Oby82GbnpX/ptvTFacJqnhB0NsVQ4PepEEzNI7zypIvEi4Db8ry+4qJdlmIm16gIKryhLL
+BdKqXQuulJm26yuAjiWm7+orNE6poRqD06hoth996tKdPvGX86syF62V+vUv458+kqEmniivqG3
VwdDK+aTP5+h23zG+1EaM8LEEudqeQsLLPWfjiRzqLRWDk1wueSN4BzCb8ZuntlC5OrSTPj1JiHJ
V3P9ULX61TGNmHKo7GEuENhJ4nmZCwAYjZZlm3vawnLXaOU6gr3nrwNVlkqWVgl+0/EVCOuGTlAP
n2YvjAc+MmaSdVqeRaTHsD32U9dfT9v3SGjujYtuZFsaA7Rp5fKrkTTRi3EptG6tNFSB5vCmE6ie
eG0JBHwhGwU5Q3gCHZOy00efkoIqPe1Y/Gexjd1JQJB7cKFYSef0kvvxCGdR3ThD40sBd4IoBjBe
kjLkkTiTJRx7uaBffaxJvXbLEOoveYp2AAsTMMfk6mD2ufgcDJpevj92oBbLf8nFLmlz4ZsgvHkp
tmgwgi/fseOSFW53F4dNq8NaNV1q5wDDGm4D6IEsM0CgOiT70U7r4F5x2ghhxnDfUcoALb38l5rE
PhQ3B7bHsOcTlTkI8ylVwwPLY2d/xurYt5ojFtsDcCG6MXDcI+UhfJTA3YUcUs6qWtqZOZ4Ln2RO
Fh3Qa+dPZVUHe09e9Ci6M7MxeuNBBqaKxI25bvy3IqOINeFTMkI8LXHz8VIIrg6LZi/hdeFL8XlU
8lrrR/e3rP4IYk7Ow9wiy1aQh6UEcqzezWcxCHfGw6dBKy0DkebK7YsLzWFPpxWLsrByefVOz2ds
41oVx9GW6a8lHdDZymxVXxni01M4TGXJr/xM9WE28Ukj5GX8deBJvZbKKUbNc/rUJGqaGhf4Y8V7
uCsdDOcRIFxQYEb3u/8BNxmELxybENb9tpolYuC1lTFQsOjyqbVcUHqgR1ItdsEvi0/nJw/tF23l
L6PVFSiyEmm0GBPF2BBBVeclFOugwFf8l1KCOQL5ul1s1fEFTSn6jyA1Oq6nD5PhBBTe3899n9Kf
oDyDlBLrKQ3FE3XYenbAB2rhfFOBfRnifF1ROIQqA9dccV3lOFH8EqnWODSJ8Qu9tMqSkVZ+9/C1
l66HMsWvrZxd3pYrPF8ep9p3glq/RNm8uJCxVUpTbmkli0rWpKp7VaS3RYLMwQwKPNUqs0fIcGFi
lgddk1JbwACEPHFqaLr5+7+zzZ598pQjKfMe1yE5zdHYlm5eocvzfvt20btMiWSME3sLr7eiOuLI
l8jGPr58dQNKfdsBe8eR7OwOD8PKBpEWvVt+6O5yN6bwVzvY0+xdGlZ8cWScJOOJDnrKMOZ6sP6c
WHlaeNtC0BpM6cXXs01pG2qW9agg2ZEFMx5tZliP5yvhtH47qCUwA7LCbcD6avftIFjY1BHkXla3
7MHz6wNZlTuBetehC9psdAG3IA7OchpIF7TQdBHXhij/f8x3k6KYQbS9YZNd7EKAJ+BsACJcz1Sa
GNKDVTFRSojarfVoUsTZ5KG7v0ADzI76I7pBffhOm7hr2TdeoLhUkOiZRoE/la9Q0dNg6w27gRRm
48VQOc571Wf9wgEwdvvLA5zivkT6FHKCjnRDeOK1h9b57vyu1mYwP00FILLMchNCwij7fGMDGoKN
b9dyfrOvg6i36W4qxmIZWlrwkW6/Qe8w8mZhevUOTsRlgCq4QSOTblzZZOrxCB7/Axp1XvYrbQqw
0XqHCSbQH7+PtMfMqbHwfKGaAMdyTshVKFgZdzExPF7v1MRKta+vQyJjv8om1B3C9U/kLx/Tb2bl
HabBRig83FNwunYyDfhbr1p9Tb3TFoM1rXTUPQzJlUtKe+MIJLP6I/94RUaeX1H1smcynsnvkii1
br8a6KBHYlTmG4/YzEsqhGH9lwiWGew/tk0ki3epdeYDz1LOUSvUzl0h18efhslamgUceX6cH+bk
OvUqkKQOlUOK2tLu++MUEhz6K5hL0NPCq9rD6ykZ/vXElu9gylNpSeE/yXqEBST0UdwQcCEXi605
fth6GvpxXeBhEHfh9tcyHWqq8afboW9bFcmZ32507xzvIhklc8R/qZAq47Sz8hydYbS4vrqU8lel
GEMtyCpA+1UlFhlBfndwA1E7YcHpqpKpYUpqUkL85YY/+Zt5Mkk55S4wI7gJ2lD84Y384xnf7+0y
l/W4tdCEZ/SxBL1tsF+ylgj6/D8QofMCnycyvHzAi4TL+BkruT2rmHAf/OO/EvgWzS+6rHp6DvNB
KSbiPJRzFgU+yr5/l6nl/guCsOJOMcuMxYvwCyBySuXdgKV6OjAui+tA90pw+7zslkiol8ArRSp4
JLTOiYgAmEtGnmKnawIbGscd8NtaFCAd9WyMRC9yRCRjhk5um3v+00sy+zB4L1VbB3XC+6ftUTdr
INRsdyMapyb4Z6R49T/T6bQ/LCk0AzboGzGbCfwtyjIQLdt54LikUpoKq0IX7+zEXhcMa6ungev6
6t4lJ5uePkFRkir+ZyKgaSoP4zwyzOxp4efd2UU8FeAsWScPNXTAUwMksPCNFcmblQvR1TNG46t7
vnlxctc3M3W0UN29BhxfczBftfX4g4ebhmY6iOvmApmk1tCJgglJWRHJCS1xpfehZw3L4QtzIlGe
zGg70dXurtO4jQ6eM/30ekXK/6kdwGu8YmQ53qiHzNftkU2efnWslxLfVC3Xoc7lspr3UkFzCaNI
pSmMp4KhrR6TVlDlfPpZCyun90r4/H46Lt5GXlBsE3mwGaBQCb4aWRrFN5W+zcN7/kkuYLN8arF/
Uf6ZM86P+4Nxw9ccPHjXm9a3wSJkZctxlvtrlBff7wFUif/anK4WWwddEEzXA9hWOCTTmoFQECc2
e36qmdBTNPjneuLJHIhYWNRVChH3iNYhJp4qI6WDwA+YyKp2/sFQjKZ33/UafiMzoQc/9pd2juDg
CJ78ECcUyUBjmMOnuYMOPRvucLxn3L4zV9NQ9zpncSVKmmQMzC5wydJremD4AR9Iuoc5jWdC4s3j
+Cj73EdoHnECwRxcn0BLsR44rTniamCi53mIhgp8QrVzSa4H0ONgBAn9aN67bBnif6uOguBHyF3K
EIP7+wkMXkxchteFoBNfSKnfj8Gd1agiguFFaeY3F3cMIrWAHCD1QYlYzBIkZQhey9OfnhpWjcXN
pPsAKMP5aqsBuIUF/x1bPAOimT30TkoYC37Tg6NSkkHzxiLl6u3WT46EpVuaMJzciOgs4Dqej0KL
WvVs3S7O+PNDdNf1quIIngSHmQgShku9bkcPRMIdn/hGt45/t/Tfn4Zxqpv4PwDyM9WyLnG33HDx
/IRwcTmghh9tmb3jmGZxqbTwGlFX2vJYcDtUAA16hNDCPIP84hTv5vuaH03GtCnZkKG2nQDZ4SbQ
ZcB+AqO9/NIxsdz5xZ1R6HR/4xua7rwRAE7wTqQvvkR8u5Xd657WcL2VvOU8E/8a4yBW3TOWTUHY
p1XBhKCeY7EyCgt4fyfo7nsrDSzgGxtkQROiEb+TIfVkd+JlfolaOM2YDf7TrNUwg+paNUcuyj8n
pSXCjfaWdsTHyauaiefAjGrnHV7klWFGOc67vggvKCOYSvV4BoZa71gshpbn/8bKwWQd/l53Q2HH
seyxjosqvOi5b9Ifdv+3O/n9E524B+LOKUCaIJTyzD+urBb3KqhN8Qzh/W5ehs/7fz4QCCjijJ9C
GTW/m7bJtokZi3lMf/QZEUrcHGIhtQ7jE9xsY9vd8aqgPf1JwnGGoMQoOpixsiI31AqKgaKC10hr
P9oblFkIsqf+gCoR601ThHrLbO4vLQLokohzdpsdlYTCqktwVcHR8FJ2sIcCWKgDWeHVioAN1LnF
TqFH0YReYNBhqxTbxXTXkn52EUM0R2Z5lnJ33tpJIZSlHABmtPsfJi+BAZM+RWucTSw+5YDEM806
1akRch4MwCxOyXUJjpaMpttNvRBSaa/1MP/zHtzGDT+CHdScEcDUBWeqGW/MKz2PsSig0Ntm2TfK
acsWoXnLqhb02c7SYXzKU5YL30CBltGbxWz6EbOgtt59hMt5bAcnRYAvstOGGETh6q8aLONUDY2k
ocyB/Gmk8GcXXfJUYpjX2FgFyT+/MiJvdqOZLaUPhYSyoU5pxdYUSnN9WVOUrShKGYwqINoBEtMo
ILYyYdsJpQ21aGdAXoC1Bojks5L4rgUUK7YICeAbSU4tBPSMF15r3Lz3LvjCzwm0Z8iLUwSERhsY
T49Qrf2GQ7fJBWZcJxjAsoo1FeZiIYgaxuF9Dvcnz5eNdeVb/lX1VDnp4a8atkvDmOe+fN8UjO3S
UWxtqIvlDwu7Gq/zDbgpGWhRuN445djzee2UF3M77ini2BPSObMkNfX8bT483R58llfQVaI42qpu
UxJJ+OhjubOzRBUu+KZE52OPmVYB2cpFkRGI5XGHsUKL3R7QGcZkDUzM0kSAPty8CUDH60NY+oue
VMAEWS1egl3zkP0+ZH2SzjoVbeFEE0Kj6IbKURwWIBDzkf5RhkVK6i127xPXi4itHI2JOeR1nIHr
8HZ/MmB0B53GK17Rj9u/FPz+s8S4zNYNIpp9er/p9clsLuHKiKtpdp6IYRoYudUmBxogdWG3AUn9
QXR+oaVMxGw2PhGYnoj+569NZ89t6ynryCUuPiKrcpuZnrTOJB+ghN2NRZFAMq8m2n5T07cfU9Kz
s9yAJuS1cv9njABp11OKOm56VT4mehTVvchEn2x5YFa6ydtG5vZ9znSHY1NjdIqqcpd5cWQNg2Qe
gkJ/ska1STEUAxL+czr2fN3EZFN8VJiqfgCU+cNs7CuiWQ3pK9KwT39a+q1l7IY8beq6oaIf23zW
bJjcDC/DQbTlLPt1hD3U08/M+kO3p1oJle7HZI5IVde2msduY1WGnzwz3ncjETRso9Hp1+UyAZ+a
lc8LPgIPJeemt7583p2WuSI38shQ7yRl7bt5mSRf75J5loBBMc3jA1CUhUimo7+889ptSlaprEoT
ljOFwY49xvQ/Ui4B6hkbznqWPnf5fdKnEDM6N78SwM8ItLsMK7i9fM/exJQth10Xe6bEvJt3uVvK
8H2XiBqzhRYnhkcXRy5ej+WUQuG4XxILWFVH7S6Vb/xBt8ViBDcniWXdSvxiPjpEVidJnrYzPln3
LGIZZFxqU+w5Q1CDqa8BSojlp5v+d4cv286DQ/0jYY+jBgKoHaViYIh72+f0shDJpksAvEGE+PlA
0yoJlt7FgHOI6j1tbsJGSEOi+vpaSRNRyo79tDriI7Wj5ZQnkKnlXJI67zw0Ag+Zp4nbotjl3eg3
munN4DDLr3J6phNsROnqsGzRgQakY5Deh1j0+hEYtm9FT3/Pjm69VvE9kSX/jfpIjwUn6qZ+1eHs
TV1wm1tvPgZ+mv4yzR24PBnEEA+hLf5nwQ57BX1f5FS0GvRb1QfzLiWHGXKQuhxYB/4Cypr+1Cep
a0HxWMoOaGn0RAKi6zMzCqO+96EvCII5KHI1njAs9YXR+Yos6fKupIx5Up1sBbKPpIsUVrb5OzON
nylCg5BdAllzHgcrskQvC4WF4p+u62Csz4QYqgoXQbbnWm3/GH4ArQIMKGprLtXNLh1caknUBd6n
3lnp+4phVSEiHuZOD97s9npCkHY4/Kw34EVdLX8QfX+W0XGhK3FNiq5fFubE7pO3GJVsAvAhwSdI
bjxuTrBPjJL9TSOFUIjZoLJE1/ObER9IiDKVQ1WPOxdb3SMvEweOyAUN8AX1cc0j9MTUnYJwRfzM
jhQaRolVTuHwHIlCHXOS7R4gUJC07YJcNMqqycPL1TAig2Di6tBNX0v/4Du/Mb8VMhn3Dkjn7Px2
5XI525UGoBxoDRq0zPKwJkgAyIt13Y4XP4f2ENNu2BF1ECgBqBqT/H34XTYk9GWoyjZ/CoSURaDS
mZKqG/1vEqmE3OuAHCH9zCqlCqjpp8QKs6CzVnzflrNqehgXUzsuWX+m30IlhvwkxLTE2MWQzzJI
oNuxSa6ZaCvm12znCzSEYPDs/1bdkK5Pdv7Ehx7SZe8lSYHXFtqU8vqPhm9u+ifk+bAhm1eBh+Or
f6QQcBXZyfRO45h3YQE3Y9UoVSCOnspFpek5HLy+KJORchXp907LIWskg1HHKEg4uC7CkhgHkVPe
iE01LraATAgLXruokkXhOR9OuWpujmzVY1/xyu3nodQgdRP5Frfe4tUN8Oe59iYOqDjm1l2oOT7W
36mQBBwkT8bLFNn4XaUhxSCmxiNRhJ3IySiDcsmJXRFotXQqFyu796qY/1/3nD65/vrbNL2l+D/5
+i6gNjK/aX2ck/MJvWZlDA2G/766gDWxYVwKzIUtM2pzsqovv44SZb1yfvzn3VZ37DHNzbuqTPWU
le/MQoZYJF3UrL/XJOGSSQsGXWfqHaTOK5TLDz/y1vWondSUlXZ1kX9DOzKgwkyj/HlQzT035rnu
BXnPLagLRe5+rTdZOpgOwyVzHxwVV45CssVNcQgin8XnFmsU5wzTdWxiIYcNc8WxedBMbJZegGJI
fEVQCtl+rNtQ/ft0M9Ij6RQFMKvJ1fRDrGTtumDn1nrFNKeC6Iq4Rr/juXYilkUk3EzGlkagqr0T
ih9GpPcR8NcASPMHJ38wNbusk/Qg+A7A8V+KRP54nKgX9PUF8qNUGtcrnvUkYt1+5lghmGesyZyJ
ftyxElFes1dRxj9XCe7VtB9QxOYKFgbu5BWrIdtqbX4vQ1dQTtb4t2tlMj7M8P7oXdYLAtC3a8X2
FaFV2N7ifPB+NHrZ0rKohrbxVktXZlXLll0h9Nhd1zqA8XJoNA+Ge6JV/P6fhREVZv6ZHJSkfzWX
qCupeias9GXXmsc20sqM+Dkf4ru/F+DVNGT8a7Ug1flmdaTfOrK/5L/8viCrq2ctAezIMWdMpc9N
CQnNp2lfUHns6h4lZ+29poUbfUUv3/2JzAIl4XZvyNQSag9vRCqjMkMNh+KWW/PryIm7UlKqNQka
frm2Rknc+FNZ2alG5+zBstdkxDVMmfDhO2JJ1KynPw0Yh3HxLN02W86czxU/BX9z5ncSTuZeyNNI
78HHiisFjFyuCYT90G9NxJuEjNGLM9QzK9UdNlUHGexawMxY4bmkcAeNzhjFlUNJ9Q7Ul+3TjVuO
iAQr/HATvxNSIECK0RUCqoPYHplhQcp99r8Y2QFswbeF5zdybOkhrmp7QLAPE3Jz/hduyPXJL1J5
Va+zK2IGMNv4lJvOEYtMsEHashGwZ8P3tu0DgGRaVv54auqz25R0XkFgsNONTjgrZpZN2JdqxMn1
JopLYEimgUxygso1YJCqVxKIIz39WoK+UBNIeQjq61fcA/xcZCoxGZwKzbeBVDwK13I+1gtsWXpR
xtyryKljzT17zp5BrUW7K4YgodrfIngYrMyOxhDdZApRLkhjSMbT2hyATKhww4Gy6s/ClvCtc37B
GQlw4kaBe4GLQRDd/Eu+sRezsClRzfbCZyDUMPrlO2a+n/+3hAV1afB1HPZaTO9QGql2YuRrXeVG
NSAzo79YQMdbJxAFZ/IqR/N0+6wkhHQkBkRPHMUzhGPfEF3Z6fHHYvt+vh+wkdBQaOd6tjJzV10d
ShryRMGMU6cGi3edWmuYvfbqJQ1JAPXfCF7wdX5puH26VoT5nB8A2SuKhRIwzdM77epgoQHNLKHZ
Js2FW4XOJocwcujlsB6eo3U6HkBel8m5SZsaYEeM7YLv/3s6AJudnOb3MTvgSBQIV+wIl7P8ZXKK
1s0cpvoUA5sJD5nmFU2URxecL8HPjF/OhXi89GYKEaVvHjq0dN6APgATAUEmukXQrcmOJmDSZcbQ
4eW2mPZFPCjxl59qPy3moMk/fzPgj0G8lIW4Wfws+MB5thENMKq7nsXNYv43dKygBXSWdththcbo
xnj1/jNJniN3wB0rpcDju8IH1BxSC/5PrjC0BUrGoSGpVx+5zE8/+5skiZ+hqFcjLKWLwwk2SfS7
rthfCgjyNnNQYljEHA7imWOf/DO8YYvXrCZ2QQCgxqkTvH9bybUk6MbMjxfXBkOGkUjcm2izCmoV
UmYH0wMffp61E29oToUYUFjEM0c1nmJRANGFnD9gx0ujYb2D5A030+u+vgmI3O/XmzerAB0ZHetS
+1lzFHeqP6tKI6zJFP9zlz+R65qh8ZbionP44gANci9a+fESiRn0z76aCNioGsZpFimBZXgJVH90
XRPMB7eZkd4rfV8pfNgr9r6sxg9Yf4OtiazTU1cbvWCVbarxf4hAO0GmUZSNJcDYsKwvxczYIA4T
iCitm+e0wz2mZ2ruBPoGXegti9tsed4C2OYSSehxlDFVgjBU3XNRe0iTOl5cYjStc2oH/8mEBWgx
Hy0c6Wp3U1ATdsh/nVlhBhZQMBOETvSFQMugloODAlwA3ZqeBadi0/VbSpVrMywUfXWI53L0rq3U
1LsGSTcdUOEx8epxNK8YgylR5FYUs8giClav6Xbq7ZkfZuINBSlUnH4NPDSK80hdctEpH+WZKac2
dtOwG7eqWHQ4vbwCqOV/6qSSen4oKv/q3g8OJZZrJvF3moPGc2P8lDXEKy0mnqAmP/HbfGN/MtCk
v8jEIQrKdRT/M4esjSmf3/SdSCDzHTm1fkoiH69o+8zmnStvtVrnRrp+hdIeuHBaCbodQG8rKj90
CAKa+B7C9NpAoUTZ59DlXbvewHmr89SHDln9ogpWTUBK+S3xvSRlkOUhQegTLCbOKff6pYSwMWOr
Oh99/69mKemy/zN5sf7K26nTVGbary4Ko9vA67FM7MMlR7aZcvJgmnRU9RTxam/z9yKCebk1ff6w
s50mWe5YR6xwWquufHAgXRwSu63IFZoMlV78JOonWeXlgASZNx3i5PzYO00Cv+l5PiPAENUm4Jmg
vnv27x3F7tiA4p/OhFBFCkeHkN866JFO7Zg0R8pOc2rw19WtmzBeRgSWoy1OVTYgcLc2VB6ZWLyT
sZBwHlpqaO204Hxqw4zeSLiY6BuWecQlQHrd9sq8rxME0+v32iZ+gFyeajltNlLcXCNx4Ovt7ZqD
dCLtLroAUpeoZktCiloGeTSVyk/fV0vMwJ9Q++3Fs2l4P0JmTXU+i0pnAmRq3fjNJWxXkg7cRRNL
b9zLsoArBdtcGVWV5PPfxuOi0yNu617FwPaGeXykRk0sLPLYd27VY0p6L18ePfe1QY50OiOKxS6p
RN7HJzkW6HXOSsABDMHaIwX5/76S63un/YWqOMIzPDMcPsuDymt30sLQkHQ3W7L2tVVmhG4rq5jn
9NMVz5ucJx8qDZ6q4wHuNANzLERxFZ78Bp1t/fUqY1AmcajlV7B5V3psCcMBIUNDfvnB6q72cK8h
Um5sjI8UpA/6IO/pSGo4x7pvAxs+whnVn8u1MRjfas63KGYE8lzLqZa8EF26rf3B07I2aSuq+p3O
BqsuiWImVn1PtPfBSJ4A026Rhw3BYL6OmfHAOkR/ntjiasbUwRP22uYYMHNtAaK0aLBz06Zon+8r
Nh9A/Hj+MBvmEeuiJmf85r/TASczMPxijrMRn5FRalpCLqOK069/PnRczdFj0RbR2WDYlKGN+/BE
gPCqcBXoPyNRw/pk2+cBQhS6BXUuuRhuDegHb+CT+KVmF1iW2puYeKpabyFWrWWcZXUczr3a+YvE
PhBS9KwUrL7dx9zpRnZ2gToGYpFTG50TqIMVotegpb0z0tn3lL9mH0AiiVzFxzgUhk/ySjdP01qI
+4CDEeA431RZV5ZSVuZ59YOBTj6spC8ArbZOFRVO5ee0VK5fL45D2RioyQGZ5QOb7+bUHpARAx7E
6mNE2dCxOJ1wExPTs0La30jIGpe7WpItpEHjXhvyItWABmhTZBbA+pX8nHtMuKCO8EjoioOG75+l
fl6fPb5/u8X0varcozxeN5zpVOPEwQOQLA9UAAHJnbelD9vEUh+sh/6jr/yamyBBawHZXvevXrJ1
KhEh+UFybzWxMvm4CTdslMgIrBqophi5EZ7lUqhU0Rr767yNNbW3NBNpX+BzVYM8E2dj7Ckk3F06
zvr+W7zh/mi+FL6buSz/OJpPjDYlw5JYFDNk55K+fOVOLX6+7Qo0nCjMQ5B4YFYXI1mS1U+6HEzF
6BKnuCWyG/gR4M1brhz0cv/4SMFFjMVssm7gvERnD2eQNzv4EJIkA41UXNXKX6MyY3TtPGquNamz
9+pQQH6lVj8YamQZwjqAfCa60UQ+d2KQZ4ZS+I6zb/buQSZa5dPn3ubclkUa5oJuqpZaduEb3DYT
wAy3QTEef03gw09Ze0OCzoArzZUiA1MihYd2c2E7+nAqcKeogZ1Vj/G1HGbuqhsCC+EwgbIK7509
klXG6GlHebyTDqYbLOIg80adJdVTgap30LJ1AIbzPfcLW9abLUFK6B/7swjyEt3mI0Or2am8LL7c
5KoiOZxOlD3l20YeN7PHuUrlfAztDoSUO8qkgi8dmaWuyIMlN5lJ86wNdRE8OE5xGDjzg/h14WZx
/oJzdfBjkwiHjJVDRW36GBLpSamfCeccjbH+V6ixR6OjI7AvWk25JgIsR9QepnbQyRR0joRPyn5D
Za6GwdOSd/tTtUCN3Bc3aM/qGkhQiJKAOl2bHkKYS7wMxylPJAd4IcyShvXTBaJnlyHWA4XP0ug3
zHEIQXSQrEg+Im4NX7EHAAYZmsyKsaUQAPJ3v8qPn8Shw32J5z3poGD98zs9FRItsQ+5ZL41ckpV
QO17/jmecox9ThdEiqbk/n2f/JEmvoK4Oue7bCLu+WieIoPdV3Nm9jJSzGULPN8YPevGs8fqd1q2
7gXoLMRGLUITHkMjUqb1y9vDuva5OnJPb7NFknbnur1FCnL/PMEwJoixKJukl406+wwLa9wYFOQW
OBkTU1iMX5/munjkpQ5/5/4jBWnbtzDNr6XFjYawOPEU7+6qRrDRnWckUCZjoqStfQr/pCJcRQ7j
n2BRMnBXCKZbUJSEzrtKLsXA/luGOq4p0euTtvbd15Cm2BnS6ovOo7U2Vy2ihCvu6/mdhkKqp62o
tf1IxwiGWZ0b1l9CD/AfU2kReJ6DSSrilwp8FdHe8C6UCFQehZ4923ZictEE+rFBsGIy9ALqbfyZ
Ru8Ll4AjmMTQn3bS0/z9x9Z5a96S2HfGM40jIo5C7OANuSCfLF42rThM2mrnxa7OHvEH3CoYPavF
Hqro07/6XZsvD87r6DgB1S85uI9IVB21vZMNKXlY6u7k6Me2CIYt8GF8AOZiXaiUqvni0VN3TJA5
zEKld9tUCNm2D7hcrNIdJIvZpBPaBZ0nklRWat86HDaclmXxMRVBLTR2DzuGq7iimWXIw4+nE79D
tE/bgVtqv9hAYxOgs/BTQqGEqsNVQXf0OT5vq6CliGkrqycwOguh+Sr+ayZZJRz6PUmAtyv9Yh9x
8eF9MKrjzV/T+kKhIaoxJ/1mxAc1W0Yi9cU9LZL78aq9yuol4cE+KqJPp5HWIJGUT5AWGfQYFt1L
UZeP1eMh8IYCNTjxYgec+kAJ2+/cXXFUilrkzR19P02+FbWKPoPKPrRR6R2MhdkDHn9k9iwBK6oW
0X1YEL3X8fF3s0DLxNZov4BbxnaPi6yw6nNGtJKWtG42TpYIQC2sHCrOiUnJSHz/XhqWfIJP4VBZ
CW2sH2qBlPHBxc2vPxUrcED2XZOlCmsYoHjYn7DmveTAfCLV55fGw+A2Uk3oYzqzg/KtQeeHStmG
ApPhgXSlytHKRfojz5ug9UCzVVdyA7GS8T5rXwfGnNZpkO4ilVoSc+A9A+ttyeefvxPts83hqw88
Yn7AT1r8phx6NC4vN1tWxB1+ODFYDJew+do/R125MNbEJhpnDNRKTkUCu1qngvwIUZqKDxY588zv
Xfq6+ydShvNps4V0kdaD6iIb9kJQaM2Td9Qfeg43A/6shy/ZqCpqduAoVO8g3OwiBW1cfGJBfwOu
EkM/8gCOl/Bfn1Na/3AsP/IlcFXjpWI35/0tyytQDDAa4jNt67yuRf9GyGxcq6T+cqXq5Jp2Jxa7
CPDHsldom/Q3GNdzICrj6vMJyYADGkUdUUeUqKsTPBbC5XBO1l4m8pfVczsalnLRcezqTvdygeQp
Uy0SUEzQMn/SNLtnjibVWgXnCexg+uK1yEYGJnTxzPatd3Ci9aFJZC2wnhxVVXJTI3gfLzqxfu87
GMH+ZGQk6MPe9QK9rXg2dxU+DMiRZNMPWweVXJkXlwIuKJu+YUb1kXnnil9H1jDkmSxB6/rYSiUE
Gjamuw8J6+pBzF0zhEAkVBDbhEZf0wWlWoVyB2sufxNDq1w9gX4vzDtcNJ1HXY7mNXSWkMSUj59f
AWvOH3NhAtM01kKzD3mKnOPKuGUjTi/y34sizU2snF/AUiwdSkTQ7PBDhgsdIupncQV5GLrlT9Jd
63+oRQM9Yd/r2SzsVRmlJygP6gDiNATwXZkMPip9K3OP7eLoiyEHRQU1BNQ2KJW0lTN6ldFWMh7/
4ghCiSJiSzy8EE/EkbrEh1AxX8IOfMM+/LCIfwedv7wJ+zkW/3CnSbUMLir9hhWLl0BuzUnQH6nr
k+wY32FapFxCVhTUW3pVUCL1xlOl/qlFuEApoXvU3In5wn2kzQxuvPVMltZdcCjQyWV2lEpxRAhE
h74HAm5H7jKeLuCnYXqBQL7/lSGmi5fgS6Jj0M89rf3sAMLQ95cEYrXqfrzGWQVrYLY1xtcfSlzx
/I5L3y66YGItMhE4+yB1XrijHE+5ZtH2h2frZqoC9Nuk1W0pMAqqzPuobbGbK2VxOCFaoQTTgb+n
xuXE9xWUSaeJEfrg3kyyn06uXyqsDq37iR09jMyELAj7mg5SJInHvR/BgTQQ7ZpRDOrTaF0z+ITz
Ru8qVDFVNA6RFgPtjCNsHozgIgfi/qPEkSXBjG9Y40Cg/QkzCr+BN3JoIKpi7b5jrhyxQc6fJSmw
geiWIJkaqbKo1qUEyQQzCwWX2zzoidqIZfellqvrDVeXS7HmnjCZY9nUpz0oHlGQXphMKArfbJhM
atvMJLEznPrcbkIMTZR6wjlqCUyv4NTJXxUtA0o6Ol/LPsu7rUrWXDTnTRNNcnfMQFdqPabb0Xwq
aiSCyTGDTHMb8zFjgvHU7j5H18j9l+Ak6UOsqpcrIVwYFPx3X5/SWbna47gjPzF2t3kCVOcA1E3b
A3W3tLRCEIfNCI/wFicuVrAuXnD64YRy1PMGwOO39VhNMbXRXkqQlvjTz4IjtEc76q4U6ZbgsWiA
waAN3itev5Qq1KTv/7s07MJPEztAQ6oJ5s5n68H0OkKU7o+KWztM08Zmxn5eg5XcpB/aLZDFT/0T
NZ0RAhdKw26QaQnpPRMyq0mkfns3wjF4h5W2taRQTlipxDoMSrP/3pzGmSdppLHmS/yujFting+e
gTXmX2ybkXd6tWs8REk4syJZIeRtKITX0m/NSBpJIDCi+Hy8EQ14fjRIQZuYq4gGCtX6DItUaQfV
A1fwKOmuTGJsclYQkt8mC3BVaKFlwrl4RjbC3nTekEJzXKQOHRURaquX1QGI4IFWso6soyevYVSf
eQGQwCmyfLpuQOfblkGkzXaZc3Na1fOCR8ddKaXNVsliWtIZyDp9XtKB8VPv5DVVcysKJNDZ/WtL
KXqe0rPb1Na+dCJep4bvtUkqXpdehotwkbEv9Nq0qK40gMUYLTVK2pKeOe18MD8B8gyw5cg+L32F
YnOJ9d5CLjFifhtLqwW29zg0OV2i8vdpkvsZMxpIN5fo+sNJhfWeiAMuB9pLVobmWLaxsb6Xl4Ui
z/KsOG8g1LhkJ+SL9r4/1UCHydiB3WoLQdSW1YAV/lGmyYdr5DFyuB60kg50eZT0f/bPrKemtmFw
4GKsqsu7Z4m7YaDTjc0A82Gzwl/tsCJsbEJZVOCM2lp1ndt33r6q+SeTgwU2R0YJn2yHv1R1WU9I
iMCSQ3F1RlOI/7quHXT3Ketael9niEZvlf4lRWRsODh3oSM7aMuLNedkGUdFlQDv3/pO+ctEaJvZ
jK3LqOGmJiXkr6gQeBiPNFNG7ngpjlSsJAfvxy6NcDWGpedxMdFKBuOzj4PErQtqmYEiU2srqX3H
MGTsZW4GQj8V7qguczKxQgLmJYU1U4XMgi3mSk3002OXOsrGDbSYgznGTQMMYfnUfdqyrsYpjTzk
enM2cVqHan7KMfSDQwVefS9rkQqIC8rlFzvMqCsDk85arMboJpfNj+Oc64quWuSPRqjlVCqGgpN/
+MYtvMLIkDNPkuahI9oLl6BgHk2gl00e/9afQ8sBuzKwozDQ+iIXkfaBv14kUsDD5m1UHf21U5TB
xaAZqe5bb9aCuzPdR1MUgBRvmVk7IQq5c5t34gwBxNmsDMwZj2lv1i/N5EwGH831JnCe4TBGnULM
p8eqmXzFLqE/lFC3/IDmrNOsokYZTG5gKga99kqfYm9Ak1/fplDXzryfczGYtnkPrENtaiKHs6Fk
2+B8b/FrOEI5d6hmpIus/iyuxm1oeKOpGVCUhJLfFeyeSWFDEqF5YXQ+JAEcDsP5JYDBrmCIVaAc
RqyvDBpTKUHU3n140DN/BdeynhDq757XyS3NiM5Hpt9UQhCOSpggf9Zhgq0j112uaPP+hJCyPndX
g88n5xerji5/6dvFdAtMg97keSCxf9PJt9j6sckQ+nZWHYI4Xn7T+abjGrPspqG/AgrwKAEZPzNP
Ro3PvIc1k70gublPakywR/cMBsVU7yZmQ4XYlcf4QHRwIVFxQM349YH4TBBlAPIIxWdPZDY5Lxd4
cWXtmzSJkQbq9Vf9OOvPq5oFhtKOGaf5aUm6ojSggRzJqZFe1hd/j7KmYDh9O2dLhVeAg6xZh/Mp
aWr0ahze9BxCyhgZ2lt71Q+hhRPsg1yktp5cWVw/AhcrauoOrBie3TnoSTQs6z1l5vLBR7fzimM1
5VM7X5KraDgc9Bm2jaemicLDh0fpzizCfuw0vweYAZ8NgJN0RK8YiTNDZ0Dc9tlu3HrTFdmRv74K
oLw29GDY7OJ92yAfh9jvIRwzbcF5b8NOPoJnJRAZR+tvdOmmJFR3tiCO/ZDwg24Qiyn5uGFpQr2X
ICUPthW2pxtwfQpcUereoX2y2gNWu78ox1DuesillkDh6gZcQQDHzRqYBxge0eF2lO9c2+UPhyYw
B/oxYsEoCMJwUlnFlH/i7bZvqxlc+F/5tFGEn02K6B/wiTdcgj0MnVSIFrDo2kXQNLG1kSApsMkL
k4ovDhsYqwDy5tiWmFnLywBVuGxCnzRc2Q4dafMNsJX8a8Qq1RsI6njW2DuTaqbmgedNNXwIHBoA
y02wx7K0rH9DYetAi8uvPCWiZQQTvjiO5xZNRwyjCktSgUUoAdlO/EDWeI9ew2XcpKwpyXCNiOJL
YLvur5OHaOScjPQs2PP09/xLtiMdirsNfv4hJmc0i8b2JDolovr8d/16MQqajkH9wJUsilR6Ez28
JHwXouKELl9Vkpd2MoKvKPIUPnTnxLy7NRgWKYYQOV4siUMgcDtnAt90bVfIQSpwZ2kZqM4KtzZq
q3cbgUGAvrgwyF4tZigC/66sJD0+gFEEzWh81Xir0ravA1rIG7l8mO9MNzoL2PsmhUSquMvUoq4e
/W4Z23C5l8DwS8Z9r+7n0Ei3nkmeZ5XzvrF2tSALbGGQ4mlj4TIvDP9onhnl9FlG4YwH1xpGjjck
F8hY5gGqX5V+LAWqbm0+pUuzq1eIycXgC5pvEnQjIEE6jDT8DQkVeagNGNWJcOmpQ1g5RGsyw/3X
3cykOLaKDESclD2BPH+qaYmZVttsPjhe2DYYgAaiysLpLMxprXx6hhyMoR2LVd7G9sXMwxbR0V9N
b3O0XAqCDrfo51NpGj2youdD6GbTgNP9J2F/IQDuxthdmvpnsYSeDI04TUPC8nVnpxJRpi+icurU
LmbvFOy+q2YcbKRLY1qmDlOtJ/5wTpIyJqiTqGsmD19RQ8GmRVcyDGwoh6a4B2OjREQf/k1DAxLv
OdyUX7WPRn63bgfszmdoBNavRVFUXo3QBof5x9TetHc435T6avpFC8lZFm/fTna9Gtk0ktlrpH+F
q6RD+ibmT2R/hgAls9epS62b4yBwgyKkoen+sfD8KOWjugSI3eRbv+QAAQDzw5HYSOBb+lVxQAG3
JVGfUpgHs8k0+itufLnoZczYZB73Ctm7RkYKxWaTyYy0NyjtbDwmDkXPEs4lEf9ylhdcsXDCxHis
44sKyjpjL7fkD70GREuhj/CpbHvhNpharAqlt7HHNLpJ991pYCxlr3MIJ6ZKPsSX9/IJbk2PmsqX
5iTxv1hvDB01lKHwztW/JOmUD38k+Xbz7ctB0vl+SURKYGjJBPo2MlSU2k5IbXbVEaZNgWfV7X/0
KAxGHMyV93JDiTQz6oPf90kXx0D+t/z083mhU860SNggwcre0xiGyafvOxbCNws/SsQFeEzX1/o8
xUzcKSqC7Tc10Yq/BmpWX9jtwE5SV4hi5Pod3nlH+IdZWH13+aeXvb40FEb25PbLt78AN49CwpXn
Tv0YbgtbMeNx1fADTD67ftffgzeAeFCUQunuaMWSHzVpzDiUJPkJx9Kzs+atT8ILiflI53nBH+85
YVqABq2KX1NoTO504AelWlNDm20Nn0HoKwFB+7sB9++ut7XNJ+rkt43O0gSmEG9SqYj7qNHr6EAs
uALWNmimZKon4OWqFt1h3aBHFYuWsFgjY749jH6n9hD6iHh+kNJlySpJdYck5ffwxX/u80ESGHQs
qOSrSy1LipXZrMCrVlgxZNzagUR9pRIfbHa9odxvSqAGk0H6zHkixNRhFY7lViQ0oB4DjGKkuz9M
n4uu1MeXMgJGPjvMPZqFbvrZSlzxZ7jEzjM2L5WG1l67EJSmd+hVXrScgpmUztx01QbuY60+Lj1w
MheiyPmCH/55mC2YhTuPcrk2Rp9egxLNmW+hN2AL9PnpWYRK/XuBFE8pKa+hDOKh/KBqubpR3T7X
BrgGdnZfUyOXYO9+7J0Z04itOueFu7fqVJAFq7hMOsCjSWSGK3ls86j/jDp024a8MBfXFDsW9Llv
ZepyKuHNhR6OnbDZMf1bru3TcZ7EsO3wq0tmdJg+wWoO4X2X2ZD9C2H4e0Hjd1Ev5MTaHeTpMRlK
+IoecFVzoxe3myBPifPj7XftFemBb+8SPixRgWTC05uXgxnG0YIiVRiPAgKpwbMnTvFMMElGCStm
xNYahVTaCMqv9HlTXdU283afCwOLL3wm3ZPznbZh7UCvAsusYPPvreyhfExeIc+5LHgtQ6ZEuBoR
HGkW6bBECTjZ17jAZxsy1t+LNycJx3A7WOqdscUGBksXV4X0hOn7wDu7irrFfEwr35DzAiIzZ3x1
DaiVg0nGIpmTt5zgxbbD6l2PmLBrlt+y1e12EL1axuPZTV0kLe51JfnMoSWAAG3u7HFYbSHM9Y0g
zIPk/kHaX0PGmsXDN9i4nNMMBDupnV/BBHRYN2iX1oKAtUz8usNR44NlUjzA0YFQSm4l3g5Jp0oc
yZ9vtI1v/9fULzhUB8PdS0lwLBhoXz+hd32H2X+nFWOy4YBTsHfMs0d2iDRHHLoWZm/xvmoc2Xpj
3xSG/5JBGkT3TDcxYXsHQ6zs0KDsTBJ69bjceZT2KGilqM0oGQ8rW6McRnEB1z1p2skCSmk0hCUt
vrmFG84D4nIwi7TKrg7hvwCYS5wm32ys+62bfHAoQUu5a2zIZsNlkSxlik3to99hMP9uaqvrnSnh
uxt5dSQBUQn7wxytjDNXCqZgVaHnee7C3314v4otCBeAJ5dGHtOvGtZ5/uH0rq6CIixAmcZazI3f
DDn3iI9mqB8CoR9in0Gj3PveKPnM6PS3ko08HaqPynuTgRc8xHoaGWXOh579C+pC5MUF1QTYERie
dJcViUgebMeFHrmsZFYDzhbTlNXtzBU60FaPx5PHv+50AsWTGkAJmM2F/oW8pBMBZNgcrQg9k5NK
ksn4cEL0IczYnk2GEXZ6cDE9r2HU1+e0csVKPUDu8HJMVbAFvtlbXZc2lGV5G0qIeQdKYsDGQDmd
1dObX1d9L0gr+RvVyBtJLaCQJ9fVxqIbJiM+W+O3hOU88OlSBcKFdgEVhzo73LJkklXkhx0ca3JS
E8cBRX/VG+CwO+lziECkYQ6qa/JCJXMQUXxu911jjOPi4V0DXFFXjgXdgs2xZOaDqOYf00UgCVGI
fmlIzlVDs0ujC+pW6eBtwg5e0fmH7J+gVcANwieEnXX6OOzCwtNlxIwAnMvdKQcY/g1bAOyeC3qe
15kFIFbaNe9rnoSFCUoo1qUJiOabWmZYlGkAI5x7SIItBdYQQ0Wy1zc4ePCsl24e8FMZlWf86cj2
qOn+78F3tWdLrq7IlaROvrT+m6NsTWJXcwFcG1c6cArBsEYM2c053KrGfNdfjltSyQ/6ePGw9Q8P
JRWtC4BxtRqON3su1Ka/geU0bx5mmaT9ivpGCAD+mjBcqxhHQC7TVZndRaByKR++eHCS4SAXtSYZ
/qxHsxQAY34OaeF7ECxuEvPsDcQp2X3rN+k3wX/K/F+yWVTzQjraT7l2+GM9Vu5ktxRxP/8VghGu
hEkPb0VnNFw/9e28cYaUACCB0AjXoCR6gLcv+AjXsgTjrwLrcJXUn4pgeoKgy/lWLmUOopu4PrpC
0FpmLZAYTQa+LaoF8Ma/2SQaZR/AnG6iHWlq7Lqj+eGICWBwS10Sil+OQLmaeKmnbtquZn3V7AF2
fOnfQq9jLPyvfIwh8bTfvEtnPE7Wy8aOH/TjeI1HU0+xxRcGRyvk3Ov0KtCedvOqA05dgAK+z1Ka
XQDQGaLN3dmdLdfW7nw/RziFnyAotlZhB1HPGwXCQKiYun8Z0cQ4Wsf9XBhUbGVnvLvItrt5eKp4
hFZa7pmM9+JSh8NzPqN9di1K0J5fR4UbcjCSvwDemTE4uSJ+OMvOwHj2ZB4waA06lDrhGxi6KDs/
7DPttfjwj/kQE0l/Ze2hELKFY7OTXNKQDBTC15FfQqas90GEIfCOI5uGZAqqlVJrtjrGRr8Y7/Yj
GPDppVU+eSL3BZ+j+7AggoG9RFM++CZJODtDTIfkCw8abJkiCM38MFuzWJbVFOlwmdzi0pNoLiXG
tkk+fEnWozQOKLXqg15cTHMRhs21cg27juodGSkXA4KylXbAg5oGWlodhZYcj3WSsWQIelfAX9E5
3a7sRwu3RsOiRtqPnEvqw/Ci0eO0HL6Ie9tGuvaFY/DmXZcozNnjvwg2QFPX/wCyc82OyTsRjX5F
s1Fnx1+RtopMXv6K0gbmb600Nj5XeeaYci9+dUBWwCTQsvKpXs9JqQNlgdNv3NiSZHneBoOakMfa
fuXesYgdyhvp0bN71Yv9sz7SMi5r4GLIafuw3bCPaKmx1ziBADI1qS7BtJ+MwPNHe9yimCPWhNI+
0GyvGkq9pVme941kAIx1vLhkBbuik+kbzN0zRssXdL8H5BGJKZZHH5u5Mc46KznHqj9Cw73V87Cl
E3NIPEIj5N7U3m9sLH2bjehsUjocKwW3HVazsFE7bUWpaYKI7gY+Ww5T/jXiSvT35U1kM01s+ftd
9vf2SrI/s2WGN3lYNynLd4joQxNPBw9j40m720LHdr3gou3WmYBiSppGi71B1oJqB2k9619P3ol1
v+r61RPxKCBOtwjq4gbLBWNWDS5KVTCLaw5bERbKZTHz9hI1c+b+lHH1E/E+ASkOyUPltAkaVY9R
OLS+5iKtxN4MiTgGvvfaMwsk20bav48SqESKPtw2tAhqVcg5/knMDU+D2jNfFKvqw3TGBAsJnrxi
/yvKLdtTunM8jqykZUZ3lKBKSqeekH+5vpZmzqxZrzlGlefHSsdnXpqp7JyOseLGGI/pAk6EkQ5+
bij5QTb/y2xT80N/eDSJH4b94i/OWqBIYn0+Y+OTITMcoTX7eIxzDd4xadodEIBRyEvwkhiR92Ja
UAr8VnvlNJrA3yBZhzvHH/L0kHhaZdnM3cE5xLvS1t5IkMllxjCSREEZAqaw6VGRqXFvX2c/tpOf
43CtdOoKFRPRA1Iz703TLRw3DFQz0wVDqMZx5uKMUfJs/Yf7yhD9vUHk0Z7m8DM2vfaXFM4J7wTx
R7kP72E1dmrnfoDQBsVMthJOu4bEf4nxGwRwnPqgvjy+91QeHUMR3oj6b8Ek6MDOyIaSjd9Btvul
rZL8a9JHhzCpxSwpyTXTC+3kfEVpIBRuKC3ersX9KfGKRghHr/EKfXzGqWSpPryZTwkquQJmawDZ
phJrqKDgOVjBPciOBNwRy+XseEATiXWCFNUuzHF+DEPzCETfTE72vTbh7xjsIAysxCk8zBK51/Xa
I6LRDQMbP3B+DcCEWEQmoYyeVpu7MQrMLnsudOszT/UBKVY+0K4b0bAv73twjr5PstxE6Mp3RrzO
ArsTcrJiwg+OldTDWr1PIhcEJDiWWO2Jq2qm+JLgTYjj2YrFe6sZQzevAh9KejJfqnmm2dmUlX1F
Rd+vgsXvIvAdDPm2bLcuhHD4xYrOKb/GyDdx2BsdYd6Sp80OwFqz5Haz7IaIwnmHxmjSJc1TDs2y
dhHyXUMWBM3+HkUHL3wq3wpat5wdWYTESjhQQ+MsQzldVjroKs60WbRqFgXPy74bDWlqkIXmztS0
mPJ6cimqyxSu6J8UDbjLOlTE3tC7Eqxbfv3RzyDH3yT4Y1kWrbmdmcMk11psq3IogoSOZnupR+R6
S9WaQP3l63y+Vh0ttM64hvTKbKzzNggvKde/puD/w2V83WaMDdyP3XvJU5rmZ11OD9AJQVXq+2MK
Ie6Sr1pA/jmHqDUFWLvf0a25V2YjO+SJ9LFI51ltbRdxmPgNjTUWt/f3WMd/Shcy4w4MF9VnHgLs
nADSKef9EJgEsg6QmexnLco8e2BioLjEXJThVFTYehqcKAxLkiWmOiz1rI91Jc/I6OBF0kEZMc1a
TbzoWt7uqycT4X7jSWwXYsb3XaMSScH555p0ZFz7mgLHZX/61ZTDmc8g/NbN2t6Gf/pCZOxxyEjI
0vlqF0/lYZ0yWCraSjLbcgSR9jxaRTUTXLlyOVMFzFIrZb0E5k7YR7SkD7NSDbIHxJMkWWq9xOM2
oKwx4Qu1WpOVQYcIr8yTfLHyCuAuvbPjwnz6mXPUaXZDuny2WkzH4+N+w8aK3SJzICeKAjpPb3EJ
CDaF38/zs8MU1cZVnNWFk+WwwdPVBjo6Cb16VuEAdEOiW9IsgzixCCBi7F2BbUrNrydXflMPEIsi
xa6kK0CGCFow2qk1LfV5tTWbLhZiwjgEojePQUPMw/kd0/j0nNvXb76qY7f3ZheTtE+aVhEUpZN9
7OlZq9xHsgj53nzAKZMK1qdljP5udkMKnieedeE/Vkq6U/bdlfEXTxenofKe4Ea7BY9otsA1YzA2
NBvsOmvKuR6SKntSXoHVGbM3xd3bOELCkoE0VCQKxfqW30DfQvSE9830A28+4tFGxHwZsGbZskSg
KkVJR7NaaIW4Swl+ynYlpUMPD4F6Z/RyaDqpTP8i+rOmAP7i6n4ktb8f9yWzm4jmnxX5S2taY/Ws
OswHYILBtB6sdlCJC1Ng9/ggUXGevHbIXVKk+C4A2Nv70R9VvKQefHzTZwylw/FVIk/X8o4NtKvg
83RXjBLEK3+71r79rsQhGWOjXMa0I3F37umuQDMDEyvSEtK/yA8WmTXjvON4ZbtlpBJAKG28ylmN
RkPoMws9Do/T3JIp1fZOD5Cb8hUktlrc56skzSS0cckhwxJ8eQ0bNCoawc6szMb6j6sb+A14H7so
N0X2eRnPaG90vQ3IVO9vFexe9qMThSiRm1sluDzLEJJ/6WdjoQIBXvfEbhpX32ZzmNuE3ezamfuT
skdlW0aRTr+6W7EHEIY/rxtJeMW87UQtJzGtQ1jrpGoVkT2gPZKThJthqQ9RbtfOJB4aI9ueG3fS
2KMrjHrByKahJlfnuRutOobvBl0jTX7hcLe/IdTR+NptE78Y31/tT4f/OCI+74SeAp9ClAdEQtJN
fcVU6VdKKoobQifHRG+Kvu/vAt3HajjyCO7pdg2UYITiE2zPXeheS3GoKLbmdWiGVDxqsYxHK+jh
0h9O1ZexfxIxFizb2CiB7lydtmShKsSePkNme90DP94VrMB8j5BZlJZbcMb+MKpijcAvYQvnwOUT
Y+alvl5KR1PxwjPmgqqM1F2Zl9b6kMO1wscpazLWMSb07j3Z3GQyM+ZuyO9UHqlpeBVB9yASVzRd
GlMPL6zadHC1B3ROsZwcBuF1iFhP4PpKf7cqF8vMZXCBfmv0m9o8Ostj5alNA2XZ+LgtQEwOCp7Y
zPHMp2iXMBGIvqp5KANfjydFcDV/k16O3KvSGOMny3Sp4JschJS4F6YP6oX7f0byH35Prbm4LMFT
pfEP0jq270Vr44Z69/RHJaKm5H3M6NiWW00WniMnyAorth9e1X3qXiCScvS9GTSVtZU0X83sPYZP
dvMNRRIxYAocwNLJQq1A7QXytx6yutwHOjSy0EtMkBeqOvXEKpb87eLmeIPCHuVcNObsx9ubyh8u
M4pcfkIi3MOsVguHq+/D11eYWO9f5GJXUAsA/bZMgtErAPAhA6A0f7sQM7JHIYQNSwW86M482Ppk
82/xImR4QFrtQU0LEIcbi73EuuYagAeQhT0aslQF8SRjdC3+vPc58VSFMPYNUL8cxhKL6TJZiLYQ
j2qqWr5+Sq+oWMPZWbRIctBZURPVgjclHnOB2I6Oe1T5Ex31EQBG04MSSo6Amn/pDjYeN9npJeak
bYglPv7ux67vE2X0qkW35h9A4+O9nhpmvrU76MbXSlVeOEJCRfkLUB1sKpN5rQtxBTNnRxxWAOqC
kIPtE4TdPBooYh27Lqb4D7zHVP6/Aa54gcRFIYmAAifIlQsHG610AOFwNJR0ujylXJwQzukRxUO7
sm8wHBaQnoC+jbcuzQ8c1216uLbAsgYWEpMnIMyWRrstLMsm14b2lR/PZun6bmRh0xYKL/isCwGg
yMbJysbbTTg99y6m4LvvysMEltSMXeuO49XU2Q4h/fqcASL/DBk5gZ6IzFdtTa7zcUopA6uQuLpw
DefRFL3eD1xweoKw54naNfX+90Y62zvMDHvETlnu+j8ncKcjPY0GDCMKLRVFk7qqfAepU/mj4CqH
jd1zN3k1MjeA5EP5SK5xK8MFQCfTrU6i5XrKj4ZrqSnSp7nIAHujoSA9dD+ZpmO1tLUy70Van3s6
yeBBzLndbRAq5x63qJ8I19e0WCucK15Ryp15FchajowBitaAaPJvtALcR/+1KmTGmoiZM3oxRite
rttfzB7Lvzt/EV/M4tZw5Rx+4fFaY1XYznjGldvLjU6N1oSiFzWOgesDv8TqCqxX3DjUKn9eyFe6
L2Ds3YYV2of3eOwytsd/5tvNxKf3xeP3W0naAFqEg5xY2f/6/E4S6Kv7Uf8Wu4N05OfD1L9dUQjv
UDoJvf8aZ4KyAwuEihept+HbdZGrcbTBU2vnEul+o7dcFeZ4v8FSEKhWO/1Yil/zSh5ElNn+Cxc2
h/IBcpd3V9s79+oVgyefeXtDMSLFnSJDxQZG1IX0TP4X0BAF6x11Y1nClVkLD1UOIKraosSZiyJk
hzlSCnEhQE/P6eV/IjJjacoLTmZH5tq/sacWmhakxXWof3Ggw28jUTXXVJXQjB8V0+Q7Hd3bwIXI
ohnj3Ole6VoJ5MRDr/00XmU6fdsbGpOKqZdTk/c9oaSqTfWSP4Rr6B7XkKZDwsH7nhAhScP9L35n
5JDvD5WwcveQG8Rz46Bram7W1LjlDO6HubvurtUlabhzDzCHPmEGfAt9kXkwWh93zn7MtgFMo7KN
P4EjNEOLktuWw444xDuwXj9xj5/Z4OX7METRcmkKZIHeuSnl3OHQWhrfiZ7D+EC9gSLQA2IuXOS+
LMmLLqRovJVDl8m4qzsRRtnvCUckhO1ZT0rTtba3bvm/ItBppp+QBL9KG/UM1aAbTW+l4yVhJYgM
cLmq47KKAQiRMDniMvijECEnKZFZOzd+jPnuQiGw6IzF/LP8MAWHVCv40rNZ4eoTft+NGAYZJ745
a3Gt20NgwAA7DFTq0CNYP9JMlkYlGO+em4pMUhNyJCSnR4IcghurL6FNTNFwh2ErxITUZbJGZxyf
pAabFRxQTWb02hgx94bfppQGHEz6rgQ7mFlQldS77Mj3Cq4eVhr6r++hMfMsSmz+DLM8NRd5RZHv
soiqm7yCs/Xh1X2PdphrnO/JPVVO1UqNbk/Yw7JIfg+Dv0NLy6mpjIDfGp4xDRvpidSdA34N3RQP
xvIjGmW35O1vIoMKo0O5BuUo9At+542oxsCP60+nCy4lcjfBxTSHpK93wKFqRqiJ7xsZjE21fjRf
AA1ZLYpusWfpU82gUSK2b0BAYZyNPS4uxNVPsV2h6bn2snGHz0A0ThjGjVAXn3Z2TVqzNcGjjWXB
k4PqMsX2LAxM6CR1tenwtT/4wk9aYzoz0glK50XkZF0EKe11UI9d+3yB8kkwd8jPgEiqLCx3koIF
xOcmithPA4DgLCcqrI7z3uEEANyvJZTRrcs5un6lYNan+ARZsH4hRP24JbuCrzblCq4B0/W/zSzz
/A/uDcDX7FtIOO+aNMU1suBqmQtMAtthxyk6jePndQOtQ9pumbh+jn9f+6MhvCXchCouJ5tBBSFw
zsL02Wgnaq3T1/DzyEDbqkr/+ttjfKxQgpbj4eZAEdy3zEWc76zycFIEz2DWIGW1OnTVETWX+2EL
CwrE9DbYrB/h383T0PX7xnzsm2i8c/hU0jAj4GSyWRvbFT3MizKzDhzxgw3Lt4eBiu2hldEuYSw6
IRxX01992enlCjCVmfUHotL55l6J9T5+bn42/aOdwWs33ucUpAKvwUkIaHHQMVxuNL80+jf/A0Lw
iyXPGJk0P/tQrW6jBb2sPBT6dw1CP93pRXQPgEXNGkXnvBfp0THXBUoctrqCHaUlKOQAWdgM+yxK
xDoPOtHBWjfdxkJksor4MUjnbTUezkps0EWWMYypj0+RuT9foPrNxvaqQMRlfCEHjJ1NNOG2Uvui
6QvZUWt2laSxXxRRDtrKcuZ/79ms5t9dlsCCzUlkwiQGaLxQvjXFGF/7kxQMB/s7cDcdJ6GyscDP
oT2lfjn+7suVrE/hWoYNpT/fqDiCCq+0h1bYNhJuQJQj7647WTS7OzGqaIfplmiETQNQHT8aEn0B
pd71knsiZjt2yYYV/PHjsWeGdEo/0ARtP3tdyMYcLbVtnlZGAeJaC/2yPFiAQ0fqo2bD/ZlTWbUI
80OTdodFTPIOrvAUUukCjuD7NycsWg0KsbgQ/iLwlMFbTOry9Sbdo62QnOSOoWwOM60Zl0KmgrTc
VGKBk1WRv1fJV/MSBOOA6tdtv7/KTOyp11lrZRs0arfygRiWrjUgYvBBI7lvHLONdHKrVrSmnw3R
e6seDdhVDWOL0iBOdUCGcpwLKNluGzoiu76xiXt0KtrPFnh9l7WMHxDuQ82KBZd4lS5eeowk7y4O
ce0RjvqNFI6u0bql4TZD2auTViBK+QmQBqgDLGWoONG8a0IHrz/SZud4Dgfj1x5sQHrfaxgMWEdE
OTRWFGLW4Tc2VAP+4kxIqxV1QRxZuJJ+IKLbOGiDK4DJT9t+kJ7l7bhkS8vUcJ/lq5gpoas+hp2R
rwdW7FEgBg+pmLXBMo/tjt9fvyyyEgwpEY4VeRLgOEOs6UmtC+fnu9oYTaeXSw/HRc1V9+Jxxk15
HlD4FY3Oz7yB28z4tuvfjjLWJcHuzABoNAVezRD6LNwNc3ri0gELzPFYYVFnJFuzK46J3mE4Dcbz
niNZdI7RS1GOZBEz8+5dzYZUm6Ok+RI6IE3DmQ0NZ78bYRbKkvJztPFqLJxtWmk3O1EU5F0D1Dzr
NJXG6wN9Cks4qJIKJnibg+I5xHEaTfJSLyc+XNnwfhmoUhByaZJ9lgdwE61MivHLSbDBdCvmd3nS
inWpFCG6e9Sf0dVplgvpACk+GtAjLtSARptbl+h4hMTnHrC8C/mGWz3LHF6OroGHozVovIC4i7ku
20wrg686rBLotGu6Bv/vw65zqfGXYW0bMau/3TwxeLXFwut8VkCkJNqH+65s0o0fi7CK2DOxyC0/
ki+qTMjorfMcs97mUNuOeSpGyL+qIZh9dcGOgMpeBaQVK0a17PkSi9ZlKtOTq5FwS/T8zmGWiDIN
f8SPTFoDAscauVkgDvQjgbYxap6ftN/S9+i40MYk6A1//5cbNcB3t781W5/DVhpONaZrpLjJZqti
4dlVZlQr/24stml5Rmsi2e4QTDGleImIIIhNs6T6SUBZEkQyErM9S+sMjagbEm7hI/Xt3FkoZkD1
DBmAJJ1ylzCamEq8t67dQU5yBjBWvqbDECnjEZHXEWRR2c8FkY77GPW9Tg4XhpYMka9Ha3Y8QoMS
YVP+hZOEUmOtaKZB0/bvTmG//PtdhIAc4p1VTMT+AynApVIsAURG97WaOIwmw3JsPBU/vsQTltwR
6WsZ1R8PRg7lYeUozIjxy1OrQ40zYdz7CH83+B0z9/aQIEEzsig0JIz6/xUvQWJUN0peVnXIrRYo
cbJj+n0L0ODKRxLOlPu51Am/xccKH2FJFG9At9mvGaEHziduTCNx2JrKMpAz5rm1xQ7EmKFFrOmC
WJ2nEPtjdFoACwl6H1MFHUMTkzQ8Y4Bt3tYbJ1QLfXIlBi8QulzJAyFxMh1QQZWTIOGDc9xwvM+v
PkJMa05fs8vMoKxVDKnncj6iDDOV4oZs5z53/pdyvaJxg00gwFfuYa2W9tIW8jIO27wV6tYmn8vW
969sp+tNQeFgrGG+Y+Lk0pBplefgdd+ZRjT087ttAOdTgqJIhsN0rW+OhudZv13lEv71RsYGrf4P
8aFTksjTFT4BzPMSzcj8kmGhLa/P71Bs/5O3AQj6otOgmei1oJH6GdwqRn3MQ1UkFYznyMswQhmm
oM0qXK/lTLQzOi4vS8NXKqa55kGjnFrNyZc9AQTrUjD9t8qIZkVEV8/IbJs/M1K0Q/J1yxewrggn
L2UG62YpXXHmN4ZU9s6UqX5NX4EofK53mkLESRFq5qUD6Fq5VjMxaFOb+W0wWvpRXzOp5p3zjcxi
Vz2nr95PjKLuZceQpi/FbSaPy5fFAxL+lzanh8Cgy9f1A0PYcUA+yFZVmxiEPbTYIwRvVrUDSS+A
OKjnd3jVxTwdpjWNwkwj8k6bSQZ2j1qqtBlDyhbarH2F45tbo167HWOYM39kNE+rtzEbGluqTllY
BuVeJq+VKKHkOr+XM+AuQIqIDgIECRU65VDyK8FEr9QfZiHkiHVMBKUVtN75PptZOieCM7OUFpYr
TlW2F1enQMdPTqagnhfUxq3W41Qqxb+vROL+B7d6kaP48pMq00tF9UdeuXWiXPfqT04m6t7KNQrP
tehHwWbR6FjCjyNQ/8hFF0sB+cgKx9X0QSv+iVqa2f3zUcdnHW1yu/K1MA0GNeCC2JMV+xyHiOOF
yX2btZ+vcpk9Us/CmVX/Dubsv04Nh+LtvgqJ7wvJ1IpVYT+H47shu9s/ARQpyfiXQglTycGA5Uia
A7LxaEzAapT2llXJXVL52NSgHYI5lBjASTx5smX+I/+qLZjQoq4L4C0yOnDX/2qTxGnIEFfcNd+9
VQcry9MJlIJRXiW53M2lXxRZhn1p+cpjFDqcYIXzOdgtllFBqaDzo3N8LnMjIz5AhC+0/NIU0XeK
q2bzwOdCv7o9COUT+84MekQjG6Gc/fPOUrooT/GBPJjARNDzId03XAatN5RSDeAWT3r7n9tesjra
nUQHRqvMlaMU0skdFTcoVretWhTrz1WG9Ypus/rRGgCXPd6867V3pxhXh37n71IL/NSm+ktKT0GH
FD9NL6wG7jCB5HXzSVccJtGvoNmnrBJgO4UWPpEb4iyaqceTp1lgbH9IHQlOrlzJue4cYioZYb7M
UrIt1gBHgoelXoZ6H0OaZ5dpqAIlF52e6DlteS74vqOmgIehvnT0GSuvG4ce8C3nr1Am9nb4z4Yo
DvFRiw/ge+Eo4YA9/0megDlz+eP1Ru5dnYsthCpYHOkqQgotneP0jGoTsCpLF5DHeKUZ5U3bZ+P7
biYyP0vX1tyMtFZCM+p+rLrv+J1ccpDPdcgKbcXidcRDCJ8AmyDG0rUCeQa9Qt0qGo+p3oqSMB8r
KA+zoY8W1yaedPjNP6lqbY+VuKHn/AeRH6EBj0t7T2HrtyaMIQP9f9uRWXCZsCIJdYMbNyIelhCW
4/Zy4aLc2+FoBYTv9WdDo/UTNxfS5ZARNxW+QuPd6nYx1rfeswr1in9tAcIoJsZzOu0Js1E6C5UK
NDCewQSQChVNtk2TnGCaetNITxPDTldQ/dVcUApgSk1gT+KSYE4p5l8/LbNCtN6D3exuUUWHVGPl
6vBUZVGs8ECrWdiFD6Zw8r61akipJJ6YMeOTRPMIKPMPNKVJ7XX08wa8rAD2Eo9d+QPWmXtDkI1x
7jl4aFGTj0QpZlmJss0fAgIaXMU4uLnqgRAstsJn3HbSGl6/Q/WU69hd/gLTKsqlMZQ5JJTyeXxP
dfE8bQWQSg3x/KNaeeEj08rnx7Kcub1DJpRvSl23sCsQiazqwyw90eNxghYgP+zuFhFvFREAk6uS
M2BE10E0AX89vKH7L5pk+6SVZJXeqlV/mL5L4ZXmHx3TRfBbxN/AJ6FejSIekriTG1muPlqi1Acg
VSGIAfjfOr2g29j0YlBKM+6i8kQlXIDWHLOkkQdF0vtUcYdepqq5KR0b1c2+PG/1Rpu8eBRxjno1
CS15oUyYX5gDUBZFS5hmK1N3FOlMZ0RgEHyvKzkKd9hPCgtUEB1fYYOOMrk90Bwqb1gEPbgVSajv
x/rvU8cmm+r5SP01MIU5a6wZqCUfLti777xBxhRVY8W5ZqFDusvikckWmkidwQf+AzVzdNYTBIO6
gc0KzNtXotjC3JiwJgXOqgp7AdkiTA9ax81QJWKGiC0xn8iIBV7I4vL7cOkGh39RRWw0VDKDp5V1
IqCOpHP0ULwOS+Wxw8fq4vISHnSJAyLkiy3KWLgv4m47WuE4K/nr5/8b79WmcV/1R9xHy1c7n8zE
0IEDi2T6sZclScad3OogVsyVUYxv28jYFP8kKfai69YLXtlKuJdlkd3Z+b5wbKzxuX460XkT+fgB
pLmj/XfO4xWUMtPEmnvAEBMOGtTwLFy2x66mMD7fVNsh5rvXgjq9NYGxCZxa+Nc/VEZnFOLHav56
xXrInHHbGvXRc23l1saQWlAM1Jb50D3f1/LJ5Q0G/l+VVZ8C6HyPKV2B1WZnkMdd/hxZy50oEcXC
LSEmn8TO2NHazSUyFecBMG5JrGrJYJLxZ9qe6GRz4/W3zc2FwUkmvaiXD5OQIzLt4MSvpIdCdG7f
h+yzxzujEYw5vsSVPwDt2X5OXCh8iueCHUbYNk83p9Pww64euOcFIooxUztqUI/HL7ttLs0qGW3z
QSnya7Juenj22EZP+zcw9AlalCKGVutnhk5fhA7kF6cbdXy9bpCb0xQQFjXDpC+EIVZoiioxW2Pd
0DPxL31GOmmHPFg4Rq3ajmgql7GkDaW72UHvbNEzmVpoAfysilP2Rh+B5DlbP1E3DQL5M2+blu3Q
JhRtIhpSX6UNVBOgAfhG5GZQeq5/9zAz/tbC8QScAnzzn1YV5/5mLs1/l6n/zsRVxrwfb5krXl6/
AAjGuxKybOM1mEj6wHoFP5Z82JttP/zwMIQ30GkP14CjpdDxK2WdtUDVvjIeRGyAN3/LC5xOYD2c
P6g1Hi+JALHYCKGqK0g2pmFUjDNJmrZds5vezIdCOWGGXygJoGDeI3zwlR7js76qr5JIDnPTntIl
gNtw8/r2lpyUKYyJ8SJGMWst+yP3O5iahzRt72H97h7aLkIiRUWx+++MZa9iapozFadx5iyq4A9I
8zABLwBDbuKo5aALfpeV+xU2pwRX4PWiOJdKH0Ac8WNW6t21AC2leF5Jg13JZrpi9aYkW1JdJ/Ws
G0gFPTUMHkCOKR29rDIwCsr32pqpNcq0TgcTe1/3OhWJnFvFwjwhTpMuIGPjafGayu3seSJEr+GT
QlUvYTXc6dxmhu9ZNVsJibfgLxG1yJua3BdmTUoCqxyMv2E3/qErb8xEgEokJ0M4znL+QO9fMxm3
9OKIVWn1njw8ANIAU3W644TblJgsSAmx9iHuz//29gWgfMwjk0ftnZBMguLbZLld2mDqlX5gNSZt
4I71KWvTVfh/f0tSn0FB3hG+GjXTAYJr0ws/8xdeN7Jy+TbjKgGykPeoAPPL52cEurXdcJYJyN7s
5a8+OCP5tshAX0weIachqqvkasOIXHrsQVv7sv42IeMbRS1zAk14Rc8maBXwz87+1w7GWH3BGwrq
Efm/C+HqSDIfHuMFiEQRIChUEpfovWPyd76ORjpTmht+2ERw7CPPQ9fHMaHIgziXuBYYv0Wgk6p+
bPfSUNjtL3YEpS+qZeDhFlIdbDKeT9IwzHOvduU514Es4v9y3PnsjIBPyg4fRhDsnMJn20mTBkfR
7ls3f4j6QYfIX+LDAglRpfn0Bg2PTsbgnGzouQLO4Mm1DP3hs6EX54oKuctgZX6evEOvbfKYwltd
WKXbcLYxSdHFmouE7pZ9Aale+0egb8AvqW+3x2kfkYJioBn+OtVkP0mSTPJZ+Y1PH9Uc/5PLea1z
9wpguNb0385WRXqvy70o/gD04brZ4hECaQ4OrkRME8idRdqxhTV3pBgAzwQAo1eNjUHZiJ+auB1E
YQqF1FURjb6rIGKEwvnESy5d6vjxtt6Oncd9W4mLlt1NxoV/wjoEFdG5Kdn2hY8CTiOGAz8n4VFA
saj3RPx8qFlbMx7S5eG5snT0qyn7DRXS86f04d951yIHAdTxN6XDrfjseg9nUe1ydZSDT3Qo975F
cig6ahjhhqi01+TW7FQ6qpGSm58iqNrCzUvZEBkIi0r2cdWZlHKIZpmq1uxO4URhaNwrtgI+1I5R
pVNsb9bV14nRD8k0qXKUpr79cLZE98fs/H5bTUjv7bAywoaec2JL1j+CezNZUe0wbyg2NQc+wr/b
wa+1zDzbljbyA2U5BcXaSP37fozbNJNRgitNIHNbJPppEaaWI54HZUi2cWNCBIEC5EvvPquaCOl0
lDzfRxsXiixVJp+z4r9BoKrWZ8klpvdnT7cuio7iFkKOgh6g2R/uxDSOMq+s/T2aQOynTZFdDa4y
8/8aR8HRWPqzD5Ms//UskU7SJBizJYsautBphKz874dSeb5ZBKardvGhLarGQmuLmC2az8+tW/nJ
7nwN/AIgmjldLWNJwcAjAhL7UniKf32khjMXGd0QDbvfJhcdoG2XEHmhqQPDhhn18Zv+VFRIKGnX
0h/xyJb0tIvUVLQoO1cBSyfsoVryHoInf6ElAdpceLROeV3kQjN0lh1G2sShs8GJ614nBwEDs2R8
dYYKZ18nLsNYIxA9iW5+sWH1jgWnI50lrd96SAp/lLkcA9gXc1t4GL0YGnuDSBrZPg+AFVCxfIjk
5tbDfi5uwzfBheqe/aBNBqd2biy8HznL0VRzVmJnIJ9xKDlRM0PPSg4cxwOgXZ6d7BGPeQkbIkFQ
MkDeFhoiy+bzACVgIjoxPv9uUJiVxwFCgtIc8tXBl7bbpotncGDQkIK22tUSacSyhHGA5iMbJoXk
2mz9gRDOI5zGmX5cP/02St0OQ3tsBLI5LtYt6fuAzc0eXjKAQlkfnsKlHSCEp5Mc6EMJkgaFIF5Z
0X9T1avR/z56HsgpUszCiuT6oCrJSLvoVgJGEAlEOCq+yJP7cr2z+gaCfCjhBrY73gysFS5DOPUG
VFjof4Q9wNLHD4VrC9bo6hr+lDA4cvuoIMjUQH4JAkyQbaLbKVAnZmHBGAoI72H23r3v4i3RXl5z
A0K2PJva2r0sglTRz18V/xc5dLV20atjEsL8Ur0o2d4XD6r2ox6pJIvRC/XHkq0SPyTcLLKs/tsX
+3mQkoaviMSAC+jkdSwxLzr+nz9Oo2z0fTkY3he4hEfEQWizn8SbXQJ5X8z+//f+u+9w0oOzgE94
wxJT1KoaT5yoAku1RYVbTp3s9dAQOshXSIAWBI6JUzfr9FKtEiwetgksAQqcSX09Mg3CmxOAjdHc
X1YYU3ypxCoM3YNmWxqzQ5O6UIimb0h/qgZ5jBWzEtfcLRrWeXdvRr+Q1DkPDJyrL+bwmtphrw+j
fxSHvvHIX7bDxcDr/46Mr0VgQSMOpxYWCi1cNsyMXD6CBDLnvaqPmIGzZuhbo5abkqglnBHsF7jf
FIJ9JhP5f29N5ZMjyaR5vGd36pC9qAw3b6p67b9GmSvIaSljwBg3l9g2tbgea1GGMTJgQE+hWuL6
xy2KzGp47ZGJ3RC8l+6GZ2F8iLvW6FjvPT9Qp3NTCqelqNUsckrjwjqAY0dtybOIRJNI7DXo+rRW
BQLqkSY7TQPT8903MR2WI9bSsqk8SZF/Yz0tG29FsDJ2Sl6XKmCD1q+uRaPU8jnuW+JKG6O36QTS
5GaCO1o5MPz2yqFYNyLrieUyV2alU2s0V7O1cf+s4YzEYdrsjMsnYpm5rtdFnCEHapcCxgzTe8QT
oc+n8Hw2T3/HudRkC/sgHECz3gjVq8md3MEzcZ1fFRcMLSsdowAd//Co3pQC5Bf9i1+eyAF7WSEa
6Wps+vEhVDIvf/npcxtv4USV+/f5LxsgkAg25j/gfve9y9tP7WB4HS4cJ9dFWHPt+Eu5YcD2V7N4
WzQkSyEsKLGrYBzME4iPF4HCtHOCUCnXFwMPenBGGZCYRo9febSeYfmdBcyJoxMckQinPfg+ikWg
uwDaBnDUJ7wXvJ7Bj0Aw4G3J84WXO5uIC6DwSwN2NngNMFLKECxPrc3Q2spPgKA0RUMVN0qX2epN
mj/iWyaxPC42bdXJxum4JAyBqHitcOzLJm2QX+tEBlCis8KBHmKOGxvIhO4sFnebgQ1dApPBEdS0
xhVZu4+nMlfEeAdVYB7oTfpR4STagzri9l/gxev+/L4s5SwiW2AQLHTXqqXWOOOFuS9dfsOLhTg4
4SnzTW8MLCnPaSovtq7EgLai+27MF2ma9joI2jtPK1vq2+Zgd1PtNSpMT7R37nDR4qe/9B+AWWeI
2fhzFDX4TNFsLc898K0dLpREGuYhI8g8xRYiXQOKgqYVWC3/8dZpVgZu4GetF9+Qf2bDqsijU7lL
huBgxeo23KZmutpiq+baJmWi4ZX24SVVJq/cfSU9xs7t4RYC7b4ZkJffgTAwLQqUp+dcf5uLkp5x
U1oi3/E34fXkmbvYL12f13ilBuqStlbu/dKpGYLqM3YzItYE0zmx0w4GOiXh3KYFKNb0GgQT2NuL
0vNfAgIY2MtxZdfAKVCMT7YYPctjsEXdIR+4Ll6mRvL7YoJBxCXjsFEL07F0GrP3MImI2gd5b0IJ
1ZQOWvy5jr9FDWY6ghMwbm+XZ7p0U5ebNTBcCA/V1o4YLLgFQsUY7alJOd1ZbfrgyQPv/jptlNur
t2sKB0Po+kWe6BMvkJTK6gmNEMcnEvM7wOPeyCoTQLdTuUsH8ZDgNueXVFSp00oR/uwjowo3/YmF
zTNOhI3CW7R6bSffxbsbyKo3KeIicHk3EuQCyVGpZNK3WAIHR7bRNLkQpWSVvS//lAX812jSw7/Q
+56IRO/llwyDLrE5pdiSSaHi4+YGQH4JB0ybVPtgKA2cBFutTdeWVmiEg2rx1pEJaVwI/3UJE8Oe
I4dvJ6PIF/75a2AC5PxMI9d+yu8yCPzSyzNjgd5pKJgKYs+YvAAHp8miNtxy8W+ewq2rql0A87VK
VQ1q2htxtcPLdN6jiZecae5o03ARH7PJeSdNk8zUeRoTBOhM9omEe3aGW7haEkhaEKaAeT86gvNo
THOgRyggFpxxIqr7w2AF/PuCmeYF7etLdKavP1Dxt9h04f+7HUyaJs64XGPy37V0rJDzJy6woAt7
ONrNJUAVwLF9P87uKVHr2kcBmdWN8swl0qU/mxVGuZX1cW9x2yZ32gxouQ2IKN+YGjsG5dwJxJyp
O/0iTx8aEyFut2/GU0w+v+DwjyWUm0tVFF1i3nl/zsCr2DERKSjqyl3bhBTxECCAt6QVie4ZQZWe
BF/ptJnFIJXmghQqLCb71Jd3+VEYLOV619pMuEPLkEL2s/LgEZ/QrX2h1J3tdCS+En51F8yZBymq
PCJL5neBswyPjktejUvssBVbr7+GdGGShahUkuvMt3CO1yVN1fqFDK15BIwPSztf5nlSd+/2oufI
LaxzwuDW79C/9oI1BIz4yaSbuFyaZJ5I/sU4l4WaSfuihMs5EwCuc/uJ1QXJFVK+EvMbdFKrY1tH
UQzLgn4YqeHoIlqDR5tQU3cgvZocrpMRPkoz1WG29yy8+KkXIDtPmc0+9tb4A+6iThv0eqrk5Qxt
Vt9demgp+k83zhyh3sUPGu38ZjiIraJETCfB7V1+gFokkbYdsDN3T2p5DTe1Y/7iGQVKm+fl7Nj+
rhPDwQOw66L5VtXBUCcAtV720H8Co6U6FvOW4yCbGbYvysvUE2/MX96li0a6MnhPesR2vxr3qNSO
Smct0CiOuZXAvj40Wtom0TxDJL0ib9/lre2uzYKBUOfZbOsWcdJKDtfncNLs02Ed5QoDDGCZ9acc
gmVqPf9INOTfu6amRuKB2xLjVzhHhfyWJa0iJkZ7D2fwVXxqcmKpT+XX04f4qyOPHUM6jwuVKFyV
qjHm5M/p1SINE928x4Kslvcaom8/oRKuLV5Flr9iz8ufWQN6ddnR11St4emsRNJk0Ia1I/uxSTCw
HWqYiOATsKP7QnkYDyO5EvTmkSkRcQoDwG6DsYIa6z0fFitQaQDqBf/7Kvvz6xOjUryE3lgO0bTi
f3FnJvB5jXUN5SfJxXhGcfx/pj/TN7UJqPBmXSvmVrU5Y5WJ+oy9C1oFTlObJoCaqNQk5SZvj9ep
/DjMZZOJeEhUoecUVVHfpojggra09+SSzTSnjbSZ4b/hMCgPdSJJ4pncmEznt/SjWFncNTlEoJFQ
J7sXgWzPIWm2wNVNFNd6vui3TrkcSoAnGS3s/L3V7Xf8fSG6GjWIhnJDRd4l1Ur57uOlvYdwBpIE
2Fwnz2qPmVwQneVnHRY05ZFdyhjEYWiWBu+HEVaCJSzkuiMlWU01OVmLveIH5JFfLMOTtoKQLGT8
u5ZNMOvyh+xB8XxLStZEkzZ3nKIM17+fSJMIduWoLbZcCw8wjrUwVKD2JRICuHKBZNrBtR938s7T
QQ3ZcGftWPkAoBrxoFlyzHO7htKTHamvzGW9YaNSmTq2OVsARxyQ3xIjh5Zi3vLR7rw4moJx4aO2
px1YJRenwcJVQIeipc4DvvDaGbf9N2+dY1f4zepOTvhIsXtPZToQpqbxJCQMR/7sbzFFbw71sQIn
P1sZyw9ngHBSrRRWf4YmMi79tkjlvdnEdOMAlqXGcNmXTlgHUCLpUKi9qotyLMssHYMkb91V3RBo
pFWK2ARaDnJWs909OL6E+uXkKxxMYSZgfBRykE2pxjRfx29jWDzI1ZFy4p9lX2NB2kA5OcyIkyJW
AMD2vaaclo26/eW9/xi/ZQlDpeDuEBu+98PFxxPWqa450gTJIiHjxbCYzbLeHcAslYfMhUtrIJRN
tT2w/QVDhVK+M2ZapKV0u8XSoEUUBAbzkjBx4h5Yf934IsIwj+kz/BuNAGVr60sa7yGDJ8Bzy26X
PasNGjI1/gt3YH/6BhdJ5HBOy0THQud9O74ZZGaG1qAc+wK+ONnj2H3ugjGIy7FcoS4d5ebp+vgr
VQjIoZUNaolapYkr2L61+ezit+pbdOaHIg0VIz90KhtpdCSqyigxFNS6BxghSQe84mGSvKO2J1H7
OxtDbWDV0+BNH+39sJ+1MICm865bTUVMDgFsN5gQaLYdPxeW5Noosof6V92kUHhhZidGZmYnEYWB
9E5xd+owWApThPJo4nswqUz35Aeh9LlHKT3mE6pwyyjdE7jOlHc1Ug3Nn5bbHnTcvEtL6Pxbg8eR
TyrdEZN0cKdWUwFjorRKbxHXZFlFns/Ytzxm8vLWF7o59IVJg19HQG/50tRuHEbCa/pgl8BRhloM
cmrWoGvkgr2ttbodl6eg7X0RL1xl/8+rGFj3xNIdCz/l5fV8iszAp6CudMfnnc9wxWKdxFG5WXDb
Nkn5zWBHAq0MO972j0SWYA9qjxV4x0JVnA81iNosqj4cURd+s4ffG191wo61mE3KERtIP+rCz1VU
Z6T+nucDMr0HtN2dla5165FKg6lLTmb41JhqbcF/V7QKs+ysV6fDNEcK6utWME8ES74WOBXb4yhE
Cpyj8/VV49guVaO2y2QanUNYjoSB/gwN4va5EVR+A+NhyAg2FBc4fCeXQ6MluObO3Pznl41YRRe3
dmc2PygjST6s9KLTlbwEQRNcGqKOv/IZtEpLWDItGnaph/UILj0g+86nA5BAxJffFBr7dlW1itXe
tiu+pyCjtvXoH8hO+mbkOdbF8ABPoiKQNm48UdIOyseleMGjY2X4FllQE764DAT8g0cCbZEUg1x1
o45idogyQ3Bo0MiQvUps4aVn3uWHfsxk8lXsgfs813LbvQleYga/Es2oUBXb79ap+5gCD9aV1mRr
5xA04yPDjfh2InMH7PktFgtAsEb+D3Kx5V4O/fOaw2bnnjHbpWtzO3lMB7M6nJ2Zx8LfWsYTuDz4
PlQ+93UEO0IZxIxqsVrBxpmLm6RNQL8I0bxgP3A/PAfkBC5ZtvfROfrBJWfcWcynHM4/3aSSJFgD
ssr8lkZ85VZFaLnQietlei4ixHsqpJxmFM/NmSlmSX53dkjqe5f3VPEBCziLmX3hP1GVr2HpcPsN
l/QNQN5+JnrecZl7DTuu7jIT0ar62iqA6GDmHgFM2YhFd18SEHHEvTVmOuHOHGBrpEYZcudi7S6T
cKJcjogpq3ebr+coOYGC7B/nnKFVxqfFm0mVbSETnk5B53QzuDllf4yAQnoHBfptgF1Xa58mupdJ
2lzBqnSoRgJMQmt7Jrv+U1y3zFmbAuPyU27tW62TF6u5bKvOaCjrQ2kYN0LcKIfSehebAZIdBgwx
CASOTrVdL2+/oU33ArWYMXWyG/LjfOaFRj0WzhNHudQLQsWEfQOpbyYweKh5TzhUDZjxddg8y1Np
YPtf/c/89R27eMoeARgxdzBBUi5+qCY/nXb+oXY22xk7fDNTKU8ALw9a3mFkxQDwT668pVdClmZQ
QHFG1OUMSdxpjReR2U4TRXLr7lwu+j3R+g0XIWavF3ZvFVhXqO6hJIda0CoOW1XxT3CbJe8relUL
cBR+TqOuTmpGXxY4xA8S1sQYAXHsu0nBYq0PpLiQVJGdZIxJVxThyP/EfXMP0+iYqCIIuoJ4mNJS
hn14fUqsb6Hv2v36TCB+VwUVmbaAk1WIeZ6huUc69f56E7OMo6/OReWGEDZ0TUo5l8MHju/FGQ3W
XrNfpLDf3Kwm60AD6ZHxwzNsQqijHhtnoA7AS66BwrLNqivZQAUhnVMOIFTd9rXQ1HbwQJcr/jt+
hyJTnwvvsztMy/dxgYl27Nits7Uqi0x2BQ2G3uOo+AXQ0EG97EeLJasXal7q0FtdsypOHFGYZPNG
PXklb0da3Z21rDIZ44ysqDOYKo6e3FgpTXDBFrGoHyBNDhtcOatVKfjKSAYQA17CPSF6W3V2XneJ
u+fwsGhjzYr6QVf1CsKA/2oxppzrVc4l5uAJArwLYYltNDTAf+ArgJiNw2vA4w32kKGzm3GVF3Ga
jMseqemXvr9ul7aMKL14JEXn/4erTYjNAPUpjQq3DuoY8liPp0B8Vcs+9fkR4wbwkPH6LHupQNoi
8B91ofobLMnZUHysJSQoVIFV0LtP4oO81p9W4XvecXB507h5MTLlMMGpC8q2HpPAFyoElOqYCO7j
432d/kPoFc6CalsLdT5ZYszHGZmlXY96GsrMvD211acI3noVZ//JUj1CzmjVFbwxJSNmvSlemtyr
ZqA7du29uUGyosfA5PaGFyijMXDxHpFisU0qXPnJ/Ju6dRHJhbwgPRkIgwtsQIUo4BKXChMx0J9V
yWTsL3ckJreDWamsG1fvzhmNpLqCJugsF3EA3VtA5oi7SxRpCkndY8bINCufAT+2ek5/JvoWA2n1
4aUgV57lBcHBO+ljF0jjnq7Auy+pyYS4FLTAyifRyBdHjdoqTz7REkKwB3JHoxZVvcVNPMeCUBIa
Ahyc3C67d1FoP0BCPQs6DU4ZTiSV/9t4CIm6mr03tCrUXSgoNRCKFzFgOLQ1abNCNZydUTS9heDH
U+8NDjiJoD8sZB8yAxdNMuQDOJePr2YTklWsrGp5Wsvv4XPU0ixjgx0zjAPXtUOQ9Xux/P5EM4cr
tWIroJlCtCBcJQJkcXegfYVCmcAushv0Nm5wiKGHN5/1tBCfJRpASJ4Df//OCDirQnOaGuyf585F
1JZTlXjd9FdLf1h3eCLsnqzS17nNnb2M1lp9f29Hx4kajIErHeZPA3t99x+mx8pBNup+R/DGtzqv
KVcfq6dmpQ+TsSwNzUs591geRQxzXTtAB6G7NknuH7S402d2Zz1Hh/J9fhpAgG29W16BMIF1NhVe
JD2Z3oHBefn0KlqgfDP0INw9yM6B+YSt+KkXZILeZXmWHBL6+rIjgkrpA1To/x13Ia9joRKil1PY
TTTN0UoJQdD1znjXYnZDowVhq2+q8oTHlsL8ZWwM2gBI0S7f2VbGwAkMDC+XXDlA1yrxlNcmAb5C
UMF2gPX1NneSvZX37lcpUJqtXQJDzr5w3NJqjN4TM/J4cQoiEJ8tgPVE+Uis1MNyLbefZIcge0/z
02Yqj+BZj2cA3bvWrVkiNHUw+Z8tChmL31xc7pwOhuZbzAOTEcBfZBaeDxCQaIH483c8CAQPwrf4
W6Hp3oTa/YDcDHONFTqkOPWCgxmtNuaVGy7h4y72cpkNkJzbnlfX5QQpgEEpTXGj7dlwNrrTz1et
uhhhPQJ4FtLEvjdeVpPwBgL8ZgsFhhhHthdtHth68mPuBGPBqrWnDHpNLw8zyxLiLoqD8QaZMKfz
S71StX8yADEdgVSkrmkSHR+IknxnL7w5sdRnBCUQ/zupPtl6CEJn9LdOYwUuSJdnJJcY6EZU8Q7D
mUyyjcBqX810Z+64/14GfAAVQyunZSwJR0x5HjkAfUfu7sHkEj0S7mE4vJTrkH/jSBf7b6qyAvIm
r8y6us1Klnkbv93Dn58zXyCIWqEypoVb0+KTVsBRQKrUsnXn/ybUB5INRMADQ4tYXoz6Q26q3+5f
nWzumeLKTTyAcGpe/l+b9/N/ZhMp0UfeObrvBrRBALHGszxrcJUAEm4X+G2GMjLXeERecPuiYDdw
Kg6P2ZxYS/vFrGu/xxPU0E2+NnBeh10ivRTPaJobQTCAzvZgybMvV1YdbeG28C/Bb83QChIj7v5w
p0Fu3t7RLBdP0LsTwH+no7K01QZ6LGxTxcNM5lxOcNKYHE6QpVfh8Au+bqW75M4tyehO9SGuAbin
PVGGYO5OPt6txwdGUX05mpriRXLkft41FFE68+hKwQHm1T1qZajKqTPZSEOIVk0hVk5BcZfumVdl
7wSh9igzfCOAKXhqk8IqS3rPQ9UzvosFDdd6OlX7Ve/NpIoozXFK2WmsnH0u4NGSg1lWvR7FrWkf
T+Krkrbc7FJRMh2tdzSE4235udB7v5y5fN7dqbG/YDkNM/nGH7dAgvGcAsURZttBUwWHPb1DrtU/
b8mOFjCyYLEMlXlNv3O0VYucyVQARwdFOjvrz8ZfGLTVs5nMlGOfmJi9usYxkwY8q7Xk3NLuh1Nc
bNmd806qEX01I+n4bFUDEdLCwSUG/AB1uoycgpvPEWEK/ehGPqC3bGt0C7KU/1vbNPMuQ4f8/Opk
1WRaMLJY14i7lBFRw8oXt+x/Co1L5a/Nxl7Sr5cSVSI5ou9EQ6ZwdWeMxfWRFDZU3mKEkTWrJyzy
MmNG8ifapVHSulr21qGHwi0fMnR95dbHljsXgxkYowwj2Yhprk6JM/CdXuV+Mh90KAW2u3nKvJN+
XhXbGnVPEbhTeldlM2vBPQVt0HRVYPoMNUVLOadNzqy+QJzrj2YOHMFWZ0c1Er3DkJ7WZeexOSxy
+F6xBQSBc71xyHL6StPZsKEFhXL7wPl7crU5tFZdsNCioXdMJLrMTbH4xRHz8rrJ/vpwGJeFtAtB
jOMtVtWkUZ9ACjfbTvJDEMrf+a4JvnNIF/5Ir2KOiI/zKyGmBAhup3N0QT/WxmxKa65MADwnCO35
4/Z4bheh2m8f/ez9xddRO3KDunN7Ab1BeR7g52jZ39o5zJ7MBmUmfa2Xx61tQwUojtwj/rX5nBmw
BxHTPCNWKyYmhTNnQQIdm1m6VG8bi0cC6shIAIoioK3SX1zg+Holy2gsOkmSWwrDFFDzUreLUwbW
rFCjU3uC3ShRnoG9ecca4Qg5jXNi0FOYu2Mc7pHsAAUMfLSP9vJh2/2sCkNup9zLXTlQcOUkLeA7
boF6KzTbUjtfasAv4XivSR+Cf1EFSV4h6gZm/JMXlfL8rRtpT51wjrhA0YnrJdKWJG19Dvvk9cbm
QArJhCA4Foj3Oq1GL1iHqsxJT9PAeA8qNNoHdqjD/A9nVKEkQnKok6ViMJ0mBuYpI8J0ZbyL5Mjr
xCVynfDTJPvtsU1P32+CtTSyvNus+cj8508Xg12SKv/9Q1t4j8ZVfs6MCLNfX1q6Zk5kfrCr4fuc
0/GlSDwTebsuXAh+IKP+13CAya+ROV3Whms/tz57QACf8LkCVDNUzthyJjutffRM/HafjPX1HNzu
Wa9ZM+FBZ7XtdI6P4Zu5olQ9Htovlv4nTGyLy8hY/Ybh+TnPWE9dCV+VVcbLOvzb5Ut2aK/eS8ll
cY2vUUp23ZLSYdvvAUNHYcquv3lrxLf6k6njqpPku79T0g/74J+s0NhBE8wS6ktS10ArI0uol6M+
3va9MQ5AUd86THLpwpg5pkgY/shn5RJjMzK6tZhmo1228nBb5f+X1kZP2DXJYlrsN7FYEIWPgCSZ
Bz8giqxjaQPHKml6mYUyWvg0U6Wj7YM7QiC+Xq8OD5GJqcWNPYRDPOxAqICMl4g/mIQ/vrE7EAzQ
bCJzAUNJNxGYHe9wkY+F6ptYXK6A5gPaImghzS70wNqtiByM9w0SUW1d9cNrMDQzvYGkwGzg8ssh
rvAMbvmaIoGki4Tr2rB0MuKQZExG/ZjOsWLEedDGPFyDKsfJA9rfMVmiUgJbVEbXsLlYZGBft8rM
TdfrTaKw5WXWU5yD0adS7HtOhoxzDuLy3QZ/PrKOfSf80eEft8bPn9gGt6RGa7rEFkumjkum3yYH
UOBFFQuoniUctWhiNlgidnNxZghtaJtMp3K/+yHYTIEtFXweyvf+HT2PhWpxTyHJzY+WbDHBPtNY
sD/EuLxuEg1r/ViHgrRDPouHhSwhO8aStlZUbOqvm9LNNFHR/2sS7mFMl7wfT6Vdtw1cwojgKj5A
CKfefNONFzMzMjG2nZzkhHWAZ2yxNA6nUI461w0Xto9tfSdAwmZCt4q4dh5S1s6RXXvA+xSnMIH2
Ci1amfGrxND0tQJWY3mJ7mfTTwIF10stehavgDEsmfzlPNhOZgPS8RCMeLRKYfSJR254nx+HpUFK
z/dIX/lGsoJ0eeC4n2dvEZo5X6ay8Yi5V2slQf4+QjaN9SldjCZPBd8uEJhLirBjMVaJBwH9BkOY
w0BNezXnga+8aWKzSEBhJPajpof9GjVQOfcYgAcPkYKysIhvCG5q/r+KrEeyejrNCqyVVXK8V+9L
Ym1HNJs5RHeFNkK866D7KZzpSVUmhANsHVZYlTQjM+rV2/GUBSJq0slQHXGAnxX6N9YNwmpQ7JEM
LTB74qYuwn7439Def4F5CEyuTW4ZPZ4Rg4rD2IxbS0cVKOjtp5TOpinJxHJ9cB75MKyehI2wzC5S
NSJK9AFxHvOJwrrP9RHeVL2fmhu7UElgpqTEed186VPOCtoabgFhnH06bwOW6fsHo00PJY2IOGNs
eCLuyoxXnC4Wh2jyGbjwWN8cDL/Ml9NmFy4pQsTaewRpyAadtQdO/RvRpKIf/xQCSeyd/l/sYNbP
tlXJoDzgYGghLfC8CRi+6LL7hIf9v871aOXlYK6Owo0c441SVZ+h2MerLDfkn8O7x4c3r0csdV1f
mL1hP4le9fLfN3HBoFMz1Xqc2/07lwo5sG+/aKkWsjAvc27HKwGksZum6DESWVHUp5E93uetBfk1
OX2LIO3Pe4g/FQsR3ifvIHwMJNeXArBXXm3JfRzFD04la1dcGIrXiByQz3is4IPCGoaGALErfbzN
2oKx9TZnMiFbl3JBmApdbjfZZSPwc92Re3/mB7xltpJK0qLkSvCIA8K3Rf88SvuGTAoNlbX3p2oI
PCoAUr75quRVgGL7qi8ew+09SNo3Fp+flnwPY8gqdQwyO/fjwBHTKdKBBPmSeYXUezdqNidG4tcm
XGAlf74Iqoljw+tgx1KvH0BrplP4TNwf66AjbSPLfJI5D7qSO2uEdyDGazMF9ClqmiCc0qKwB+Ft
gIPWakCae7rfrCEZ2VUdIX3hLAtfemIcP4P52Z8/pEg7qqw3F9CFDbReLRmvl58ABt98ohOb+9IV
ox2TW5e4TfovaCCRny8KCkpwRYSQSt8sH5qBKOVgpkuMLYcJlItz+naG8iHorJH4NdO9QcYLkvJy
x3Wu729IsvTMC1ZajUNHCVjr95nsVA7xqAkjm1D4KArDp+qqrgupQSEDIL7ynV8KEC0Byy0JT9CW
RGwvEYnDmqG5XYnTN0IIV+W6M8DxoQ5YjhbLVBmCExPwv3Gj5EPBlvNSRsGbiNzk5UOaw+0h8mYP
HdXFo90Z40XKmy5wguI77JrX2tZRXeV8v1UR+Pnq+mdvdSdmy1wPy6iBBL//2ARCT8JQdQZnVEXI
mM7UbI6NnIjpBM3+FlUYXSxoY7z5uUxD7/Oe4nYygT/JEHdHxkIbTEqW5mvGQSxU8AmuBCzmJ8s8
vB+X3LcQ3JyU54aibWRqXvUfiYQQeiPsyqsRKJtZjrc93c7HBFp+pjdZ8dyGrxrDDcy62UGQrkvm
VG2jq9Uklm3mC3+lB0u7XPwyfytd3ZNlJ4fymtx/R86Vnv78v1PJS9ReDGQcdyPuubc6LYpCAdsi
RZVMUbB63W41zKnUPtMjztYTsZAvVQkZY1AUCq/kd6ct0F2U7dQSMkSYvhgyywETcTDyDbi/uDXQ
dFeivuhVamAnVEGZV1T5y2W5kZzgDO6l/vdsncgcHtz3+MUmxhp+WqEGjHwAVVDYCq82XNATLX1K
GIzfxUGNRYh4Uj1gNFE5IsWehT8rBApLF4kmdXD8K7c5ioZWUfC+nvOhU46SBrTEy20w491R+d/B
8rvsGCPlblkLOxz09rer5j5UoU8E0kGqGy5wlSrRUC8hDxDqn42zfUxDekOJ7Y6snUq4/FHWro4F
pbdsW/CO3i9yvIgbnxzJkyKc1tetYPHKzKOdOdU9S38Ra4cZi8eOcOzPxai5kEStSe+54FXjHZFn
ocgrSiwAFJsp0iNnBDflPYDE3AJmdR9MRLrdt5N4fsgICEIEeBe/TR0ynI8k4ujgaLizSNouISy8
Pi06IgdImV/8kuEn7sxkQAPN6jTi2hTM2oa+xapASxWdLRisPPGh3MEEaTC6fGEcYw37eE/sEeLS
ZupAPq9Y4oRwH2QodRMcXKHNk+YXP/N1sGs0ZUN/Oj1js1Kl3+E7+iE5g9CLL0cI5TJpI1NR4EGm
ChinAG9lgynGa+ltF/dJEpkv9A0Hb6t9dFAaSmaISzlB58C2rBtW066uqY/dQO4LfDsiOQqqkocC
fpbU9R7S+GYZj2Lw3Dd8eb9ry2ac/5PoHWGz1tDq3CDruG+GD2CZU7QKgYwvRxQKFAZKLHA8LG/m
htwmOL8OwaryOC5GvkMqHTm0UMr4EaDBu/sfsCC7S2/dbS8/9lZ27yUqlR3SKPWzEQ+M6yELchfu
vfabKFx4gv98AWh4fDdd5OisX6tlqrYMa40/tUl/0pTKPFzCxQe/+yH+NsHx4hCsOldKOhM1BRHl
jBvXXt8sv4zzbGh23QhaABct8V3MUMi4tG1k12UZHfRV5+INE/RL9D9yxPUMBwEcmERI1AXhNI8o
r5INAi0L2nBZa7vSkqWS4ckb025I30fs6NEH+4sj9ZOh+Ig6E3GNghjw8GPp78uZYKVxntyjvgXk
/D6r6e6NPzBKITCHLmCZPVGT5T7t3dQlhT/6iBx+L8POGNyVmdkAhEc+AV2ou0gXk/CMQcHqzBlM
7ZXin36H7EXB93iyV+DDi2MtZHrvxULUCJld0bIrqWeIU9FeEkin/7hC47abddEQrngA2G544vnJ
nz6KJt7QdoII8B97v61tgYZf7Egf5TaP4Y56GgLSM+SWeryOMiWaFosmFHbuAOl3Dlfxu277S/6c
WTR0Yb401jXyAs8DywFtwDJQLI4zD0GgvqdqGxMANEgBniQfkZxK2UEw/S1+hI+F6A04uyNx2/Qc
gK4yImtOnln5assGwyM5WvY5A6pSAPz0pLziugCgokZeSDZBCrS15BcJt2RnEClP6M7WDrHO7wjt
0wCXw4nkkPW7OcSdOwEa6n3+fAubUjEM+0Vm8/+mTLnAhIorjiHMnuoxsizgwegattYtjhwP7wDp
RamMtsZzH7fQZas6P6KA4WMtwL5tq5CWbP2H6dxBg0yymCQjsR9EnAHVk8rM5EVEqwmVr420an2f
xJj1ivm1q2L7N70Pvo4xzDC/ghfFv8B7LCQ3BdyKZnGfmJzCVuRj7Xcjfqlranvb16ZV94HG+l0l
lz+BhA10oWjsRU6Mm6Nmpgk2KqNQ6/2yxI7tYIcXmYPcMDJYOne0yrAX0+kiiRvDwwDXztl+7w5I
zKReLodJpH5UhUPxJsVQjZRcBd1LCPvFbNCdKBSePXApEituGjrxFiFUKKksA7vy4eElvNpQMQUS
/frROWv82O3gM754nCKOk9xhJn+U1Elxv271p6IbEHyM6assz2xv6C8jp742nfiYUZmk+Cy9Sl/J
AboQlgQ/dwaSVeIZACzlDzrJlyIW5dxnKLj1v+jIXo9h3LJqz0zq/kt0qKg7npe9Hqsvohn3YBr0
AzdnSk0vDFgdask7KmgK06bwKzGs7bmwrrnmsgZhqZihd/H0Lz8uwL141SIW0bUAUO6E2Lz3IG/X
aTLXCbhOgeW+8JWFZUhND5z/Qgd97GNkNEBV/bmfeHV/o5z6YV8jkm0uyPwnbfh+F3V2Ywjhsy+C
Wg2M02n6h9eINwf5ricGoP900eQ9tLnsG44uUB42fQvcMaOJ1FL/JAzslffYxjgOwjk28/Fb6Q+x
Hkk5W07QKsIgFAOOH9aCQvqtB3QQMDLzJBYZqzFcLJ5BPCi8XQm9ZgLCxdE9cqq3dNXXgGxdtwQs
Rt8fWAT6B3bCBzcjc3gwTNxNAzrDvxZ606CzV5fCIFeiMuV9AULnHGqtMlXT5XveQXq1HYd1IdnG
ZKzCRHFT1FhrGtv8UlHw0rcYfvQTh7QwK8jAjKeRJm5ENz9kAB/o5PY9fAsl/IhmuWKoQqim3P4a
qtw8QRm3S43Kud7fyoLByxMv/XWgCakF4uhT2CrasvpIkMZw9x+YVdYt2Lhxy/WG0RzA4T+XOMii
d+XmUXpAWLp9jlXuLkE3Xh2PrQJ6QxxYU3g+dw+EVHbpvfzY0h+/DSOilMbeM5M6u+RX+fx+0XIR
IiAx3E7LdINTBGKOzH7R8b6dI35z6b2JhO3iaP/eBTzbGbL/mDa1G7maHjdQKnNFxNBJ9DZNeQoa
4s/HK2m6uPqkgXcgDIFvBxcrMFTeLwQN0oM486JIrs2bWDenj8vZs2HvlrYp7aiZmezE3mroTsIm
y+y/gQoevnuNGU4FYmAvwWNtBzofuiZhHFRGFFDvVbm/8VvwgcdE1L/yBWaTSJ/Vk0gc+pxzx8+r
txladhS6vmORAt9YSWnuItfOFt9wZK2XESus925V8G/cD1Su/aqs6+Z0APLFi2eqD0iUG9+d2kdu
M16u4KezVLaUTlVK+l1O7U4WiylRzdOp3in1UdcPeqpW0CU9R1dea4cwMtn2exYmk2Fa+fSZ0HOs
GkfHg77Hwd6B0+6bwj7O/1NocDwA9P3bDmGmiD3dOSRJGVbc4OUgF1IluFV7OMEjj+IufaiBN7XV
1fBVL4R+0vfrpP5dbOQ4JGSoyDLPMqxXaS3bK/CaUec28V371Vm7LKNhTx/v+t1R04blIhaqZQEq
UTF5Bhjs8qvZqhzPMl+vd5T7xKi+INpCnpH/TSj48rJS9O4NLvU7ejWHGVb23nxa353MIsBB6n85
tE7DkvVayEW6DhdlnqS2t40hJtnt3Ah/zSzPvtxFPGxi8Qenv94cm17CFjFj3s9Q0S3hQ0vHxXIQ
nl2BvSiFUVmCGPESxuk9kU6RGM9rUuuoJpYB7Jvme30ItRzxUt5uEVNGstmUwcUuiyQoz7aide8h
2yRzYuJyXNu+5UodwmFA51q3U2kcna/TYrYFL7O3Qu91/oicrGImE0fEys9UKCNU13mjHYLnY2AM
wuitUgBg3LET2GB+qGfwBuG5UnuvXaHbuu8axWTagmo4rEI2sAwEQqvTw5hEFtQTiHlmGHtnnpV8
Y2h+3Lfd2+OdC30klFazFCwmU345F5h0Tx8RqsNrYctr1uG6s2XjNkKdEbjUnSjj0l2JMuIulb2X
PMAO/CoFLR+UZfV31I7BFOzhghRzIo1cmo9KxmZ8zP4cdoyW8YDmKEb1vWeu9VEh4vkO2wEpcRMc
4HCAYlAwqnUgEKdDdksBEWo390XmobqPEjFYopLwfiC/QitXcyXnsk4jKFUKKsiEqcun5Vpu5F9B
KL/DOS9FcedqnTYdZY+KsyCiZ4snTMea3yEsYyYsvYdJ97nCKgCzcX1t+KNkjI0pmAeKT72kYyhS
29VEA6ZMY1Jli2MyqdvFsvVkDSh4Qg2mICdJBTIlxN8fTH7l30bwtZCZGFYq3yzIywP+PReAm6F7
m/SchctgtT3tiBakRLFHcjQn6+GlJNmabjwFsICaaUmpuoHTcyRTI6k3tfktLrBqix88nnKMWc2P
xK7WPWp2Pw/sGUty1eaEyyHqQvzxgejaU0jEJCb2IHvdvW6oW4J+BcgG/PVF8+445qk+u6RDJ61z
oPEKIT1BPr2rh23HSKneTLp7NL2MS/Wa3rVApAEnqr3WfwI6rOscHFItErNwFqL3LmA9ZCWmZH8+
QVOPBhJOmHZ2JVblZtXnRcaNJqWGxhZD9rHl0xzqboVbt4+yr+z81sGl0WGLgn90YQQnIOADaVV3
hTSxFwlLA8wKm48j2paVnCzHHiru5elPlqW3zJnLYLkGB7cZ+AaWFvDnaa61N6SKY7rSB+JagZqM
T154yX64nEAa8EPKo9IS0xyQE7AuvSVicZoG3OeJWu9cwYsEAKBxXoT9FIFQn1swmvpvU6aeCGFj
+DuNFHvKM0HhqdYxEgTQrTjCqYr2qakSUcMOvycKPsfqFiQEjFokNeci7jHO20wOiJ2SaD9f1KVz
BMkXbu4LQFVxHPqFrJo/fUlYPyzdV1QQ4tj1xv8IR8meA45e9m+NkBsIEV4sv2KJf9GAF2Byas2W
UpORs+bT9gy5ctPFRFp0xJMDmUmWVtTUrL8T8kZcm+JWKOfCl3yyTZvs1U/e5KSHKxOj8zU7GgSD
hyhnVH7jXbfZs4Zg4aTClvHGEx6oTQUsCqjFosGFWlmy+tKeFca/3Wdz3xxU2zEx3wTSElcjkKxX
U7kHAF9ZzeZFz61rRFvgdfGDVgV93KrmEH8t+w937Tlu0I6p0Wkfukuq20hJvyng6dLyoirscpG2
tISfWY/gb8hcfCiTFHTMN2GYKqKKE5AHb+KhyRc8y3913hJ98YvnjGNh1K0UTfvHCKPFGEBt931a
myovDWhb9IdDn50egmgCIvsKzYxlNTZYBRDtHz8DWNwBglqRgDHg0NTG3BMpiIKqGP/qjhz2Nx2y
RdCyRv72mzuReDjSa9wig8YKm9ErZ++ofjb8ON1VC7t9l9yWn155PDLO/Bnpjlz1kX7mkXS4lRR8
jHwT3tcm4FFIDIHB39w0KXwAFUA9L7b3rOlOviGVZYt47rvGXmmassXv8QYW1OUniY6Ssra9Y3j4
nG06vqTU6iIacYfbxLm4Q5bmQf0l+KyJRqnIA528uJyD5aNGpbPgl3tremMCoriVOUHqKDev6qyQ
uOorJzYkODBYgdnHekRWFNVian8mOm3iMcpQHR6BwFXOY9qoQBomFk1oCarDfSehv8XY6s4ERjIy
OIo45UUgdd1qqGoRZs3t6/dbb301F13b6xqSPHgrTVwqHqOohdbK1UV/p2SG9cM1Gb+ZE5c6yQ39
eYlRmUBO54IW5vC0E9V8LMuxwVMMrXFYBaV93fEaSubkTIw1Hn04028n5Qm1pMuYlh9W4lBBJ5NP
vE4IdgnHx2qKaspvxvCyQzojYGhwm7BFZsVGgi+GPmY/ZNGJxhtdUR45NDsLQRPvZ3ROTZ8qmszA
EFwJBh8kDp35WUjYgkq63aTYxB7Ow6qnb08+dcJea63XBnXvk3c73TjVRpGHZ2wDrhzL6an7tFE7
B19I5ApVryvu/aNh0hcNemhl4cskZCDO2nVWCEp4wOOdCIhDBiBqQoq3iO/tszG4tQVqHhDoC7pS
R+oSyqKPF14gNVGsNCslCamjD4koKOV8k9Y6j0hStl2/XjUfGcCrk4r0gTXkeRnUnU5THp+5rmhQ
UlCDfgS3oF4rVYmeG1Y2hTwaD0GSjNUOY9ZLPvmh5OgAqs0ZT4zt2Ea2aBmpw2BSC5rlM29Gc40/
3vFcRfYdpXax5OYRFmXu1hbzEiUyfgbFATWMPBQ7U6jHtKrJomOV162hHuzueYM9hxMbh3uDKoJ4
9X5ABckZ0E2y0x6+BSKDmXrdIISXBWAa/oB/y1IqhVnR/ASeY8Wg115+0Sujm11TCOuCMxxXnUtv
97ObR5i6hXKfJME7eX6DjlkUpH6DJSornqoOI3DDJm2I/KOvfiZrslbUD6QyFoyKXgFI6pAVJ859
StNc/KpRmvDMjxD/05egS4ziSa98M4vtTVyA38qZp0kB5gDPeCG2933x+ehbDseogg90CwaYWGgB
Mg3JUX8QQfHiesIf2R6GWT3JGbVbLaGUw+MM7hqLKrJH0iFeR32ParOmNfKlnAMAAoPYFqe4tFwk
ma9x+P0hzQLnWjOpjjJGVc0QcxkxyBXxfUOtxeGwnnFIiol7es23At/sdBjwhNsg4wMAap4Kp5zH
abZvWXW7im3pG5sJ+N8y9/UVzvONjiygQ53UqdMhxpd0SNaJxVPNJu/JLoxG1rQ+sRdCJy1EzjUG
pZ1uxNiGDu3hoUncssSOtUXRXlgIJYwM3OcLS7JgKNM7Jlqi1fWjj6gqQhDoA2QBXHhxvp+aFEKE
12fSFzzJlMvg7mQUt0cnH5E/nX8SuU4VldrW4/ad5m+mcNOSkRra/yoZOgpU3yIsWZncgvtz6ZYT
Tg9tYc80BDSAxQTR6TOMEWyV1Szj1ziyWtTNZdsy/VvTFC8HW3yvaui/12SSFBqF7aTXaejWVmnB
QcvelbVMQgIoQIo356NY5IBlaHNgMh0JtMy37ZXrtSUVItkKfq+xZ86gmZlNdG1R3AjyM2b40DDn
N+7sQpJRfOBfM5dfdNWHiAuBfhFxis5DHCvH1MqHun9yJFvNN3yTBdR7yRZRYeyDkZCz7arvgQf6
kMwXrpceTZzyqwyWBhp4h7VyQAiH6ebaRbh+OFZoLW51oq9+EVoHI2z4FC/L51cPwoUqjzK2kfN4
cIbPCrJ6WCPUIeTutFmL5Gytkw0fhLor0gOt1v7n2W8mGFTMhuK0saG+O1IK7KMY3BkWKpcMcj6H
MHfd7BBV9vCEp7a5QQV3dvpgw3iaKoMRqp60FYN/Ykp6dmsaLBEwAGC27n0byw8oXBZsRwe6W3T7
4ps+ujo2Fw6YTWAsH5oYp8N5SkN9C4IRau4znc74hX0CVFkh1jIJzTh3u/XjMNfuZMildHdDGrqR
Fn5xWdJHzohRPoqbC6TEIc3fjqKcVfX8UfA1IuFdHJEaJslbqErM2cqX98kxlYxfQ32ak5u9qj1m
yYvBAP+fq4p5P6dyb+YnEwiFvv2TnErqvD23XH8Tl20pp+bqEeuMGRyCal6s2oxpZvpB6ovptlis
4+wOOG1OyHlO8IStKKHKdm7+k6g8FVLSfWZlZlSEa5ner6xP6fXcb0YmVezm6y97F5jyUBHQdjmm
dkEeD+CxYqcWxUn8uhW31BArjgPqmiJqhXwd/DMeK32sU2IZFyFW5gQL99SwM0hf6jTNEoGDz7W8
+ui7/kzmzPlA+kwZgSay0UDRP5lnO49s3eghoOQb/iEqcAfO8Kc/EhlcKkwfqV49erfiQTBWIMkR
monfl5poTLvaiSN5lrF1hFCN9ESfBUh8PB2V2Msz8PDZSWInvDFs+NYW00sNMbuDU+bqJRlyDPG2
KGs58UL/VGdgkGFc+BvssdxtFMizrYjZ2MLwmP28d656gB/ellK4PKcxrDwlhUWZrMtgs/oD2ltl
zAHThxgZW+pWMvvp1b4bxaDhsk69GpROUcd2rYTc30/guHbs+spU+fQ3JDr9fpMW/ZLcKUMlnhQq
s8UykOeboTaayJHxkNSqpjEg3Rr/lLRUPLSspbBZcW3cO6kMRefIErzlc90FdbIbngmLf7kP+mM3
DDZcso3jJkKtFbW88cwta0LZP4nsp1U3g6gmeQt3O5zv2T7GozpxHyAMMmg7PuY2mZKb+ytBW/fW
zPBQ7WRipcY2cbb2sTSUCRZCZTVNy1LX68aXqYbJr2BqwgancACevOW2xpufuJtGxOyD81sIbMYV
nSJCCuBkkWB+criHEPFOdUiw9OTfMqFrGZy+dnIN6GMtjlT/7E0FCFsACWZ1l0btD6nAvYlEinNh
Wgawxmo5KpYoxtcaAExrPUui2118pisJDQ9djt97kg2IOnCGW8QigHt3GuXE/3zYzSMzykGQzXKQ
sgvL4rABAAPkCbht6sVjxd5s2yteqpoHd3UcNtWyK7ekJlJG1xHfZY5zHa7VRvQESMKokC4r5Kzy
mPXa/U7Fkuo5ldf+ch5WO7eAcjzzT/gNNBcsxrdrJJHy65hTDym0LG45geZIefAC1Eth1WkaFb0f
iQCFYe1WGLAAdzKOtRfPTfJbHVMYYBwIrBAfHgsfaFOllPbb3IkWol8iifFzQ7az7SgsgGEDJYmz
JgsQDGT4A9zIr1q7VfoyliwuCPN54tCUYoKE7a5tLJ/j7SsX4EnlM9n5QFnfgEU/DQp0KQA6IZQb
fo1KqKyP48M0aGTe0VwBeUY17NMoU5Q1cLOObLq0xpWA+qCIJX/hyKSOeR9DC5Ga/TOccGbKk/px
ozqDeHYgbV0CR9YmX/o/Yp8v63ZvrA9LqVaUYVGgMhaEajUg6Elbr3YtlrMfv4fI5sNjrkDWrubm
vwWqBHJnFypmwerCFln1IGV79I+389z0CV0W5/jHB1Ebz7TN27S1Jb9JZjD1XoWeV6dassuMZMKc
VDN/qOkQdxOmQT8JcRnhyD81PBVuJEAwk8Y3UIe8eCncdtmHtXIg/toaI4niKKzAScB2+ieEGQ0X
PVWdUWBuO/C4wYYf8MgPchXqZ+LK3Y7e/0yhMXXspn8tnnJczH7zce9KKV+O4Gh6OTgYT5RAupan
19VjfuODPgaHNFavG8qxfBEcL2D/TcVALVDJjsl0mBhTlCCed1whBz0EP2DuzMlVfQ1taSKRJfMZ
8r60z2wwwZbLGyxraelh3w19UhQ6kJy0yVOLjPC5I9n4Q+sZfTQ3pIAhveUr9TDk5kjyv3IQih0C
e0tMTyE58nrPI0iEdlTOAc88a/M/bXr9B6Qpac6RyNDlt2WieHP2CQMGuQehZmckF2bk3A8pW4cT
ju1op+px2PtIErBkQ6LacAgoLRe0Mf7awF0+ppCx23XalKIj3L0eJ10t3HaniDkU+BIdOTDF4qgI
HZ9BX/mSLFb6fehdpJVtrqCfNBJ/yyO+MvX9D5O3IB7/y+5+0Wek6+qpMWMD1FQnFr6NHeBkUlAj
2yUKMCEVOa0ZRCpB304IwEMHRKHzwGcODRUjkkOIWdVgWxqMfHxXswsrxKD9kEExdPqd8x6TICIG
Y7MfehaIRmvmYFnkTGPw+W2Y4yb6D3C/ceoPrpWR0eeu6WXWU9d24dcCf3LSIBG0ozXLKFtJtJ1N
FP1Uw19Ld5UgiGtarFzJd6Aha7Wdc9Ucyyl3GkX9q4+RFokJLeeW7unhHAc/uYc/XbXjuOGGk2nj
wVpdJ+jp18m01h5/jDoYHx0hm8Pg4zzW78j9EkKMBKaogqnMWJJA9ND1ao/J+3Y/i6mYFxeFpfcj
mXCkuKK2ELnTAzah/7Ezj6pYL31M059yzu0TF2OsJ5epw1HxsFOsdJZQoaVzV4GLDboPi9N82g4K
wodVwui/et3O9ppWSES0r2yfdqBmIlvCHwYM+7L5jJrXoAdRH8kn0TNeZ/LEwHpX38SGJfsu0VpZ
05j3uXS/YRgNTY07Cx6A6k7Iew+1YHcrjUba8T/BNc90vZc7gJBRF5aE68s+tgH+fsR2YVY+hqtF
hKD/UXNaAA15z+xYByIW7cIdWYwnVtttnIc+p7thLskgcL7pesP3bW79cr6nLnMtVR0KJT765L7Y
HnT9bI7WaYLTtgCEb7cjXCcRntqw2rXjsjjk6O/wT9p736bF2s6CBVUSCOqPISNDyRsouy1CgMe2
pk5fs/SpfWhbUKADIzlf+LGniVQVBTTPt92k+drBBvuM33VSKnwaBfY6+fmOrqImfJJHn70bdHdK
rDCohcudOgKCQmYcFNIyFZzuxXEmrhQ5KsXPseXSdCiuGEmg8ruGIMD0FpO9PCuNAtm+NM9XzIlb
RnMc394ZuUOfT6eEEHkk5ItD9zhIdYzi97IIbUpNQz8XTNSk21uQrAd9svK67e1y9t/zw8+Gujg1
FHdAWZoqdMP3tMZzrnwLHf4fkGM2zcn5dvkeGj82XLh6Y5cWF7jBXVxym2TYeCYMbWtpzYH78m4k
xOKZEQQy1dZa2OWgksl47rvekx1eypFJKWNJO9mUPH8ZNevBXN6BcuOUi1SoJVHb7PdU7hVwG5UM
2zzFwPXn2tZPq6i/nAXiTQe6TLw1XIJB6gK5oVBo736sWaDCUwUUZxDO/hJkiP45LKrCn2DkRDG3
EyDMHl9+VgXplS+e5jftcmkGhK0Hf4svmp5o7mQRm08+bB8W4x0cHLenUXjKLBpZCs98r36vJHB7
bB1T9/EwERCQb72MgDSY/mbDFbAsCzE5kMNVJRjEcpn3+RYP/s82a0fijLoGwmC0eP0IE89csbXY
cb+spsaDTtPp89J9cdpUSevaGudOX3/2/H9I+aRlXpCRkSvxjKUMupx4l9McsJWtVaPYGvFrni5L
FGnrRGuVZ7UU+L4zUrLQeUof/IJQXsXjkBzSAfhYd+c5UrOLZa5JHiI16G+MpKuIPd/y40MbYMD8
Ljry77zlb6LS1jCnfKYSbPI/+knm+i+flwkEvLv2ZwFRihSSeCMPaWP/qXa1oHEzgkz1W7Hcoro/
AcvNixy6lvbUf+5HSQ3IgFElUz3uzP8ApzQv1bbDnCAHMFyydy1cIP+KGY8oMwogCdSpGftVWYK/
r4uArqZGw7HxsKp9ZF5gYdy4rkKVOT58ZYDKbADMKN0pvaJCecycHr9EiC8VCFzpreooN61b6yyS
K7aa2EmBNMdTtv/XpyVfR9TUztYavDXNvqLRK1U5/FT455h8l8ELYzPAfZ34xGk+uiKfBVFACPL/
GROBm+LYy4pT4QkG4aX9XfgQmyds5bY+/xVPoidGNNN7t1add2WY1kzOFc9fvv7NrNy6sn7XKySz
VZieCvVK7kXlSCU85+o9GigFbU3lGfx8p99FiPptRWih9AvrAbToaI/2b2dGN7kjlm8WHAMckA7k
ijmrNRRXLwvlmilQaVgblLP7nJ2PQADVKczYi1u6qmjHLKTGrNuaPAZtl97MwsktzJRnMn5l42Xg
E2FSD1vX53llA7yg1/8goE9Ulvf9g+JYGOymyziJ0bully/q9JYLhEprvak0oLYornyH8nvD5N06
bF0gBkO/kf0iTdTJCBkox0MGO+PhRa9nKFvmZ31+nxfZHQLnz+XPrxPSMDplKIkUCI4HRnu8hoBB
cQg5GbISTvI2tbxvXBSMjP4SqsP5jIg9EpTT3GCBKr5Yoodnqog+yuQcQHICnWc2bGhu6830r9VV
SSdKIWhmvzJ3IhiBUV+6CgShRkJWDEdYR/8kDLOp+OGIxJ7stJFL+sLwGDutPfvIN/yFB0r4ejcY
NLu5aJ9RXWb6gAnzqhFsE3jh4l2Xqqr4KEoo1n/4gs55dTZ7SKVAytUYLc5XpDbaUAA/XfXVb81X
UsfP9UQEXEfxAwkPso+Gs0zPBBALp94faNX1CqIuBr6CiAYRXsTHFF6DNi6ndB8PZ3EhUnTUdpYX
LsircUido9R4Qq5NIWLN+w4cI9GnkcPun1UhbMfTnVBy/egUZU0hZnwLl5rseepn44lY0XuTYEHT
JmFMcRPh+qe1zae441iidGqIvBRmSjYeKrNq9JPrTe7WC5jKOe4llci0fqW00yzwCtUEcV2DK4pm
mMOPHE7zs5ao7irKtBEgzl4tf5iU7hmuriXZc2I9NJ0SA71h6tp93uAScLP4QYj8d4QdvHZ3wG+1
lTCs5KnvpBe8sZFlvKA+k6qSNDGKG1Rc2kWvsOOL7OhkuHNGwwhxi6HoK7rlpuQgfwPa/ItPqSVE
W8nUl1so6X/L+Al/qV1VZuV9rAREuHtBFBSh3pjQ+3KxF0D+wmA2UfscGaxHGYx96nTCNktywKmT
eaF+GKi9GlAah/5o7S4zsrLfVtCsZ06QwUyiGPbwhtEO6R+Kr55qmYHXsQZSL3p1tLt6Zaz+EKK4
r6tVOpkcs7d55j2KwI/8MJ1HoUjbSLBFg/V3Swfae+6GC0LrodFjqqsK1xT6dN7Q8XXgssnUOWCe
dWrpcxCY7VWubkSESeVTDsXKA9Cr8ioW625MMSssWao3OcyC5xw7sptwur3QgdGCKS5Ga4fpzo/1
GIoxo2BhenIDleodYSiY/4BeGLzgK/iVPTaGYesuBiteWr/vdaCbKq1WtmAZ0USLMD3+3+hPVEjk
Pp9bOmrNBvHnFMSpC7fBD/bMJRlhT8TqXM6JkCQEAPxISE3rzCx9LgpBT2rt+i+ey2MaK1O+xBnp
TKHwuf/DFcCOBphs+mRpHg0z+URmO7p6jfDcMihhuLPKlzxMs1hmLj/wTRRlUl75ey65dOg44lRz
0yaV9EbdDECywLE18+f+WcuhfYXk/B62oB5EA+XVXNRha8BycNi7kmViP3PSYY2BZK2Wz4ZTD8FN
UkDTub2XZeCEZxcJhgbdwFC6AQPN2iWcGvyS6UUzhD3h2+JkNIKR9/eF2hgkFlAhzdhrI+XPdHiM
erBZinqIKO55qPyIl0w5t/DOk4T/J6/UUIKePh7XX29I9vr3Fh8apGIwDuPjWAGMREpuWSHvsCOt
nRI9weIz9Kp5l1MkkNMBIyDRgDwr4qNqwxpRZWThfgeWioHc1EPhJoBreOQkoRcVNYoh+Qwz+TUb
oErMfupUEbDzXyCV5QKXgSli6ZswezSeZ2cmyNe8fsBb/jahq+GJh9wV0k39hV7GkwCGQrQRSBT5
2S9AfWm1UnxkxcadyMC44pWt/M5Q5Ke89JFyRSoHfaXCj47cbjh62oBeWL/tAK6pu+KVz51zUzAV
b5KMfEB+bN8d47hJiWHLRz8sofUzenoAe6TAwKs7E0Vimj/x9s2wygu2klE2PDP6fjQapPwuNmsw
NKvwyw7ycMhXsrVaJU+Yv55VIEMI8/KISkClBiW1+MC+K54DkfSfMDZTbRcX9HcVidhGBhixYDQA
de3IsAZWbrTA0fPZL+JGqOt5LeF9I/MZ/RLvKIICa+Q0Wk3xYxC+gYUSU7Xw/rY631FCtl6s0OPz
bitvsxHvKcntuXNbzqh7EvYBCLDdk+oYTjtOtKmOdSNXv5C5hsIPt3DFWvnyS2yPr/ew2Tm4kbRF
qogngaGPk2ahceIQtPHMMXIDpWS3qPnDibI2gtVTgXh73LsTVUKMm6gTFCEcCTSn8UfwwRiWKMID
L/MEH6SVL7I4w8W7Dy1FUBjifPRJEJhkLPMgsCdPDjM6uq9SjPLpAmTvhgfsKSoItTL4/5yFSoIa
BVrYBhOaVrf7RzglqkIOV1CpRIdMgXJWQyFCTX0AmnVV4a0yvLa/13nT3FrLjM3hMaPcQHkO1HRO
TtdR3kmNv2beSUuwDpmeQ6eIGiQUJZBeh4aDrObL0mYnKfS27fv+y9ozQb5c7rGFOPN5JP8il1wi
CV5ORLujaBNVdzFY15/EyywCW1R7agpZ8cHv3qe8U8veeaAww2HpWh4x/AuvUwUcns5qBQJ/AZX4
4v6QYsN56swoGJ8VT54uqOst6fdE0TXAzXnEdGrH2XxxSl1c//gm5CbmLfYF+Un2fHEdxAA/3Boz
t01V+BqH+endzaYLBU2VYG6OHtcv7dnIxvjbhOKVwG7CVoDfxMtetyf9RtKvUmRhF/+EYHQ9VI/b
X0+t5IHBPULmrmKnin6JiVgPQF+wX+7kN1gzndozG9RnnG0IT8Phrm8NCb3wn7yLjNy0yO3TukdN
rfmWPa9/IDsa7GFnp8qFo/ZT3id1nvXH/ylRHkTul7ZtDgWPSHgt9NsMueiDTyuOdvXsG7SxbomM
/5oRhIoDtV+5LHmeXNLLBRvvPBIXgpOWlzVLIpNltb20INonGJEQnWZrIPxGI5AnjL1RBToNCru9
iRsFvSOyKlG9BYalwtwJPrGze7KFtrrEO+MiXP9uVvmi8ov9OxmYjxY5+oEDztu0u1fn4KGTW9rd
8CTCfcXzUvE08L0hkLV5n/0EVJ3AJEzcCXnVg/CBiZ1I83aeGK/VSMwtYJ8nmOqptLAc3QmHYhJ4
SSQcDMm/mhkddTAmm3lTrJs4nICFv5H0bKechG67Srv88FHtPpgO6XSzts8ZF71HjP9XpGUNvMLW
28NDxSZ9dVwsEW4S5wMcG/et/nuE1R4V9RLsmEBvyl+LfJZiFoD+/8NYY9ZSYP78h86pYcQd9mht
UD0y/a+arl3VYM3CYVeNLYDvNKF7Lnw7KSspHLPfbATFZ63Hy2laeEkyxaxpqevLP4fBzLLn3MAr
ep6jomx5TnlqQUbv4b9I58GeVBqVFYDtzaNrcfm5+mp2F7zQc1DR/xRvG5C46HTp7ONEv8Ih2ap9
CV2w+NXNK/cztI63663Npuiq6FHg6yL0lwZ+xS50KNNc5cR9nhOUjXO+t7KRF8DRwoMygFdF0mRI
TormOClS93dHjXImcu39xJOv1sr/dLCOVDS1PdMqbJz2xMpa5sxq17mBsa8/3zF/UYfID6O2CSsy
+cLrDi3Kv4mZoVas7u4s8dJ8CMR59K0wvCaD4gIHo2lcw/ipyvupBLqf8yBgI49hpdVuWi/LXbms
OIoJwWlUwvhAYYaHSi7P259lwCGQSiAN0l47LEC3Y0H09m8pj2vSa8EdUMyawGEONBpUkprEzJQt
MfnJ7QMrQVz4gI9juz0y9zWSW65v+l3Qg7Ak77Wblg93ssKzYBHWrFT0ZecPwIaU+1ptf6Trzz/d
WusMKmgVIdWm+T9MajsWDbkL0xTSCUFMWpQSSld/InxBQ1e3INJB5yN95WF1+0ROopGRmS74Px+D
TO4R7k4ZIzQM3HJh70VgK1CnXd0JZZNvX05yg9dUp8fZKi0ko7aeOpxrhVHVIfDceXmD7x1aIZod
c5YlR6mzJnpFEHDIGD96+RwcBUnb9KoFYd/x3stp3fDs1HUhxurcV0sw3jdm5C8fRU6evep6k6fa
nSy1/mDCej56MNuzq2772+odBHT5pIhngTiL2xXL/eWIT55uhFzj/AqspdMCDtt/WMZ9G8OdAl9t
UJCM7DocHDhAtGB/PaeBZcOtcxTZ5sOtddjn3oEg9kwi4E/1ReidOodIPGPWFPODMFAuWMjfJM19
OU01NCnzCHxTjkWvWjgPMGGi8qdMHV3gTOy9LQNuXgDVLzkAN4CMWQXiryxTJQfv6slpK1LkCjfy
J/OlTy1EIJX5+IJjiRoj4gt0HgGk4XiDeKdiVAhmLMnSQUlR05ykraWCDKhXCQA1RMniKunZYtO9
d655Dm0uwf7GtN5SrbQ6zAeCOBVsABBpL1+3MJFGOpkAewNOvFwx9ZantnWFrbqDO4Gv9KyHAGhw
J/+mz8f5xujmagojR2gdratwlI/Fn2Zy+N9aaNfDybm/GQMdUJ1MEtyN2vg7udljbBBNZ8kCV+ar
k4Jwe7I7p5BIxM9qE+DCvHt03wFhCX83ArTA1hHw1efqTTDmydAy0rXENWfqk1pU0qwp4uhdDGTa
bt+FFB0Rjb66MpbCzu2XNdvUocjtTImSrI0ZLT5Fy3WWnf+i5AMQq4U/n5y0LqkESL1JNz8/C3HV
5JI3xirr8TsO/LrUji9SwU09O8RN8KQcZ3EKNCwXi9PCYkdtVQPyLkAxSzGbPBgZNJ1XppPFLHjM
YB6drzwHVHz8bABsnVN0SU8Bi7nKdws4lDBiP+KdZoPZi6tjAG4pKBY7bYfOUHyPX363qGsJNw8W
osa0td2NqqdmY66BnU3N0IIFiZffkyoFHHxQlz31G1duBZm334CN5r6//15sYuSlUGtg+XOOBMzK
uBHJ2ohwKendtWthh086a0mOonQk1nC+BIj5mmSvrfPn/2Cz3Zv3RzY5yQHkh/jrVIGs3xeJTtOt
x5yl6YZ9XIhcST6t6xTJi/z5akdFSAg7XU6K5FxuNiV9lj7IS4ZceEjkeOoh//8oAjKi6Te9K1ql
rfXFLiZwC6Umn2fugnWhNauTRAntFvBVU68tdproZIfJMwmfD76iTJ1cS5XlSPukPZcAkdabEX1j
u73cV8jFgizTwTwUbguqN+c1KA9EbDYL3f++obP0GUWMuGTuLqjF5yOtTcn/wvwFLxquhUov6KU9
sCzJ+P9NT2Vv/qfNmbEpqFYEcuclpzaC38iqQOSTJr+pvULZpgBl5S7uuHdVIo9LIIxEjWeqi4kc
qb55yYrosur5OrZA9LGxpBbrJJm4kX12Zljq/OwNAJlHlURhMkJzc42afkyGj/ctj3YWXwwturzA
jZFugMyS6IdnNqj3N+DyHrOg3IfkUprzMbkwXI53qUK1PjVQh/LZ51T4WdnhESVmqBIkmZGOuu/S
29QtUlhK7Wl+zXsIbAqESveC4dPaCz3+FjasWaBuGOavAevGC8AtdOTfnfdKtUhBgy8weiVR7yKd
XY1D+7LmNj0cbRz1qLLNmimnYYvsU5XIgCmsX+nAvcu/1eKiC97y4cAZmxMB/VjGwUTaMezMET7Q
j8A2Q6ABM4x0YXNvMZJWVCJcONCBaDY4dLnyvZQhWgizIXOVaNt5LFgCJC89/6PJbNLQezIv1qkD
F1cQEO647UJZYKu+ptU8xKyT7Kb+3Rxu2in5YThWfhqsoHJZ4Gr0w2XwOZbG3eEKxdPzEHGcy4/5
grQtSqMv8m1JNBVyAw3RbxlqWOReOow1GsQrJ8/rJtjY7C7ZiYCFuVSOjL+uIATioCpxf5T3H8kQ
OBerkcmi4YF8mLv1A/8Ye9eZdjij+9TIKyK0JJYqoUgqsL7Atfv1zLfSFW+T2XbTo23fz1oENL0+
qEUdqo7ShVBzVfXEkoJBPK95wOyvvEzS8OeBhtdmjQvGa93Gtj0PkIMSJMedmy512ytf5MbIulwg
U0uxAX6R8xnDZ7oCg0gDsitePk2xB7BqNTF/MF7q5KnK7rntBcBy4Rhw1DKnP9x/FkPZBiMpDQOo
rvJJyJVjlpPQAC14OY3zEXYJ0IylcsL3WCHcSHsNNhi/JwVGZfeXLMXnFlIqumhSjKNCw4Lc+TCf
q5+YGWUqRqyBYRwUeYNIhks+hL/jzHZn1LikWPwwbX+oJWQeaisUyhd8fTDWhcjyhO1UqMBqjr1A
LuUFfKLFiu1tUaBSffDxhQ1ev+PxgH21n2+NM+/ojteO7utIDpThrtJVNd0olpCUwMdG32d3vxYp
RDyKNwg+nLGpBN0mWt+AW8+v46hczKF8rUZCBGRsACsUk1HfEGMCeL2Kl9BkN5voUjlOtupAXh4N
O/F6gbkQ+yL2vuv1txJbAnvPF4JPsvrawYg4okrHf3BrSMOGobDvv56+jYEhHVLviHvqUiSnzUX1
F2Kaqt0AmgLiUw6zQVRVTicFO7/EeiuujF+xIJCJ61iL6Tkz7vW68UxNqx+c03NmyNfZLGMl/Uzd
ng+7EVz6HGpGKwdgtv+nuPSwMxq5Ca8MqSyrSjCCo+6RKwkdmpUtPBsz8nGSP/TSrogeqEmcEV6l
QLkkosSgWpin1xyRtoaWtfdPxpgp7HidYsrpOfseGsLaCjZOJaXN/+cLL0yoRh/natnBaq6fq+rD
A1OJGQU4LF3z0SLsP7dWRYLaSb+bumpFn62ickyBWAOX5Sr66Ho75Tainnd1ayJ66LwbIpd8/kaZ
2coW1riHywiwGmIDcANlcqBjQhBpgNW3nUqd9koTdz/pV0IpvrrU5SQ8RH6aVeKY3YZzEco8w50P
L2jsrGx+1IFYjJJRd9XIU4E9ql5/7BfcfiKiOM/ne+xOYhJ3CD+m+SZvFlIWZVFMt1+WPzVJjIly
BDnOr22EpBUJ/gNlQXSqPU+K0PolJW2OVzRWaVdudgSaznUt3f3m2VkvshNEOTGd+qbOOMc6wvVZ
jk2+SWAna0CRLq+AyBcST2hE/GOfAxozr3uUUqZ3jj3+rc2whXPiVZVBevTAQlmhmx6yntEtJNtV
87qeVwShj/zSHYe6LtwYRLnonuw0aJpqGVg2WisPsJbfrjtUXxWjSJGairnoScC2Gkw0zZ+2ukkN
7Ba+k+nVzebTRDa4mM6Z5wtejqslcwpAgIEpsXu09d60qYQC9eYYBPGFdLOTCLFFgvMO+OOhG2IW
OlGR2uZGjIBSF4esmDrrVaLE5GHSVYb9MhqSVQaFbTVUtff1jRWA7DqP9ZLvDnpFs7ecauWmMrSA
0VFYzn61DDKKlKOWWJzlFEfk/gxUPCzLqY87BO3Lxf4kGKq8hZDZ1hzEq5E4RBB9sXBNo7lejvMG
34cVxEmLkA42HD7RqX/OrYNrRJV9DSVS9UGYrA17H+yU0lfsOzptAh5JhJD/4ljQw1lw7PI9ccNg
0Zf12COVjpDgTBQiWHP8O9uqX17T8ymvjF5LOEwSfvf6W5cFtSCe66S1gT8QCzxdZ1+Kz1npK/uq
V5NBCcICMiabTORZo/X5b4W0sHG56hoiYXwWtchYCRdl5H+JW0RYIKgsV0tfI/9U4wtHhTnYNZff
6TSGy47OOlLZrTOul+mL3uf7ItH/MBEv1p+C1raSyY5NIGIUXEX6zYhyP2gsSPsx08eSUnOwCiSK
/UwynEnwojrnlp35kXEuc5I++N29SWpVssU6yrxWSRji5J9xyZ7OpQPDeCaC9Xq9IZ1LE8ed/+4q
eR4Zx7jZUwhgQ/58zSn9ENYReWVQBDfjOBqYo2YPn0oewr34XQ0okrS69xd9UFd1jG4bncr1FMDT
yOppvezbtcMcw5BUNjXJUCW6hiI5+41Reib6pYcJnBZwXpQb9lYdkUSgNpZJ34HxPPH2XyhurW1S
+9548Z8R7iBEuyw4gDUuyETFm6Nfw75K0EnoAsD8pbO1qgxJPto9sFNolQM+sJXouWywyKlsngEe
Gq+NcsW3v4coPujILnNa/r+w4npIZgmUs1djrVaTyE1HCmeSq5PPuxjOWBpu30bkUlfVkRKiBG/p
PeVwhRCIYV9vLwubWnU9hcSr/krAdI22eB58fZV9v+wNrN/9X7AEL+SXzv4TaA8iPYsQB5gr/gkm
9HbKFrCdIsNVdWsxoCLsO868C7Z1bzcsuqUStNxo1wGOG91fekakF2DtO867Ksxwmd9AKmWzsYXn
BxzjAMFxSbWZiittl7uKu4dYn6o0Mg6X17yiaNpycDX79DjdvxaIgi/afFbp3vVWI5x7BEF+GlyS
rnTJSdGSoN4OyRIRFXbTf5j2JQvrpQ187ko2BX3g5alsM9SkRPR0a7fvC1UEDmB+W7Ee+G1sJI6N
9gwG65ogxO1aEL5/z915PDZwacrt2iXWj1wsNkfMMq/1B4I/KsqeaNOL9GrQe/29A99GUrqFNVMh
NmErNvIzLV/he/l+30z+UtthBlrap4vRSoV0vtvefjorfs3WL8AnYbzDqqscq2vJEFFsTJwRu9iQ
qQPQBovOkeUVp3vLlqt7vKkEf6EjCg/Lt9C4thyqDVRvfhXTcHgiRXX02mOnLBmummHFpkbSML5L
l7/KaHM5zhzFunNdG3QwP4OVZg/f0hEGrYV9dMrptd7RrajnVO/iVCd9g1dpLhLP9MX0COTnPkCX
4ymFpVkwGcFvpBh5BiPKnUEb/DgLVVIvHYgaJZjx80yuWzg2hhjEW9SYoOxTxAWMEo5edHWqkflu
T0BjScy64fUgxdxt92XGtruo7BiQCBRXqDVeCBOo6OSTVLleSvUR7x6na7M6MZYeX9Zu+HnW+z1B
5a2QFL2peoiVA4KSEcwIJjQb0eWqKB+TcfMQ5nCFcv3Hu9BcOxHkakWIM7i1mULk9nufxKCosCpz
rEi3FYpKfJLX/BDLwrhWTWI1FHgr3Modjoc4mRgk2ZIaPY3KevhhbTBkUMKETk8yfh+OaTIfDDQ2
DBOnU9MgP7KpL0xBgZhLUS6uQa55uUFco8aH8WAHh9+lyoRVIvoMHJH61qFpIVGr8rtexC9/EXVS
/BiSA5Y1p5Nf6DXl0773+63DPHm0e+9yA4NDUropw7LwMW128OuD2UL3+OSKDFGvhRSpOWDlZqZI
rR9gC+gKzuWE2NyB4FcQjaNOO1PeHL0doLb0OoGAqRzc5MpBOEnmkovdkV1XG0DXGTxQzQB8OTk+
mBptj2k0NsbHp3U+MHE5dJPP1Zspi9DDlfrxeorx5b3rpzJDt+02uDWGQNNS4E/bh66yI/TBZIGp
4+TG5k9s1xG63KCpsM9T9qJqbUMh0JtIQgNGF3tQFSLZpNSt6lqOV4niuRybcdiWC7Ay0F98/zzQ
yAW88iWXpdBJZTXbsaUL+Cptn3rjt9jYozERD7AWYN+3CiGlojfdI6QgbH6hKTZRACqcxTc7PaG8
QIrDFdNVB+f1Cye4nX91ieLcZHSZMAs78sYMHzvc6nzuERluD2XiF87I5+CzEBfGw7aeeNTewbfm
3Ppk+jq+E4xb6gzluXX5NEiH7lQ+j8a3L7eY2HL9a2i7JUuLzJQIsEH7qImztnR88FThVw4xG/7q
OcdRdchMKHQtutq46V9ZVYiINmj4URR9vp3dRU0wuF2hVk6ub2NcUq3CppTXrC7TRM+/rraMU2l9
sVEoU/1m203lrQydsds6YqqYQRTyNLtO0JwEjVhElAXjErw0M3Ag6tgKlzkI9UQLmZCSY7u5bQ6f
1wuBDFL5101v+UO8Ms1XF7tCT6CUDfB3OkejaSzTi1jdwh1gceMTb7xbnZ8iWRN+boZyZ/Cb1TH0
rKgg9kZdPYguD6oa6BxrWdErxUZPWO0PdQ/t+1lWsIyrHPhk1YsY1Uif1F2etenvaz2DYk4NK+SO
APtK4hjTGOIhTbH++pgW+roypYW7feD7hXK5K1jRMnHRQGoqJxjIHzaeElSpubcc7ozkEbKP7KJb
/zH5/AU3pMyQTEJSrTEqAgkMhc9609zgU6v78L4jRSoXbpaaDGv8FYvve6Dq/GU9e57pIsaP404f
xCgjN/nQkeQ/H/rUfrAEW2qjK/0+6XG/aBAfDoe/E7CBnPM4/5MYdyBnlXB2L5nOGtuP85dUZr87
q6fe0PCj6AZmAuFT/3ks6KrV2tKmTNBNXIKus4lsmmXTNhq16B6e25gAawP9GB0lspHGSxL8oQ7v
mi+EBNDoSS6miwoDzEOOWAoUUO7fRGmGwCUdYfXu7N7hNqY+DZP+tsRgtp26JPzxDramJ+jR2W6H
0H1Jh6kzOrH7kTIpYMA28UIjcPG25/Kg6TCwkug4hTLsk6qtrqrKYbkuoloxH6EROV30G0mmodsR
gDcmGWrCenr2wT48YHWVYXxSELC27rkFo2Y/DS/FYclYBE9xOQ1pLWurzYPFeTkwfuY+WGGiSSyv
4v7SYu1QH1yCgxHugCdcm9jgg9lqpKw762MT2jC6Sp4Tu2ayDfuBOmFYbB4kw1Rq7iBT1nYUEQvI
hQCdLi4+4wI1a1xv7qQGwqoaOiocFULwCWt+CdbsvSiIiBgN4xHewYmBy7xtUlSwSbL0bLvy+SUY
qs5pxnQtHEwLAgCPmnYMJB9g5I3d3/EK5yrKdOCF6lqgY4zT2iQVYpH7gYPvi7f2q9lXl47E494u
9/LxxeATSIF7OkWcg8jNHj1tDFeCn9u8aZavesrrFLi+e5RYaeOXYLN9HuQQ9ygOmuZOo0UxNRfs
MuFdwzjyP/eYfHEe8RG0CkIbpXxeHGdm9GGgjD2zHkTFtdCF39Uab+5S0pRTfhj9Sp92KnmLkVbT
zVwMvjnRmoLZnpXs+89QxiaRpfGar4E5qEz/RvmTrixiE/Zmi0g6PC+nv/uccqX/HnvRgOwVOV72
0sg6zSzaLSn2B0qcdKS5duEDa63qtJBGwcqKp8jH5WQuZ+D205bmicvoTJRerIJSxsEqDteX5ddl
d/5ERCd3H1lOVsYs1w79scMIv+UBEQbIBUcRsmeYlykde2y8IX/SlPk2JdKlLU9fmW0ss/cA22Dw
8l0CcLmHGjNbSXdobV3iXT5nXcJqjsyiafoLjCwo4SvtS8/v62wo5/f59GTVVHdv5iL7QYjl/DTb
57BsdEMIRfu9IYJKLKxh8TJeEW9rT7hXBzvBteSXV68EGxFQjrl2plcVjURjKop1alZEClbWeI9H
0fA3UsAN4n9dX6Fq3mg8Z4IFdc1+7iVhgmfLMlgLxD+Ahn1WkIzQY6nEYC0xs6oFhwWwjd/bPYes
LvK1CYeS/pUPdsH9jznYg5F4wEKIInoBWIBkz4JoicTyyAzZNlWosz4FZRaj52m7CIpX8hkegwHC
b6FMM7aqA8omZaFu8KFKtUsBhj/w0GlNOsJGswvsrwrV+qW2+GNKEhhCT6MOCaWBFiHyAH+ostUr
cVTCOQFOLX29KGjSDZhOu1XWyabY/HM3bx28yu9lNww0fFAywNnqEdl5NPIaAPAr+mlnX4hPRoyI
OXjdE9bvfvn+mVghqbtTTzl8h3E1LwnKNqz+YkaeIqcSAWqifvX3P4oXOdLg20ykD+joRmSefrXf
B9ApwrPxjx1hKsr/UZLRe2EAEcVBwG5nmyniNMLKr7/EHC9LEkObxm1qw7u+KVVTGkqmu2G8TBqy
p5KW8stz4rMK1CVgKmsHbAkvaVdDYsqIIJdCV+apvfrzGuG6Ysz4PgetQfIHej01MoUzifpZG688
P+9H/rDXGYLWzYQp495pO4Tj9SoCEe4KmSyihwzu29fnbhYNNnWxPaRp0/wZMvbdgME0P63kfbGD
V1PR+TCr0EvJCG6L/sRC/EJpbLhK6k6KcQXd9pbj8l40hOtZckgYm9dH5wtF355gNQwCiU1b1EMM
xzlUzMtaPa6P/FtqNfRby5zZ80SrEwx4303/yszzdbNSsSCZPpVv1NR53atkm35sKCvqh1DHvkyT
x/eslnT2jKXywt3V7T5R8S3/tJ4QoJuGrMBKEQvSWlvQtq7E1lB/oJ2MijrdUGlr/07YpBi2++HD
tSWaf4f3K86pt3TeFI0djDz31ySLSBDfhLstfjoXtuYYAL/p2crbHwT+KBoJdBliti/IylPlpJNk
aAdK2wFYh0+Z2GODDjAi4auwYMO9uvqb2Ybc5SrLOzz5yz5vK0c5GD0rh2URCetCOC6K+Iy5dMgV
1hfy50rlJIi8L+sWu6K8du6q7DFfuIRd8RKyysSk2jEi684CWoAmOkuDEdEMOsvSsdXNrKERRZZP
cNtpEWG5pk24YZm63VaCrApOr7XUT3iG7s8u+gifgm5U43hAJT1tRigfLV85octsxtD2g+zn9B3N
DzfOBq+tPleskz4w3nnxzKYlvkEw6Tca8J7KLA5h3QDY/UUDh51uLHY4DB4VuNYP78u7ALamcfYz
s5z+uKu9eYd4IkT3xFxYeAiG2lHRxqBlgf7s5uynVwrOUl1MAprXwTxbgpeYCVEVTr3MCR7CW+Le
J6To70fAeMA7/3mZcRzkv1xBzbYxCbQik1Q6Du20qVqYg0zC0SdozunQaiiG2FP9DdzhLqneMcx9
21no/Zm4gREZ1VOKNfkShVcooUfpLKxoR8wne0FYsTw7A6P7DpaOxHPh3p8VXbDqM76S3/1XDeGj
gzmHA/ATagAeGlyYqvsm+bt4LsxKE6EhvsDC+ebJwgGpkRcRC+S479sxmHLl9PCPHrn8Um8VUe01
nEzj9Z+S2yJ3hd4BbmrUot5mqwekYrWCXLKLf1YdJhptyXN0Js0kuwbZqgym3EPhCBSH7XsjYd6x
3EexP71wHFfXi4qVFBYPaM+kUh1z4BUgqH8ho19I7TbBOLvWwXvg9dvzykiq/YxCjS8e0nRpMNy6
PAALjQztNrgKvS3Vcg+hnAFq8QFRIcVgQxX4UxbjBnfuI85N3Pozh9Cpm7sYXGX6Pem3W9GwxrTo
Lf8854ctEFySTxr9bhk9daPAkMqetyEPNCjPF6F63HJ0uq3PBNLJhzZ1p3d1MKox2gn+eZ0ScPbt
jcpu/xJf089dBUxmQbQN3416aOUQdrCyMehoPp8RXmTdklXWOGVJ+1TGtcD0bQERXBfPXakDzRo4
PRs+LoP4eV3CqMENtww3Bcm7estASHMJJIsNDy2YPqanvt7HQmtIH75P/JHlg8HJdbz2Idtt/zB0
p5eYvxIYXV9EVcko/f2xCce4HXAP/lhRNh4GOKzdXkPliO7jZBmAj3eJpgtHbVgVdd7Hh+AHQ29r
kOCHB9mVryp1WmUOsyKeSM7jjYqr8L+39HrOMDbW4u37r/Vr+WiKTzZJQasHZa0/EVtT9c1G265l
w6/1eevyeQB62bSUokXpamhA/v0M632lkJ+B49k0g60l6G3/lkJ4nDkCkzctlpeJuRQ63AqW6PST
kmSYmMzIpOYzhbSTzUL0bnqVXPn9nyVYLqAtaW5OaVkSEzwaO8M1Rh4O6NgXK2Y9GVmwsUC8xvss
kbSXW7FaLND0Q3aY9F0r4VdS5w+2loA5inHfmxfmeOdsA2sHOBdUmQEiBd871G9oQvwdXYAFBpJo
fvkhvB1uPHuOG1dTyrzADPLPo2tyrvyHP6IS1MEt4MDyWzSIslat9BDFnsIb8RmngKN6nLNssZCx
izVbc6S7Kjv8KhbXE2FvrUme67FCJ5Jv56sJshr9oCJ6vyWbDe+9sEcOr+uh3zrNposVBNXtsqhB
/duxEEthnhzDlzdnDU1TEJV0+ufnetHc2VCTekHIXUWR3bePnN6JbMU5s/xQgWTPfYhx9SDOpEZa
QwWUaHE7uTBmDaocLhE1rlkGIV1I8locMgaZji9i4NdiNvxSsyKvjB17aCrpbESKdZ3QS3OkdWV6
cM7pNH8cbAlhgsaMz6dTV7tlsSDlusuJam0HckuPuUnoHPrsqOLmBK2DtLu8fnGYxac10F0JKeZl
g+Ji8Pn79EKwE9760XUqGtRcZP1EeiL/n2mygOmr1YLjazXGjWH/9KDs533sByDHsT8cWS4U3Nf3
wypEWhCmYIu7A0qp5yvTy0m4zbj9R19e0NNwm3n0InXIJxoqpYrbBaSKkil2lqbU3Kh+uOQscoNf
8FOE8FwdiCUQ8HIuT+xh1MZ9tVqiKmXX6U0j2QZEde8MrJlhlAPV7mqIxG4D5KLoBSWlJGOYVpFW
qxgM9AUvJPtEUdJWYmrthC70oI9vyxecTrt1NOf9guOfxAgIajxpQjg3fPtjRPmdo1he3smAGwSD
sR7ibWU/y/0O/8Vs6CL2ITlTCBWmJ+BbfwMp7DYr9upwzyimmnTqP3Nfh4pShzVtSmX0EUz/lRj1
FM9pIILPLa3iwbOHpjQHddpJc9bismpKUJ69qJia0NSJCzFwtBwggce0t1K5G+CuHqu/2lHP0cJX
JZ0am1opuWJ5ILNAkh8LyTDeMZ4YgwnPzQqxteiDTqYq7rdmUf7ujyMZuBCd8jP/z72ZIPiRlYc6
lXUBM/+elB7SGolFI4PGzzvqFArDtQdbjgvES8Jyk/qJ5YXBc1QJdmqqCXIwS3Sd/rtodFafHqP/
KDuD0RE99m/0BpaQE5yCvcwIeK/jOpM6rEU6anJlXg5kGFMa/VUokRHvAE1yDnaUx7kUrPk4b4ku
GhwEQasy+u//8y+3M29tj2q8ttw252WYd/7du4p5wFI4G6BsORmnNrkV0bWoMyJkrDLzGX1WMbn2
VoR0fTSPSVhk+fn4d7l7xfyIxwCccoGQdND1rRutCdBrma+iyAq4UJMryjfVYePC9C6q0PWzSwXf
FLcVepvPP8dVAGzoihB857fQCMoSNxBOniEPk5s/xn/fGMsBYMje76VNH3RI6zDbxVQbIwnv2uJZ
qDu8Z0QcK9sQ0Tk/xFHmDM9tB4HMsBjxQnvAq1QFE6qY5kgvW8DrN9kkrGaQj5eBHhk0QiCOHv20
2LsCCn+oU2eS5KrUeYk5oNhJ8/+32667hkY34+Ht+PSegUyNZWbVWF+i1P5TfHqjU4LVPOEv2KTm
G+/AODqWcPBhESORhYGbwWyqqE+szGUIEogffnuEY+i925NgsREgDLl7t6lO6My87azuRWpo2jpY
R+LAcMrwZvjw2gQwNRHMfyZV2uocxcz6Yw8rEAveJ3VvA2x/tpFtzMeQTKjTvKFL+ZkQjO8CCXhx
/9m5BtuZFidwNgDJXZcQJ0FZOkQwmlvhSvmbJcDpuE4RErb/+arVDU0WnTzyC/CsZ91CVdf6vpHM
7sZI8w8j5SAtkuQyXVLc55JI7dja4swIdW/yqhqlAKNYaxJzdu7ptvcoQaZrYjtHfWZP4PrK32dV
dnek9wEb5FS9CFAnYMqJ68ok3oAZ6Wxr3uT0rJ6VeVV1hO6xLkrMiB1kwLHUyXyMY9aANFQoZN92
GyydBGSaM7SRA2OU0tABRTZ8DMUGUdqpbU6R1iPnZ5I95nbLUxXRje4gk38BFob5O6J55X2qxjp4
fGY4b0ylkFG2cbMew/lM9lGzzd6T/OvKZYZ23Vqg3lTsSkDrkBCXnU9MFfDrUAsxmPB93UesO+q6
X2+k4GAAPkX+4QDqLzfWcImNNFJeCeclyfAnRpBNx+wL3OXakeOraCEokLSy0HjU1VU+jzeDtygI
7btGkko4NG8N3dtIfFwrTZnhGVDjZwvTkS4LCd8fHbix4Ejm/bgINI+F5awcOQEsW4zN2GL2Lz4v
pebZByXD/wiXtfjnK4IToI/BKPz9Q0GNOafhmg4btNzzmrQ8IgLKKYk2cnajClTzRQntiMgarJNg
erY4WdVdTSrBMyJVetGcyG5OcW4gq6cUoLBBTE7QrT2dETaR/yHm0zOFAJSwid7CvGEwQboMGUJb
zR9+rFfFZmdg8sFpAl4zxfpzJ9SGXQoT3tkkxtqmsD8yPPGqVRFoFbkhpNvjSR0ygIJU0NyOwyCK
JnYM0wI1IOegz0c+030QiUWAFStCIUVz2pr2QK/BvSRLPe2JklZDw8Ol7lW/MYYamjeVoiW9Bl/7
WDcs5dlbiILuys3XSQI8RhH1wCm5WeLH5fh7C2g/kanudqbx1ZA6BfUqKzLxkwfcvgskUhMO1BFh
H3LWIaU62kuhTCsG6/eYSM0zuxHZDneVuK74nKS36HwUnqgy+c4RmEw1U9UG7eFrUhZtKs16abkk
xsoWiDVUJEiCfvUADgD/huOntRBZ7vvq5P5/f0ToMtThAx/EInKGz+1cLwKR6U0icjWqKlk3e1OD
77OTM/OTLxWEtuxqPydfUioExsWf93NDZ1k6lhEV3g3nwaqDnHiVyyRpAM6plbTO3PInV39gTCVQ
D+KDCADp6xx+loj9mGbcv9fWgzvGu8RLnrv5CgrQF3TXnJ4i9p72KTu6NNsoFs1zKnhEzaF3IFn2
om1INW3l4+8J2H0/Zn2LCw1LRWwP0VAVxSk5g22UZroFlAEnH5eQRo0+rteyOaftKs3vCDta8p/J
AX+7qB05mtJy7o7eBlo27Vg+4jxkAjTOPWSSIbFRjG+8ne0eTuwmsnI37LpzWNg2H9ixosIc91M0
GSZXD6i5EGDkiohGQJWMcatPG0Sh/E0CrfzjcI6ZsUHC4OUKVOu8ydthlX9V0+WMbp5ndw+363wU
N9RPJEbg+oa3y/Rg13TGFQ0AMGV2ADxq1PXB8Fkh3uaxGCzG18d5tYeIvv962k9jjawJ+ABZlaWV
xWovxuL4s901PibMFRxeDstDtzMVZop0Z54GJPe7XNwck7oDEaCkiy2HNCvXVq5P9ZpjP1qCcCgW
Qicg4uNiOEzydgUVUsNKRhlAGJpQmz2TFM7ejN+r0XPvVVeyieH9kxtmnuGH+QyMRv/8FI61mjYz
EQ30d5vKjvlMo4WugQwqhb/CLrTmpUR0Se8NwY1MFcYpUJy/0NP1Hgnw3cm736SmzII116r5qUYs
GYJCNYfvMLwrCer9NZXpp4HhmXjOPpX4bUUQ1SRgP3ocSlC5l/8QwwkUZbAjM5PfXGh3QHR6+e5L
vQ21TXIERPGaCIP//31jbl6eSv8FKbYwfU5ztplczn2jHZESEJMa9eUXqxOX4MUB7sQSpVixhiCI
+GgmfLmVvdlDLL5129FXOVkrfXk6DR0W6Hr1NlZ+JMdY3E6F1Kcp5XTkewo3x2BYw+qMzeV7h+wx
O3ChBEflne7xgTyDPUhCaYTaelpFePrY9n8mHpQKSjSqkKzJy3FqK7SRajIB0mJh2DF2r5ruXdoh
Bni2YC3CPdCkpbQbCVUZPeEV9QbQiDnIXU6MoZXWHW9YAnnFPzYOi9FDHS5TF//Qv0zjwxLd0ODB
YGSTQrycautpIVgSk9flS6iBm6DoLH5FnxiyfuhrTeAVtPKj92MjfSRqlyCcJ9ho9MC2gq2xYU3c
3GF7v437qSZc9plDfKxdaVpaXCE3CIiOVeul/+/LFZfmTYv5ZuJPVspA/vpOW1d+jQoOwjW1nnMU
rbPL39Bb/lZTgqPAlCxlGh7WD36AeqQ56fD/DS5/Rw6i8Jk2aQcCqG2POQhzqB/BvB7Fhh+xyxPQ
KaDTg2JC8GUVEDamFGE7TN2diLjxS/Ko0OYPWYGGPAoebi6WXoq+Z3mdHWG1jzBg0ryCxXV78xGM
KBTPz1Gecgqm13wBwnxoLv0p+n12kv/fD3JV6Ob4YjmgeoYIeeYbvO7f0axhOXYEwLbMQKbjhJaa
heQj2HnwMZUoGsraH4pp6UzIp2eWcYhiQRsE7nCylHwbOEVQsoVN+zk4inLGse7bI0WjRFFMoTP3
8/IjknUdrXF9zRdd/w+QP3Y8CGtwjxI1bQdNrNa7NH45NSMrTSiKLI1DmFU5kjWEPZ0liUobEhkR
vey3y2htJG3sf8Vq2N+Sw7IpcbldQEjppATJwu8qC8DMOVNSNqSHHfoQekYFPfRz+kTI2Z9jS0PG
ukTmMSV71YM91Ev1zmNJZ00qxbFW06tNuKjh51eU4edj8qj1YxSlBXlAPJG2mCo9ac17278apDSn
wh2UZyfbH3r1PQA4mmVdYhc+P7bwd0pOfj/owTiA/RCyDNIcAAc1cYifvt8DkxUXY+aeE/jyiu+r
a7p9ox0aHz2cnhadG9gFrGJBJzoqeWDgzhgJMx/QMCI9jqbM6cC91RUhMxgiiToK7/iftWXkI85W
GfOYKttOyoas3V4LWvwZfnPFzk6iq08uJPOp1FulRDRzz0H72YoJXNKNDvlu8BREu2eL3Q0aFGi7
ibyPue2yf9hmvCu167qWqCoKyZarZRn4+87mpm56smBoVKr7HWr5CaR+OSo6Nse5aEzY0lTcEFIu
nirXut0J2Sa4r3JolCKwk8OKVb8JiThIZSiYJXR5HMaLlPIYOhdTwdfATsiiMBjP3tfvpKMhPb4u
IscMgvBWeLB/ofc7+OJVcnpGdgAgiWeN2ycsWOrYChayrJlRdqs6bltYs4uCMKxqORKvPjpCk35V
8IYstF+eEpolzrmP8jd7Qjkvsc2GcT2cUJH2yORcz3gwx8y++1w8TLofwGR8YSSzjlMIXzwNwtnh
5iO4JrxcxqV2LPMPC6Z8mWyXsHzZqqafA5aFuYP6HhHIIhjHUMGXpB7FUiCkzRt6UwJFnV8fhHsm
QA1ZGHMsI/VqoNgOBGJ96jmzlnDMKfvsveuRwaoDo5+/XoTsKHbstYFB4nTgRA4xEUsotlGKou6J
7o3PTGTQEynwYyVujB5wiXKgmmUrXqZyZ0b0SsLoSWTCxqaWFeOmsD3ptCe/MGszg7OLnR/kh3J0
bWD0OCzvUSNFIxH6D80gq2egaISGvwzmPCxu618M98Pt6bh1vuvvKbosNanBOVLsteLc6GQf1sh2
G0rFpDs7r3aL52ahlEWo0QE5FPcHhOLndLiSlTFCvelLTWYxSONiZ2C2gjsRumAsLIv5YCTk1TrY
axWM/qhJU2smBLaCPfcQ340f7cQuMOhjmRgeKPixaUXlXtzkjjxwQPAAEQn+qdhA12CJrbOPVozP
enVqjUEMfWEWlXVSbzKdGTNb3zq6wW64mdQHbNDCXMMjS0ug7T4eByZeasdeHn1D2flsLr++V6u2
P3m+52adwzTWpfwaGGNl/Chpis0UOKBT5fT35aK9hOJ6gwTfP7/gOszAUyceVjfbUKF1uZNYwIin
VeokmrHVF+/gDrMYec6GqNQaxOLsZ7fk3dXp1rJ2JmPinutONuY2OKSAyQ8NQhVgF9OCFqr1+awf
ITcTX/7tOrzulO1Urb0D9nj9QpUNy/1Je5TqIK+6DaQLaRHnqtq62Av6etI1f9R1IcFBXmTWkD+D
B4aJg0kHNgZFDrJyeZQxCoAnDu9AaPduYvh39/kS69aYQTIbB2iYpN8G8UMoYVi9DjDpX25hVQ4M
z/n/6b57u+OsSzm++Edt/RRcmfbYCkpUH6+3k+zrRND7qwPhCXDh6YTVvHSbm25lDxT1UBf332Af
8rYHnDjwmz75g+zVGRc5Q5YzGaiAG+MwQblB4lSt+moQ75ijptTZxuSe2vMIdxnE8JoUI1FR5Mzk
NmfDDRuQpNLpvokqLtctqUuXKhKrlJwqYJY64O1grbYE1CdVgcTJ5mg8TgD+p00RizNP5BlBezvl
zET0jI26JdyevI1Vc1Hp6Wwoix+t6tik4OSUt9LiiI+SJhfl5g7R8ZnuRuaNEdwx9I0OlAzRlwRN
PifGJpxBihSu9hGjt/91Wr3+kNYLhgDL8XzZ9pzPoRKHEPvND3jOfhM93ewC2UBkaFN6/nHyFR1z
eGJMjj7N2ILOViPnDFZM5ETkqA0hyXZW1o/DN9my4F3qbPqCBUAAnXIM3505camrfcAZMp+AP7lF
A/IGb55raGJSn+sPayC2Rh17bdaId/WmCXVlJS/DP0vwh/rdKe2bSylvKNiZM43Z5+k2XjgBPjTc
GdHy24N3qCAbHYqQpQwvgaUWxOBPZlQoSgzc3GrkUGKSjW7U6E47QRvPil0dGn4PVuB4dhFgE2ua
cW77UYtRdAPdOMBW8qERIjtgjGQq/ShSTaQYITZfMnFFV3HzFacHIY3xUbwxQhT2yf7cyczyv86N
TsdeqduqoBzIDPniLdZcjEP45qUEVwNRYTNcVgfeeg3I10+3EcJ2lDRamGRY+qXAcjd1jqjClkYb
6eOP35dQV3F+CqjRsr3W4lZ5KgZYBT+lOXCHYujCUPzyjOkfdjMWRjvGXkk6EYpOwzFpsh5xhpct
KwP7z86Nlq4IQoXCbIBOPVVYuGxQUjtzXWQKwIFHSK9NB14xbxyXlFuL/sdok/1274CQdwlMhurO
G/esZ6ihnHMP9L1ywwphi9+53b89Yj6ZdK2pfWwKiweKemsFdgxQ2VGOqw286Gus3i6OdAWy3bhx
ntZthoFWZHf7xuu0/Oa9oeBoKckFVkXb4+9W758jJz17oUTagfdgEr5xhbVW+fcGJuqoHaQ+q6dq
x2Yi3dDU4jHXmjvuezMVJ3unZbrkXI8hzkPqWx7U//uaOPmWh9sXHB35oEtO4Mfa4IuqVFEd26Fr
rUbPCg6fCk4QV13L7LGGvUzuZ892+bDZOMCuIHt5lWHuMAyZJ2l4hroyHGy53rpM5sffS/AYHWx3
K55jZ7iMJYsDZus8/dWJkf/kL/YXEH4Ax742q7zE50+4oHcvMhyRFkFTj3TY14druzcBWrA1G1wl
Z/VfOmTYIST7rY7ZzeXoNHYp7owlo5XZ8pt0YJQO2f4FOWC9JOL2Q7Wqm8I/XFhcfxqfvHnMjkIu
MqoNanlFgA9LYC+YJyh9x743Uu/M9KEr/bkDC1K6HwMQo6dq5IKhGybwyxcLseaI7YvkmHrw+FR9
f2jchvkH/K0wkxZRA17lfETAhq3xZeiAqe79ZRUHRCdFXULE6ITY0lpf4eKRdECalgEpHbEqBpHP
mXq0xccZjNMB195zSAiJqCvthTx/JXOmJCIw+w4cMQxPFwiWuFo4ZX2QZfClNPRklcYqyqbDVdjQ
xuQazbEYPUc4DEzf2vmhqTYs7Rl45+UIjHEl7qkZwchXhv66MDret266cea8tKU3taEMV994wcwS
oA8YfiKS1MRISUEtAtEbVsdvS3Ib2fbViIP0R8CKB8Ws7D0J2TR+5pKXM8AI9rCZI8q6CgVWF+aD
l5kVXhqhJrTWIeenaOXKaihvjeoBvcsS68c5Yu4IaibDjvwORFMoyyiFx9H6HCI/2rZOjEK+d42O
SG7L3CcgfgHkZoQZnVeWiY2sbK2EHOFVrFnIAsvixl5ulzTNoALJSlQZ48j0aVdfscZtA2ZaEHKD
VMW64Z2NyGYjKtU7ElFaM1Za5X8dJFPB2FkEjoD9CVe9Fm7MhkAdF6As6ssHdQkzVeuhFMKj4Xss
opJ1Wa0A3GUqzqAzpIc1Q7DwFumUopSRH9zHVyGH/NqhPgwxPZqHZHIN6P6Vnu7Y8XourWA3xY/s
3MxY/NNBAiNt9PLAGgo5TXQhk9EPJnwU0/lyreL0xj8TN9qdZjLRnxFLsj8DQo50fjf2fjxZG2Dl
0wF/SY/d+a+x638+3Yc1S8v1RXEWrKVCOG56Jt3CPl9DoGj2qcv1Y99UIGi29mtkJ7qtJVtseHVi
XIYK/Fe02XIykWBDHsruPdMkXwltWwFj1KFz9fXwJWR0MCvmEwhvYswyPGWWZmyb2S4dXeAu+suX
VSgfAZo/ecdybkHPUZ/Y1wmoF6p5dRxBrMsLXEHfEOJSpu0THb4ySXcVQDr97zBuD8LmvmddjYJs
OJquYIkd6iUmkDElACD8QFzyOZiu1UWJSg5bwIxjvgnhAWwYOrq75jlwFekEUAIJmBzhz6Qzrcdg
ovJDRPMZAMSR1Sk2lxJoYU43SIostT7o2qcila6+qqITIsKVzFx5LqHoWyFbxnyA7ltkH+8xngL1
WVbRENdHtDylhP2iLTgS/8jLk/EaRbNgyFSzf12zcNzWpls7bUMtQMrmphwvVf2QO5hmFviKMfRV
UCFo78ME1fGS4KrOVsWqu6iDmrcg3zNmXOMGtmGnwaC7OJD1++sVbe6zXnZ+7OUgH93GEZAhEla0
ve6L1cu60vAcxRfcGQgyUG8rJdAmiWSi7NSs7FlLrJ7FZY+bXyK16Ghs9fEFop24Vu1NwN8WsWEb
JAwECn0ETwzM7slpiAjkyxLBcSbC11JdGRXTIw4xOxcWTYAT1L38ZzriHbEUTsIoOSb/am15FNR9
QEsUrF/lbeD56D6Z65QGAjdDWrTHM22mDY3SKYuWb+coymB63RtOmMzM8Zu/f+uynEb4CRHvA/iE
obO0KTGOtL7pd1yHwGTChYTbfL1v7OHeJ0wFhahOWbhrM6YhyIJvVcvfvvsQ6c7rcfCSTZOuSvD7
vJEdSkaRBLB1YlQOxqrXKhpOfzgEUUViCyiYaX8VR5EPRCAnfADqMuWmZMxj+YFdIqr3eWgxWOr/
f702ga9ZKmVoepNagThDkoI4tiirXYOI9a4tIz6W4/hvXWUmGK6Szo6OaDFsTNOOXYX9ETwCL4kJ
HyIxw0d/VDRwvcIbo0nwVR0rrox7nL1WPdyiDmvn+P7L/tyVjU9pugJvgWz3Z+Af4wSI6YU+hYtp
NGwboirUwHHjs+9en9oPX0KFsQBe3mzBzBKvaSvF9adIaJAOlkYgY+GIzLFkJh7AAtHOKCuLU1Uz
XignZaoqxy2BKc56BhBR/jJOpwxLb0RldKLkqhQEZ0DHLcfi3CLlhUpfvP5zs38Lu7IunRWxhaJx
GkGfNsvnUkB8p88cZ070NpQWKaku2HGeytjw0TATpF12cb7yFUisvxRG4nvyTsFZfaLnHM05RT/o
akYb+Xz0flQM3J0o+HI4ktoMVUyPBz4Q4wgwO/osQb/srHQYZ+il4na7FEquwldYzA+s7QTJ9BnC
Cn6764bZ9zFv9VoQI8iPxY+OstuX1VPRQOqHK9jsfYdXhe3IiAGkkpB5x1NkMgAZHna1kDY1hRz8
QqgTJlFxYkk6hi02vzaOWepcFKpCbuBcxlaL0GVNzpDtZbrWcDXIbhTBwaEw9fH9/ubdFQU4/OMG
oMHG4BiQSVwE0jLf6nkg65CF0TucBJ2TxlZdIDApABVXMJDWH5lwDQE2Jgy1uaLqulaD5xjW3BvU
HkgzylvoFXy6W32y1DLQ3H0gHc43qvc8gF8oG0ALvafzgLhnwhayHcp0vltiLC9Fo2Mkv00WoDAL
gFX1vKFH8jHptyZPMBS9hjE1P11wJ64f0+spI67/77MxsHv2H699KW3E8HnRiEwGtEJibX2h0ENw
pSGi9DJ3gMUkolijfOgoBqI5oGeZ8jMg4qsR3oEdODi97FIUxjArRW9UkSCkPAOIdiWFVwdPEU2J
wSPASv9nReMm5OLgRF1AAV7SYHZ9Bijar6prxduHR8EuLxh58LsvW/Pmh9BoEFwiI/GT5tC0VfEp
upSEgfKm0koRB4GsngHkFGMSdhSnlzQBzjTEXBixLOMo6iS84C4oJKOdSPpHlDddNsjwEAkMvChP
LLOd7SXJCuz+VZBkYjlMrgm2Eg/rqLw7+RN9GuiigaDDsS/mnmOiNzbVfmCl2oj94gBWTJ3y+KOP
EQoB5HYwp9Ye7CorLcRs/4V0jP1JNa1w0WlTK2frU64YEd4aXpRKiyEukdS6Vu4KjyoR9awPd24Q
ckztdUBVm3zoj9MoYupFltCiqC9KPkijdF977fC0y6B/NVI96taJqmpUHil8kDi53W7JOtCFGsky
EXBrWr2LBq3eLJTD2IiCkWzY9+Tw46vVpY/OIS+vzsl/xCjZDOIe95cQZbIuVj+e5Wq2szEBzIdR
dq/Oh0uuZrxaWSh+pDGGqcpIn5f4VbuFWEtiImF0ZLimSI5XnMJcgjLGLd5tlUylwmivp2KrdDPK
g08grxnCJcUzbtLz0FVgjJWvB4EvRz7uS9b7Uu8tF8isHA0TlgDBzMbUAbCM8QAHy/9G/e89Ombm
NpJJcew3JhlJgXUDm9S3ubHMXt0Vao5AIdTzclsGyr0aii0W28gUEH+PoD+8IQh0LjJwj9aKqpc4
gfLsK2qqecyO6CK5TZMxm0q4l271a64GpRuntbUBJ57dyTPQohUXR91kM+Ycy+5GCy1euPCnGFhN
PYIztg8CHhRXv3LCwbXYNGbKBIw1zcvn9e9XGJMHdEu50RihfwRSznBgKeyyu+75ssmvi2EZcQKa
PraFAMvBAn7rfJeWuk27wiTPpxm+Bh9nGIcgyt0iG9UOds58t7X9c2mKAybeJL06z4Mi9O1b+0Nj
hTXbHdmFL9sGq5r8v7eGqk+Fj3k+FK2LYxurdKX6zRBH1I4imjxLSYFX+PPaphrdSgIHucaqgvEP
hsxiKeYy45KCVaanuDD/0umOe9UATA7xfp2ItJ9AuVFc4HI3FHJSmvYyU5GOMvur9R7TFErKUdLR
E3fSDL27xsuAKD5wWIhzeZxEIvbOAMk+gHBeyVMaWnCJhDR5xWrfhxj6n86tOuEFf+3oNJct/DEU
8zb5m9BpwBLmcfpcomiA6TYEa4pPDV8ZYFLg5HeUEB356Vw2yfBeSjdIX8PK/fgzvIZ737HBbvK5
GXbYQUI+6NLlr6tNvV0nApypdZsrTBnmySnIbdi5f2qHfPaSyt5WxIowOJ3iIW/vMEa8O9Oxre6g
GEQUZgt37CoVa2nuUaN4IPs0XFkxAi/WmepdGDfq+BfHfBoZ0uaGL6gPnGKNyj0IR9vl8yx5PbXS
1NRtBhI3jNlTq2LJgpUeZU1xZSfRLY1td73vkiicpDhXqHolSrbYLpJfdLdBH2nQ2XWpfGdlIa4s
jlfRvc729DgQsPsfjtD6FXoGC35mATYMqctQJexb6wAX56Z0gPkahuw3WCpElHJtvfixY9iHA16r
jGF21+X2LpIZqqVhO2Wmx1kK90QgYx9vnN8V4C8b4C5ye9fcQFm8rkRdGwEX9Kr5uYW54RN3Y5Gr
aLhKAsmXsnfpwhlMFmAE0GKrKZX3whh43DB3HWq1KozvAcx/kighgNC0Ia3zaXME8xb+pxGFaIfs
Uh2gyfIP8cSyk8+aasO/mptmPFm83VzBnsKsOdbjdau69eoEm71BCalNEuNnNGJt8lLdvhcQd5Jv
Qvb61Zyvmf+bL0AtOhFw9syxBVno6tXpBjOjS60XOdWNpsWieyzs9x5R6ZZFbPe95zkztRxzsWiU
nOEScuX3068pYNKuJu2v+EkZOnPyYMV2FVU4jOeaTLzWvVIaEXdVg4q3dCdps1NEXdSx4lDNXled
nILeVMfdljhXbKR9P2hti1Ua/7aP6i8RnYkG17zf+pfc0Bmq+oyMPlmhCDT/QnVDpr23H8oE3UXX
Z+oUthZW3TgGRux5FjYjI57YIt9GuGHwHwuC1kfFo5hD+k3crQ71wVxfoVxFoc9rhfWHIDO/Co34
JoIMwnKEDUr97duwiy3t2eqF0XEWjeqZ3pq9N+1LudhFxBp8idPhYzWVHEXqkQO6A7TGQ7n23hIl
8XG5R08leKEeJf/8tx21wqTLPAI+fykxBE8io8SUbRuGMIeGsaxtbMcYdhzt2H1sgyxuJZq1pydj
SaNIluu0XQDLpMXHQ5CntTwsKJi7y5xML7y4m9fsg1MGhNc/ItrdsWt919O98k9JEYHovABKwl0l
V0WnC0hR+Rhon0gPBcnqr2VFw42IdpI+MSTR+fSFrG2lUx1O/Hh8WAv17oO8Q7fL92m/AdaPXkLB
7BBvvu2CYDFAmjh+Vxv+Vi2wmO4fD+9KaHEBaF3Iy1D7dI0h6J3qL1o9Quw5lSeWawKKy2rToULu
yH/qErMinaYbkmr86oQiDwWX9srStUDxJ/B43GdZd+M9fKAHFu1LWhDImJZsGG20ntiCIb71Wxo1
PiOvBarb6ZNIFGKGy9FnMTDiPDgJgDLchHHgY6kY1O40yRUNmToG3ZZAv7LJ6qyQ+3BP8fyEeCZI
lTEVzu4P5/DKQpN2ymUgKgd9UZKyN9h7jq6sNbVnFbGT3kOop/avA7xcfaXR2+mG8LdrRDuwoaA1
Se260z8ndwr5MMrOHxa0SAg+kVVSMOu74Na+/u+mR9ig3YyZJNUSkeswSO745eg3ymJSgXLGT0D+
3JHMvzhAiQHTUi64lfdzqMzrQLr6zdXwW3Z9CyjpKpQfkgSIakK3DVQ+C2wtrblSo+XgarDguUQ+
/B1twNl3URUdlWqmscKSeHWDJ59jaTZoFyD/3PX9l3CDvgcR1ctNAwK24rsOVIh14N2iLb/LDQEQ
MLZr01D9P/FZzTs9NNEwEeMZZdjZca/FtmmzWigUBclvb3tLFLBSuFqGpu9qu6ZIuZLE7XCH6sOk
2ZtYAbbcJ4s52TbXwRoZ4DB076aoVgMh4i4u8Htf9VMKa/5rvNwAE+p/KK1UqETPlXEYjxjNj2cq
UPNdhk0nnVxXWKyH7D8orT9W/4TXEaUS7CHxq+1o8GOiQxoMq95Va69n7csg8F2MjK6tyGPahK0z
Xjzf+1wb4pvXoFQp6Whkxg9zsmu1SGwZl7rHzHKJtx0GdvttAFuypRJd1WcFo2aTmZsF7DX2Qfow
qGgjJchGexO4BzSppGV/oCAdcMJNcdQs15dsr4Z4QXwKn8ePyTd6LaikJg2s0VJhAfMssHukusei
adeLdW+e3idEHm2VfGOklxn6XMk9b15qNf70e3Wlc6pd2fuDjHwYmzfngmCKMsc3IL+la73ulaKk
y4bVwITkZds9QfG7bMkbelZjhZnSxNpxMjSmJ5v7I8Dy4jnXf/Cn6csV2CRgp3quZiCxiaWwTclK
jXqImEDol+F1WYs2qdt1GKTWAc5yQQo4wXtI+pSBMzoNzFw1dZ1CGmn1n8aW3fRBWhk59tLLoNyv
5nLtLM62NPfvZMh78/PUrDZE9LffxRLyTSV7qSwbO2f3WtpkA6T3F3fIxWhaMOcqFHRCggbxDqU6
N42oj9FS76g41wn8o5AY/aKXLZo1IUd66T0AHZZc3wtKGjKRGPeopozxHXvPYJcv4g5xz3BuTb9B
NlGZy/lhmfe34jCL+ZoRu2ln8g4XJXbK0YJUZr2mqORU0q0pzGOEcPovWQVwaBZV1Z+xXpswbGpX
Nc/5YyFlU1XhosGeOT3PlffwXuJRFhz+WDYKWegIV60a2cQpHZE2otHHmPQo/7929r+l2otntrEZ
esk8FYxmetMJQM299KyjpvoLWDcHbE9dNlBBsk4V6OrMuMwQwVBB859TDVWehmUZVYJiMmDO2eqP
aVFhFRnlcd3Y6FXylZK2JAKaskWucXNCeDfiB5OSXu1VtzD6B+3fTlEPzWJfl7At5Yehfn4mRIYb
a+0lFKmRuLu5D707WZEOhmku6wo0MOrOgfiRjHec8oiIBaA0TzaKmwFGGJ8yIqQJPH6jdE7pgaN2
twGjHbWzSrp0HzA+1CDoNWrPtXOcn/ERu855LX2q9+HNBNHKG89ObVokK1mHiy9ZAQH/LPURMqPn
xkeGd5rrkhhE4fdiU9WBC12guHANRY7carJ7lkg4YWRxeRaQncPhhNhi/qgI/N7ZQiF5CNrqugjz
lbReKBeI4hkP7Bs648D/V/cfw/yHIyXh2beKH+caRHe7Dsg0lD6de27J8FUzPsVPx7j7neYpxjuS
+UE6rqKgG18eIiv5ii//Sysmn23Pj0117yrCFbCAeBYSC8Mgp+HS7+O7DckAICnAE01YDqkIAmOW
/r3tpW0THNP4ZNbCQTwo7czkD+WLvdOEPnaI037WzWGglSJ7Q2mH3rs+X5F2OlJ7vjjO3ByC1NDm
I10f2SJgghRpPmf09J/iR29gBOM0yfFVhmFp4yTSJJP7p35YqqOnjJsIVoQQb+wKVa/G96L9XF1H
3EqHKxkCkYQTK+gyWe1WMe4Q6Lvxm5BIWosHt894KwA48r6XgKzxXeK8MJqTdbNSsrFzMlp0ideZ
8EgDn2muMH59/c/1yqzRzrdPeQyXRC79/Mhlbuf5GgcNrvRc501sBMjp9+hBGn4MXfKy4fX0Cl8N
xUaRE18J+cCQX/qKz1rLt0XulG7n5+bLde4hE2dCiY2Q4lznEH/UhPqFaTXymeCfKtFZ3ounyUaX
PeHGXFBEKeSSkwveIKvE1dxFp31dweC0YeL8sTAkF2XbCqhgmExCARPrdl/uP0hp3jvOpXd/xpKz
WBjsFfPZk4YSXrxlP8tPmjoDPHp/JGM/QF3TzaHMjR/8vdqYt/883oG+t5JTgEUFRJOPFbLe0ytm
oUdpTGJqGoZBFEOPrkOmEbLIGjWHl6yU85/xUYW/A6AwqTFz27/YQYA1Hp2ol5QLfZCMDG+IZnve
5lqm6MLR7Z4VDll+0kZ8SSsMR1i9L05mjfOffVQBOcDSq9GzMgGL2nXj5ea93jfHq2Q4sZKIKudd
DKzCrc8Ygw5puGqfALaPTEusXYHHAYarcqa6pAiXO0XcR5taEcPBB89GnnqugLPDO5Eu2RRFLt9G
8fy2y84jgiuNDuBwIEGg3wuxGuNvycFACs45ImkypdV3lVTXJJsnjeSxEorNzwxo5DyArOLqxUce
aHWLNlMrlMfez0r9lj0FkTfBD0c+ZZ8crj89MPqc9qC9lHGIBWjwyYaCDSIQTHPEUYCrGu9sB/ev
SgwLLMXph9PVsmfKyTodGR9aD15om+a2i6+vmV6I4OL5hWQIZFGQ8+nqRfThSN/QJ/c2FdfLtD/C
/ef48rbjAQ6lx6H0+P60yBd6Km6QJmJ/1xh+pBM8/dTP9M2K6GsyINUiH2wq58ZwLX+96Iw6u19o
n6FkBewfqMVFD5+aPbqTkplAFMuqqOimeAIXGP0tgRv9gRlYfUUGJZ+zqSux8hkVtaVv/E5nfEZT
VnuW1HSz48MSRdgvzDlro81wYE/arf2WPiOi3GYLJ7Sd9/JR3xUWIy50py2BKOC5wyXmhDMdjL5C
SQkRsS/9KEq+iu0MghD+uArii0NqDGlJemL90IAt5n0ux48OyyxsUzUNBVWbwBMUrSJrcvyaJs6r
GjAY4NoTakKlg4xQ44BKkWfVw+wLbnjgf493OKySR13eCAZ8HZtMnmRcfFiU8XPlGIIvPK5HXqva
lPm2zpGoGIZH2DP0eHshuF3SVfjbXtZA2qQc2yBj4jo6zZnVtrs9ekmU3sVhC19ma8tOjeYI+rOe
sgo1nncme4RHkfnekbOAlqqpv1c6eItI4kdtG60FO7TA+WR6u0EsNM7KCRcx9THj3ixP3Izj1rS0
khA0IEHjpyhqOj92kJfSw5b2q7p77ANZxB2Tzpm2tg72FhccVgRfdigHxAVXbBFSRhE3r/1Vhot5
eGFeCkqJtNjz7uydY0ZuKw6WEmTBjQAFGqBYNjRNbht3mcBcIeBGA2Xb/mkz477EJjT0PNz5oQeR
BsMeNmL8hDMY4AyH5fgnbwXdhXNjV0DOsjfuTCsWaeIGzKgIKSjuSAbq9IRNokuuwKKXpeY5xx8u
J2M8lQZU2TUTi5YzFz9hzDEAkGbxBfc2w4DkQOQymKvdMlfJRNAbxiGNxH0l+gTDJlJO5C2KqWhF
V8EGVEEJOsyHW1ex7IMCVNHemUGKYUeCxgpTwm05ZbxRCKNiPM4a6GfeaHGQSSefcw5MyTlt6cTi
i0iaDVVWPKAnlBmj5gBiKEmXjf1XwQDuCphn71+b18s9trLOXvn3dpRDbAILIhRFoQc5jfkkJGm3
GT9rJTNahEfRyrNHwcqVp7nQT0E3H/7ICTM9K5yAU5vNFwRDDpiICMSqZ/mjVqByaAx5wifePBd8
QMFFFubjjvjWDFT57M1KX94gInFDeGhsqYq2CDYU2+0Z6GSKTZNn10wVWWe6fVLIvhWnwr+gIvuy
hcJyTxhHqFG/SBuU/UAtqqorUBuqthvKZFr7Qul7fM2uSwiOrrW683pWuETkGcNTRSC3sf2rzZV9
yY0QruYOHt9tSiYQ7iXHvTP4JJFO2ccM5VJKKLMlB2qEad1nenqQ0KJT1oalH6wBlLABixthdq6x
9MQiA+Tg2uVd6zhd106iYlnzyHZILZWOXwhRkUztuygvcQ3c1i04q03GZToncDwQTJN+szlS042X
8lJ22LvdZBNywo4tNzBedZ9BF8FZlEvvg0XqJT2kfd5IbfTlKoui/xz3O8BD7v7AO2GkBmti5ioy
boNP97tDFMsf4Y7Ms8TVOQ4QoBLpwMyZve5uAUjKYSC3p+cksoMpwleqsK/DsvU5pJhfu9KHI6oj
nnWSYxXNSL+RXojpq4KNydqSU98srVXh67dp9mXgiMhjn5xqgaVZeYSNHci4BRlxrk0FKEMtUet2
lHQqjLHvyV3iOe+kFlWtGZEOJkjtSmGZj2Ui34hEezw2ebGPXhbsSaa2FNu8UkCYq2wFtwC+ijpr
PzOpvoto0Nn0rEpp2O+6aiEVW/wLD028hgt1Y/Svii8zH5xEw/j8gr6LDP6bnD5zJK1jf+vu+IcG
5UsFjjl5gSjvU0pOlKhM6HZvwGATU8K9l2FZuw8riiYVM89IGCsPv9pIofwBBwwJ2Ef3Td1XoOmZ
m90vOO2YeAxpPjdflk/zYCMqG/cVN/Hq/Bhuj/3eqZrPGPqSjSh/zxX9bsW81WIXkZyUmPJX2S99
luyFD6N9uq9CZ0dKEN6D4wTU+dYfHsg7XWGz3fgI5G3eWWobunzoNvqBkRtBixJ6fceMg1NCGufw
AcxGhdLKUh+LXpF0112CS6UPNvc6MDkolKY9F0tjB8RUSLF2HPWBsO9yRvSQcm83BU86xSoHK6K2
A/Jp8iKGVXbFmvcZEaRrw0LTV3JLxLgCUzW3w57GEm1thQMe6eSWhGdAwxOMkcCp58B2MYUqT17s
+R585TlbvxXOFHWG7tIRs0iRKDACWL+3FrzaE1U2bG678BQcJv5XuHWTv0HGAWhm4xmc6RQqc1d0
AdyzhPLCDf9qAocHasG+97sqliyIHE9fHRaGmlLXiPe8xyW7rahVM2qt/z/rHAT7+5pqYjg80Vlz
rxb6rRQ3zNM/oP8Hzm0gHMddJZvJVuv0zAX043SbhPDbxSveq26aXD5U3xqJGi/v33/ececLadJc
6hM85ZfJK7s69d4DK2h3u26NBdxAHKYZMJlPSA2rCuoPm1ACCCfHvz1IsMk2sfvuxyRR8I+6jSB1
Aw/G9wWhB7kppRzzRuOXF3XexaPlzmn6aA68YxRuEj3oslX0SQ+6SV3DakOMUkWIAG/sFatvVAog
mj6/SdsRqGW5YlJM7Emvu7W30yfdL3SpkVJkm2+sUWaB/3m0Exfahp0IsAVhVv9LubFDasS07JAY
WEx50f2QWh8gfzjOCyhbQRIhhTaaAUwrCbRuWqUqHrBit9yEJDY4WvtSeeKHtdma7At+Zx83kIhv
nRl8XAx4LemnMMBm8fnI4hdpxTK2FrKkDGKXFJyJ4BfI1LDnyd1GyGHlfe7ytghPqysu7gh00Oms
R9h0G4M6JlfTRDNTvNQh19UEtEJoOXPMG6BPqz2zqyh3S7FZzlwWsjFu6ly/u+QXO6oETuDRCFaS
BJOay8hGFBez0NQiHIBLKtVXJBTg4XN3lmsb+pMT6Dv9tSvXM0YvICK9aQGJE64NG2jXmpiK57ob
vMCD3X8sZtORzL2fn0qiwCGDATRs4pX36JJqKaz6N+TLvXDdLmkVVdOxHqdinmQoE0AvZpK9AZpG
E9E64ukiBIs29NFhWbw37VR3DBXcEkbNspsFFoNjvXjaBz4cFQzE4otsO8nEDf3pRXbrqABIDwP/
3sJt894h7qWAq+tt38wqhh4wMIbM+0sgHqWuJugTaf3nmLFQ1iEHhT1V/UgQpDH/tOPNVq8hWorz
+XxuQscJUrh9uAdAyzdYJRF9M7eElfOe4idFA7qig3wpW/qbhJrii9VADIq4gNsHnf6g6kY7GZR1
ChyL6HKZiBCW1brty/JsPLdOJCca/DnmujPGp/7ra/e8tlG03vKrZdBn5BrQyxsTrgmehpYFqcZ+
l8AiGJlAfn94vVEWjDtnwMfTp2bV38Z6di4wt+xiqE0OgZNVHMNNybVTp5Za4lTNTUnTaMhPNnIX
j/Kpjw4s3fnPmfwQCASDbnHI85ykusGVyuWWQFCzrAAQ1c58F2K2y9IcEk64V/dILCmQkEWzOdTw
3cM9k77kmjcEOzWMcWlORcJWriso96SYGHRlZI520OK3oGIVUUTcTFk5vBtVlVAYJeuuCVOsfOgU
QxuZbxT9drtoO5GBEq6M/ebMEYDSqrB3BdbvQiP3obZr7NdfGahyQnoDu5gtMjWvpC7un1mhEjWO
9HY4jK3p5l0Ab33MrHgn/Zmf9ZGdIgbFUq2Ji2wPLsgT1qAjoaBvO76GTP+Z3BcaebzKEihGrB3j
4AyR2mr9kK4SRXRYNsfii/4F6H5n7EeO4EuXgMgO+cjhzGW050TAPBsrkEHK9Ab0vSdL2vR22RxW
7enIkhNqPvPizazjTxnpqSzhJn9xIJUOIl/nkqTCX67gsaDTQALwRqxnY5meS+rX+99b699/JiGk
Wrj8Aaol08Z6NjHezw3ZeA/mn5vp+HDERKVc160C4l1Y2KcJOoHPgodr6V/xlklM9Alq5tgYo+3+
igEkAvKvF9iSmNhQJqMg0pvRp5x/V3U5AQ/gw9FcMcgpPxD0vxVYIZ8FqPYme3BaUDui/eXfjCKQ
X+/gAdRKnHtiDFf5gByUMskpXqbachmhqyiAXMyBtq2Lvs7Yw92MBuwgRbE9j6OgU7rt1KnmyMss
RoWSg2Atasu8gKTeZSU9gbi6H4eLz5ED1oYhOn2Y6iqUinZWOW0/W1VAZZCZ2tEBjJrap/NTt1rq
KGISgGNrVjOT7R70uP4XnqnATGGcwsIvs1Xv/tntZDNGoIgJhNm2eiSX1HZhgiy3PzuMqqNQUEW1
kFBdAIr4+ZpfJbhxVT66toEnmwuwEbF6yCCpzstyJxbjtWk5obr2p9beYmkBpCVqj3dE7OZa7dli
8ZuKNLNFXRBiIsuZmKcjl7tgNsQH4Nc872OA3huCOCggfP4orXFfKll+/bPGESUnhWY4HkFmOKkr
5XFgxjteJ2yN8p7/crKgjRwlfVNe/z+nAcMupJlwO5AmaKO4LNNFkSvAgdsGcfDqBmnOKuA93nF8
GHS4ryKNPujNr8BYEHWK/UhPpkJebk7pWzs2PaXBAmpC2Yr0PSsFRuUZPomRtiUF5sUQh+MIDsRX
bE3Ex7lV8Y/CRTKoEUzOAVNZgyLFEANtRQe96ekH4UpBja4qPajAqWm7fmTX8AtWVMFnLui9tmlv
JSFIEKKB4BsJwr6mstyLTbvBnnnhHcEzTX60v6Nb27k4AWZeUFVV0SmhbHGdukPbvZv2tSG4X86t
eMmIzh1VaBBC8I44gCgzaVJZD/1l3Q4nByunWF0WaLCHB2B37ULvLyt61AnKaYRs1QnryU36ngge
RnDOeDojTsTvaNvf5AjyWxGDNy8uldWa/idN6MhRBwnlB6FkccQPrwhm5JCbrwj1NDAL0H14Bx2P
BPgltrMTBCV5P5WTbXVUuD5LIP1oYVtxWdF9npvmJkZDfuWEuA4UWetlppuCDKwXUhzFSez+UYAg
/up5+Wzus/gL86CNVfB2LGCnb3vNsrv1YZv3BvvOt1Qb4L9jEfgIA4mCfn1AFIteUvj57srq60J0
L+EdYcwV/o2Grl4jzr+vjNktkRuUmSKj+V1sW9des0HojLNqacZ9K0bHDnK18kbFE9iKgaJJEPkh
v7wSG16Ho+BP89SzXjhydRo61IFb2Bq51be3tEavCWhUH/bu8TF6c4KKGAB4jD9g50SH+XwSai9t
5asQDOPuO3Pq5iu648zytj3Rotyp2QslzAhsX9oqj2BLQ1LJsk/KAB95hUtPCGaZYaQ98iHGy7oq
JYed2u7U7/c60kkSinbYWz0mEy9JD+Nd69EYrGrm9SJv93cHvOIT1ofpwMIWXCIqePdTte1J/Onz
H7yKRi6UdFpEjrk9IQD4OIhCBr4QxX7ulWx6BGr626+j0jh02j9uPsDZzw8z6tANlJ15K51toy7E
TLI4PFbtoALTcVibLgXYDkBHVQh5A6CVChk2a8H/8saQphfCwo1fjmWrNFwVdxJ/id66I64SA7S0
X/dfiSyKUippczUYCqd0+iC0/93yh0AvwT3wJDLrv939tBr/tpmjtqWxdpkuyGq8DIZhvv+r6TMu
xmJOGqs8bbV3WyH0JBwdOG8C36kzZ3NXW9FlkJGipXwFuSadpBcErTAhOIcM+dNqM8ohiIb+6Ztn
3726LIgFmnq5sUfoY+p46RYx37pKJY5Abhi9j2NL1FHvL70lC0DMNE5JubSnsxiKo9i4a86ew6vY
f339khS+rszYCT79lIBSs+WDWiuB4aGSkKnKHgGEA5ybdC9hFidj0JwC1WB63nYpgLNhVanbYP/U
SdrO8X4oGg5bs23EM27SLGsptMdyI7o9QCkHYqj10tKCx7RdUpOeEuyw0Ac7rSn+T8OEthlTHX4T
jWmBsKmN3bJ/7KwCLWNi7NGafSu7MIwyYtxdLuHoKnQBR1F4kRSB0ikO2On2oTWrA/72ibV9OJom
spd34xhj8pkvg9jf+BzfBmehYRsoSduxp8i9dUW/NJFihBo39e8FQ4E2K9BNrCgXUFVGCNzg9J4i
x4fKw3SCmDw0dEj0LCDbsQTbeMcCr+/NqwR2Rved7P2z0fGGBr8Ol5s42qvdfhJ34casy+tYpozg
bonrRIfhgHnfEKZOLLBYuQWF/F0SKl3uSybZXYhqVBSBsln73VLXx6tIG2keKnN2XDPKFoHLrZpd
5w2Ivfj6v+StNeZ1B1fyNJT3+xCRraDygIVB81ggZY6zppsylntpNaNZ8EwDasC+9mKD4kApF/8A
cLRFBepP9r7VrAUJ+uKUDm8hxCu1Ih/8g6ST7fYzMdPBwK2GwQwrmsi/jE5Ye9oq8wzAyUCc8DOu
Yy9OMindGAgyh7eR0uacvjYLVEKYwFzReFMfI1/tROTq7nmBQNPs05r9alzswxPmyDlvDzPV9uBo
pwAo3Q6Lx7JteZ4Zl834qt6N6hvQwsAYCU3VFc961vm6iqAT9L086nnbBbjJ587c1OsIOaQpjwKY
QxWrbjSpwejpjAtHKLL+DBNmHTPu9bLPNV5tZlR/r6W80UmkCmaDTxLGFAog+6HRPUP6hKB5VS9P
3MYMSUOaqY4k089Wma9VGWM2zIJiraDpxNrZ4VLVVy3oWDP0wm+DXh2VxwYuvvS6bx7nBRtt29tC
uLjc2V3OATuLYIHxANwg0LgFa0y/Hc4q07Krbmh6xvq+Tkcmbm5zjZjnewB5FdK9lSwjvn3qbyqM
7leRd9ploe2XVvN9V/SUm3dUq/iv/849B/0EcyjxxTZASFLkmg4QIVE5WZl37v8DuPCQsCUhipum
0o1mpmn2Pz+SkXkG+/uFB926rsKZyVSgbPFW7OQRz/3y1eczmmUEUQH1Us8/7i7Izx4GWaIPYboo
7vUN+kElNsv2GspZ3T4VDB2dIza4tyx4h5AipsbNys4zNDHuTFBq+xwKOsofjYbTC0BIpYx+Kmvn
TAUwbLUG5QnQ2BVhO21AM1NxO1TMaM61UyvwneszP3Tod2h5qA0j3GYn8CiGY5VgqU6PVFCPJ91D
GTHNZnXzU68DKd2nmvIMxPaNLGIoedg2jwd9anctNzvgC1nY44TglxbuxckTiD66J76qoCh4xt+0
n4ZEcyNO36G1VPoH8ZMVQcqkmldmzd8afmHHsDVI1ccicy1Z5dmlWBfTAQX2By6BhbrJvw9QWhg2
Hm0sBZJq6fyjpn6qeJu53bd5gTBUk//TTFM4yA5t2tKouNFOmBfIF3St/5HlC4AOVNxxemsi71KL
6KewF/mCWRjudAYhaur3sPrfBhfjIiBr7+C5B9fwIoaRr0P6FjThOOaX4S+jH/Y+li/XRFM4OrPl
d1krGaLgEymslgogHhpoYAHeaVLBxL++v/jBUeT9eqrZ6hm6r+H8I0nke+Z3aUABC9SCVbE8dBIT
4TrA8eZyZL7MwI58uAMiBY24+J+PrzxqDUtNeGZXdjIjPtsbU52BZ3vuWEnKxpV7Mv3ZRjCMhH6z
P2SiKrc2dN6c1Wwo8tPTfCzoXyPLtGu2xXduKOta2IUNdNnZywa8MJlPG2wdh0eDL2I8abIEdE9d
wyfVqPm+2DtBqW/BE1vJhujPcTsNIB1vjMNY+WpjnBDVSBkfTiID++ceuXQ1Eu+gEkV0NxP6d8T0
8zzELS+3jcHcIByR6g0nDW4KfuH0Z+yk7iu4l3M6gNKCfc/mu/7rDQ6C1aWLBuP26mERGXlpIPHU
WfLQ3IyRQLdLA0iEeB1bubM2FdNLbQBoFxbbiLOvMK7zuXLw/1i6h29qjlXB4JrEPuB6XMcKwi2Z
USEQKG79IPU9Q72Xo0tl7VERdatpwEUsJQCjgKXt44O77WeY8dVt/RLFXENfLtzBU0K/O1fgzZC8
soBQx3/0zteCck6z1RwFWcqnHHqFVB9+cms7KSRypwh5Mxlp+2X+Sv7bot99GPZLQoVhPJYMBfLl
TXc6U9VEraUxm1CIzKtnvvAkEmTHzjzF7dqGdCTHQXv1XD3Poq/d56IN1Izr38i4EsTq7ZBPFif5
c3l3MIziS82jUneK+0Vv64lm5tpbAcQwa9B9AsSVuUdt2wQmlsJuEQQExS/P4XnRfogtf58H2+SD
IqET+t2wISSe2+tIum8GzQRMdwnaESCw05EeWOo/wDWIzYka42F5b5DeQKi1CIzwOO/p9knpczMz
hzCvvVUDv+QRaKLodIDObl7lIRvzaDyALpVRYFkaH1VucUFcoi0wX5supfYdDF5U5/VgpQwDhJfu
N+o2ExIEyI9GAbbmIYmro2KNZd2Tfhc4QekHeG2uMgdFRuA0hnvE/HSX2sDzliILwB2Oit2CztCp
sda1QlT+HhZmKbk65Epwys0CFymQpQqk9QSAenHurNd1xXolSmJMMFTTw2TuCSGj75sYw+T74cBJ
Oc5LNqB0ZIqVMerKizbeVDiLoWDea5oHt2GpUVJz0KMlyB3K6S1YN7BithGFHATJitrIb0yMc+xo
MoaOxV9/AhnfJXLHoSgxh8ncShecWCkXL6+rAKPEzeiixYB4hUUaWKTzcb3zfFbJb03zHNpFIIC3
WH6lI9ZvVpCz94JyAevQI+ZYxuOOODogVE7LwJnMMVt84xB5TIUmt6E6EyxuKdXsFeZedUOK2hoU
nD90AU3dfqf9pW+BPSmdkjvSITwCCK09VIfB0icczlpMfEdG1SvWlXvnigB6omNapwmUNy356qf9
pNDuiiJNXxIdi5w0OoMQpJxyJI/xVUJyyQTXI8zk76+lTvzTYbajgLkvbnPFdnEQlo/uoL9GTu77
SK7MTNIbqs6IKuQSgY5A5HZoaTNonoCWszEKComdUh0Tmywe46wFTXeAyzeo6ouqnZWInaNO2nHd
b4qmOpCHtzhiBac+ungVM1Vye7COH80Tb0QJEDgng7CDrYsDthLWw2mjm6hotKoxQ/TbJN/sPNY2
HC3rFT83lomuuFtouwumck1PjcrbOUPPhDb37OEeLoU3p3MLCXu2efo31s4tQJRpmJzvpzJl3CnV
TxYfHyOQRIQaQBsENrlLVmRqgSlEoXXW+8i+MbzmxMqSGfQ+FdEOIIBX1fe4eHV+RjSoiT3kDY/M
rshpdF89UyIJED6wESnWedOEf0NYoZYpGm+05ncL8fC7SDtQlJ4/iGXAn+ajd+K1XwD+qlPvmEzp
+Qh1yFCDZoTruDWIRgj6SsC1/3YhnDur8SAFY+MScHTkf/WNhEOYU1rb3JkbfJWpP2wRnRbtCkgg
6qcllmg36nrQ2dAqSwn/D5FCtR7T34Ofv8jD1WOKzGkYsvFTKHccPt1G2TVzpLp2M50weFWPRCko
8E2F1gFD+szJj7mNvLmGQGYr1A+8fkgQacb66F0OWeTrq63qfGdo8kfvBN+rTqXpq/JmYb9GC+C9
NbNg7YiYf+Haih84IR+qZygGDWCzTfRJDAztIkFpoxSTDM/xM1Yk+MES9IqOFOCxrPTm+DG9okkB
yuoilLwzuloXw2VzJuWMETaeYCWvDrqDx3CyDpVX4HLv+8t1yKqhcBApr0malYNCLNO3DfbBEX2o
61vLzzkv7a22EIU4xdhOi0dBFzu6taHxjNSie99eea068v4s3CN3lAbIrkxD5KlciUQvvX4xjw2+
ZLx4Eq7jh3GyuS6RWbGWkjuKFczz9dM5A3TfYL8jAVLHODSTES8RPjzeroaQqTpF+sz4XKXS8zre
6cBBzO3T5wlxiiX59OCNYoLRB51YClSsCCVWABkAFcgL8uvIKdL2gYz0UgUCtYrJu9NdfEOLJg+a
TQBMUUbJeeztEsuzJSskHdS6mzliVE899A204vWey929BDx6Fl1Xy36/LKQUe46BxlPqSgXP7Y7H
SlPLubnGS8sJJBtYIy48kOSHDHmtn2/X0kBggw+ZLx+1swy757odxdge2SberVC6KGWGwqhae1m1
mDgDBmaDr6ro3QyDsWFpV6CkNOKU822QWESHsZMEbALrcIyeq630naIoFsBi771V1+mMhv1LRt3L
qo8cwzzdKB1lAXQEsTGs19JM9PoWs11PzB6VhCfe+D4rkw44o+UgEXHNwrYiU1IulSNE5N7NkZDu
pnunpgEOKjm3R6Vc2vpkGlJjYBjbE0oXwXO+TVrjAHkj+lHgCujxT5dR+J1eEVmc6Ohd/NHoe2aV
hCOxj8Mw4kUwfZxZSA7Cg/Vo625dlBmhz+Up5mPNqkwphJDuHOQ9GOPzCUPdHmG2SfedZj+ifGxS
X0R/2nFmECigYDBGbbzWwywtKLq7E0M6k0nj5IsWdPHbeyZqVL/z9ify/1EM34kk2gtL0kwtUAKP
qNsbGgs+Kq++FRu1DqdJJK+qdVT2i7ho00arEUlRLUhx5lkdFZHp62ef+4Ck4/w0o4YWn9nOrSVr
WXJYiSV4ZH4AKPv1CI6QvG96kNuNZKFdUhOobbimBCrsiSG7hx+4mGXq6dz2U64y+A4GlKGjwKLx
+he+doqF+XcDb4qn37hKTKAFtu4dRnjM9xXTJpcDIBi2QKriPaLOS60iDHeIkgkUdqp6IPytkEkG
yjucxGnTl4/SS2So/KovGjOUMlyepnPpvEtljQnfrwNcQaUHeUtI4v4+8gg74XXYHbpKjzIKl6bY
GZ895zZscpJOFZaDUvfrBYmNrG1C0OLQNkQErOq50sdrVkup2fcP8ZOksbVG5Qw0DbrsPBFTzTrt
KF8SsY6L1G5KmyHMqgtAZpWBLmFXrhaeJoopdMXTpxdQCSzniaW0kWKaiPQJyyuW989YibK1hRw5
EIWJATmTs1jp7vSBozF1Pa70VYxJBLM7HemmPSQ5WMraPcrbBRylmGWe+/M2VTBdOVjrNYxhlOD0
poMSEEFD7EkV9y8FafgNtF7qwaz7trXoPH7NlGv5vGRLgNyxKIVBc0lH3tE3TnLPCDw0Odcotdpw
E19uyOYlZx0FtkFMarvr0fYUp/9hbuowT3kcms2ChZvIhjP4q9/f4/JhQIgXGqv+gk4yqHlku95m
D/hcWjmY+gXrDkhFsXwc1gjN3zH7jOCbz2H8Wwn5+NvisUhZ/3kKqbBEurH+YFqOiSeuqEaxKgsR
BFgUfrrq8Om0Sfk+6M7zjbe57RCjNrhzKksqc6DhdXjvNYvQ5HMHtzop4aj4/Ml4ljHD7qAbo5Tx
teM0ShTSj0RDXekYUXRTbXjxvKBwgpcoyyTBKqUytzcEXUKEj983ikRVw2ypxcEQVPjOZ0ruWn5a
zAzHYrQC691OoyQqKzfkL4EGd+sRbMxd/f4gGXLcbc8PqKUJFH54jD+uZpwu/bIT1AHzWqA6MVCd
DYDXsozY77tdj8ZcCHpxX/9hnjymSesiLiY9PMxsWsQzqaOiqOeBtRKEhzPMKDy6lQ5KbFh7Un9W
j6SmJtMGhrjIjDPkqp4qdvQMGi7j/1/N0KfLuPRga4+X/BgPOD6e+BVE21cixEiykw35aJJYyUP5
7JXY00qUfvjI/l6DMNDj5qjXrXg27uBDzOHlzI60Zymx+VulOxn5+5Vc7EpJFzqL37baX+owzedd
5GunQ6iFDZRvknYRvbvCKp3LJ82hQUBvdU1Lr3au4JAoRsxEhlT2IT92q/ueUJz31OFoyk7vDp4b
lLdlQ33LaiCkSmKTvnA2gTl9n/US8XZpiF8/AD51q2h9qBpOfWGesSs5tArakP9YGKAKB+JGUXLL
8fbbYR8DL7tR7bWff4JTTcypX5n+DNE87lbHLELgMwGSi4XeBPthgP5LeCKSZYnodyzrB21cImMs
NC4so+mbjIPp2ZuzLnwvo3IzAPoIZRfLnN3gYanjybfQvceq+cQkexzUSpiHSB7wJqM7I/p6+3hl
BGzgFg+r/CiGKbQF98S8rm3a/7sjD/swf7+orMqvz172MYJIZ7rqOzm6vslzhVckqDBLO7V3kblr
T+NhYNfA8CDKynSmjK5uRZd96rTWzwssj8Az2s6H1z7TbGTHbkG0vaw1wMsAB3/3gHSjYJqTFBU/
K9unNzEkcGFFkbVwUwyZ7pduBhd6O44+YTt9p0yObbLfy/mzKYKNbfE+aex2sPhQRXR4HwD5ZgBj
A71vK4LWULxY4shmKrIo5TI7F3prmyUeFsQnTwK9giH96SLzowQEFqhVSbYz5kW3xZZvH4UTQZ6G
Quvqe1JLn6xbQbfKx1XRvWSi2tyTYc8hfTQ30dpI3VbyBKQyyCnQDbxUnOpQ7TuFm2EhQVaHdp/V
O42Ljk87iude5nAFZOG7N7Ga4ZL3gVbz7ZiBFcqlJIdgbpzTRVu9bqEzzgmRs3ph1FdOlgEf2fep
ATQqJtvGqRRqUjwiVEFMNLr+5VqWIY38avLfuOv7nCEZ3lAUllc0GoXp4tgc8tFbrV1EtgTnVCeF
/boP8IRpMvEutWuP874CjQx3pjvi8vKc1kgrX/QS6Kz0EYi75XSs/0dPDxdVuGxK43TAd+GNNJul
ynRzG3kZEKpzzPrFbUfF7SCzDKxXwodFwwEuVEwn8jdqlY8Z25eHTuKSY+Ik0W3h65qP2adr4vt/
WlW7DWEWW8thYrSR6BsDLdVb7Yx946OAFVkGNGGoiMCYD/kMdm+MejcbHxLMbeWwlUSBff/aZk9u
hNvgf8SUq7sAh0cRhdhw9fIjCdc/czoDchqHXMYhvAyKrx0OpX3mp1lm+o+urrsCmeTi2/aCpaWm
Mt/dCO9U897qG8CiDlSf2Lmyq9lubq8p7CLLGZqaJk+cZO5nCIm9NfXD21M/CZMOZzng4PFB5qBZ
Y6T9VFyVKQQ/LqiGLP8k6q8yKuj+BbBS37mG42zDbhhJgd0vSr3U5AEAxNI3xPxz4Z1HnNtvFCox
JBOzdyDmBWA0odplepBfG9iQTtoAiy1RcKcQjbjDdROYdXUZYtqkgIlq4+YdT4BREOaGBusF9xKj
8icdBwZTLiBlQl2PKgTanrtU04BtCBAFiJBinvIAWB+pU/v4LvidsXTxX1zgDUDnQ8XQe4OS9eFB
OlqNtCR8HPXpSIZJYT0c7Ovhp896uiwBMVfJxt8zs53jRTk6cTxTklnK0OyTYduB+buFU/hU8gWZ
5h5wwkhfgaQHSuMdz4Wesfq+OehtZwg3luEMpuBTdfedfxxJmp4Y5+oLpjFQTe6faDksV/ztZeDn
u94oLCA1jGODS1enwBve7oCFZG3IMTl7Q/r8oWaEbuM7gP6k+ZcuYuPa8YFk4miQu9r9IXvYz3Rv
Z60lOXHN5vIBUzEDWXpsQQgfaSAcxnp5sekGaJbApMbt4q8gNhx+TUM9p6wC/fBnlglk5A2U4x0C
YNNQOrYgL2LazfvsK5D8iVj9fLBCaemCbrO5BeslDusDCKwoQpq81cHw9uOtdw4jnNojoG8B2sNJ
NGvNcrOl01M9/MTBdlqE9WfVRIrBzX3qWt+Qq00vJERyapreOLz1NyZVZ7SwhWHdgNkYEAwqh7aE
GtUWsEN3lAERwZ9k6FLzPDEg66woQtnLf6dEY9FTVIJso4NndxzzkMehpF0UWnKLpyfoarnMDc6T
Fnsk1J8G/sniOhL5udPI8UuoMyAhsUpcdW972jtxxrp74Roxfa3xbjxiS99wnp/BrhCe3Y8hyFUk
U/vr0McYWPPEnQMcBeGYjN1uiEHUQtlv4wERUI5sAKiGi95b12nT+Zq0Dv3R2cU86Kw9D6nPRDs+
yTRAiqfIgQuRP490qVm9tJEf2T1Z9fHzpEgjs4trQhsHhKXdBHS0B4diKq/nLDfV3rxyewDehPIw
0IJ5ZuA6A0Ewk8mjF2daNl84HBeiDw/8Y8CcyHsdWYOiwJjoEooSi21jf475m2e5JR+auAOrKWhX
DByc/va1aUHnGGCsUae4qf+dicUqCePN9dnzBQPPL4N9AzdnIHXdrrN0K+qlEx5oeYGhYvpkf7KO
6BSBwrG8saCemdhzdCXKNNKqKGj+pqkrPu4Gjfg0MU420ZishotDxvoVSbY6ubiM4w21TW2d6pSh
X/K92NgN454HhOcwSx8aQ1Yf07Gcbml++xBsHuwfshYP9GmoxOmp4idyeGZKrN5kX5QT1bctBKJ6
rV8YULg0TfY72wnrP2ecBew7hfJnL9S0MhVlfPekDUYIbZqGhutZrp6LBiM7tDd78HicMcCM/sbj
3oAVZ4gimKRA1NV3iCpX4WruOPE8a812VryGWDxWeVnPJ4NTuxIZLBXnSe2ME41CT3vpIGqo7cq6
dAHk/o2jxKUIpamQ7SXqFTYag/6q8npy9bnP+xw7cUQvA7fHSfidbesP31+XKSs5mXl0rdVDU74m
2y9/pPxL4HvOSMKxRyzJCYaPjFCHB0y2Xbsq3wnTBbq0afuBY4FPKip0pjW+xQk1uff1+yJcMq1O
j9zT663uihzqel5EQUgAakz1jQIZ+nrvKeFIF4ZhVMcOubM7p1g3JeDT4lRem+ejWmeAmJMAaVTp
rrpFKcYsDh6iBr1YDMC6DwZPTz574WQxA6Fen25kjkqJfw9YciAfxiirmX73/glzVNviKN4s1jeg
0QhkSUB91UZzFAW5CXyQbsLMj0OS0QVQXQxCxDUnw2zbD4oJJS9oxvOjO82oOqyrxq1wKSnuSj9H
yT4pGJ9hsTYl+XqRfvUtzOCuvCkfpnaN7N81MyUfiZ2sE7q7ipif2V8TOXQNzgVR/oP8L6wGS92e
4JgaG8gKdj1j6WLehV30pLOKr1r58VFchj2qRTG/SEE1tts7EYUJj8cFpwKBartNroqJtnIn07cP
KA6EIS9KsEfEi8b4WRRqOvCEkoLunxLHC4Grg01bbxOIytHzJ9YNJfRxTr/KvjIAmX/OWp1x47SG
9qZtN4aSZkcpoDoI1dOb8Ln5RKl1lH0l7U+VFRjEt3ju11tFYhL8SK/fZtww88CHBMePHMCGI+v/
nnAZ10fQp59iAQRgyTc+r9L1dENC5CoTjDTi5hPx0Mim93vaNTbMVBSDqDG4MnDG6jNJpdrwgM4C
6PDYgTkJeFz3+M2nP74sEpgBphYMFIhtqht/26yxP7HJg01dp13ctKXYmhRm6/wu8ETEZ819FXWW
tnPaodbzRLMY0yL6qmUXzxTOaWTDNPzE6EauY1SLBVOJMKFZOqK83tyCyQMXNqtIslDV2zYbRFXm
Vs52FzTPkm9Yywr9Xq+LKpmMTSugfiTfZc1WWqa2AbwJOU4r+C+we/GCeiurHpqmX1mC9Ai4Nwr4
YqjhHExctpFUzi/v96s/Mdx14jqGeLBfIIQo5PUa0RRwFn4iWhj9e2Ug6XcXH/eFGHhGVV/AzM+1
Xjav7fwhLcTya8XTlbuBTbj3p/eCDQncC4eeYngl7XqFqcEf/M1u364vSpoyHaHqWxEs+hJgMNFc
TWZRTWuFpd0wh9A2TNkSsN/Ap/RVVYxUM1TdCAym0e1rZ2DXwo7mhEiFlnbgmLf/CIT/ZKMDjY2N
2JpKE9aWbmbojp5RwWi1N6jan+hEMO6KXKi1OOoykBs+j+P8ek49c/p52aGvbOx0JyW49J87OMD4
K65i/lu0qOhPaszuPTMpvehHCZTvg0NEdSotz5ZgIQL5HmBCIFwWQ1YBw6gAA+C4B5pvgMZkDLUq
ppDs3w1OgdezaqhsO7P/xqV+E1qa3HCgwzbnr/PH+GJBJP3AwoQp1Pas2gDuFSqUqUGoV8FBF4sC
I//oua7eSk+iaB2xyC+OwAKsVM69XG25YRhJe4ltPCBAtiJCSDhR0T8QMWWNOW1pSO5ZtbhhrX47
lnYhq00brWy+lXKZAKQl5DdL8YYLVXSuAdRDnGJdkcs7P6dsdq4lIxqQaQUWGA6ilX71xTN4USTd
Ujst5yOrMKuGWELLDrQRosTAmxGRzpIFyF1FwfLxvjvORZKMjBeVT6ouubjeqACr9jPQUMcneGix
p9KWS9wpURFF8+JzHvnktsvfuY8Mq4RGTZ/SCteCic8wbMciIKx/3qP9RTZ6Q6C7oiemTShrbYFX
WzuHGGKiu7VVq4VB1j4aYLPbYvWMzZawhXqVKHdl8Ooc308+y0gL0TaTrYjsR2DVLcNLLXDfRNX1
+FXiiHMqCeNYHHNHABdMwgKvP3jQB8OCkh8XfF4xEggGlMD/VW2czG8wAkPcNQ3I94KkJLzpYT0z
+2nqdRxaquu80ukawD5RfS0bqheSfRmTE9DBpaXsRpsKqhTwzZ6ZP8/3FP8hJMK8JkY1+fmdeFwD
rsqPW/uT3zEjOzv1ubH8IRMX4Vh4SpHAWl5Iz4pZon4PnpuAAH3YW9lddB/9CMdRy3yppICIw5zf
fqDtvLGTlZEFebH4vCfv+2MtmTUOlU/SUyG+bzM6e/CSHTTqdgNpPYaNBCvX36o4FrMxnwk7MMU7
lbXDHzZkYbPPvynbL4ld8cbKkr36pdmPS1avc3yWfx4dW7ZjC2Ecs7eLPA6+4QECRS6mQB3ay0UT
NzXvHJ81hpSgV4tiia8SPYbL0i495UQPBhOfjkJYrRiqK1FQOaf3mvQ6O6+12UJteXOuTst3N/oI
mR6FC3ATY+POdK3bUPWe8siqB6i6I5yb2NRw/oNdwAkFlUKzVcqY5rMzwuvV6PiSG896mr3X63v4
PeBE9o76MwWOvRV0ri8MDA6e0VJXIn+GDSmXWp65Vhjv+xt7gUL0wC6x9zSfn5oBEVcG78+OLSyV
oIsq0+izIjDzhiSrthmlhoKr6rygw/Jn1GTEFFqmfxkvgLIF+hY64RvllKq67KRrqmqOPmRQ9QlL
dmf2tteQHT8U08GpDkbMSe+V9kXce1Cxi4n/IT3HXfkt2gtadVDhs444X87QazDcGHkjib+6q5YE
jd4b0HM64gwH23271IzBrGNmgEZ7i0OHZA6wWTAJfI0ka9/Usp/7f3yYpRfjwJmsrPTsQyAWk9iq
5FsQjl1ilaOYMpDtnG21pKVablA1EXvWYpl3eMSw0xhkAi5Sf8lpnrCaaa42ch8/NobWf5Fas/oG
o7PcaaqV/bHnKrQsdNctI6d5YZHK6RQQL/ggnMA3DcEJSEOV3ApG6Afx8GlekxDKEBDU2pVU9Os1
AIICxbmhYXcUgaU3UtgkUr5GkgSnhLPvK05DRzxoKcuTe3Z0ey2kjPfisA7R8swwQDi1CoHr0PQe
Gti0P92aji9W+bKLlEFJ6dpZnkr3KmKheLsFvGkUUXEXdbRo7jq2BDBTem+UPekC1mLJGLAPPTFN
3sLanYmtlMm03U0HmyhDbh/tBckBsj0Xzu+5KkAPmFsbImlPXpxQnssZGasx/aP6R8iz7/npX+xP
TwTJsOXymWz1ZIpo1bUGDfek65p2s5+3nE9ftCy0sAfLz9ESUeN6XfJv6kaymvz80uKnetFyjp61
5mRbRaSnr1Av3vnXLEifNt6IqeWZeHN7aALcsy8iCJVEg65DvpyOZB2lBoRrGxAtzLixz1lZn6VT
8D6f9TN0bgbucOQ1+cPP//3RMpWlTnrawp4tyQXMsdrX0ZHLvASIsCzKuee+/7JqK8tMvzmZOBb2
dqWbsXECZMTM3PCf+3a25nFM8Wcyz/3kCV6GKU/cE6RnjJW1PlZVYi01nA266vuFU3YlYaJAWi3t
Hi1LM8yeZsKeqAq18Dg80xPzZXwcIL0IGSaw5Cyu3aMNOrvYR1rQRTM1S+nOaPKl+qcXaa3Aum3c
/VTscKOuMCuhaFqska8hIJ7HQAWYVdoc++w+HOag/Y9vKPw3Jv20fINx9d63Gb6Wlhw6X4d7FoHw
rWslWyfjm/W4mib5AwH5RBHErG7t9HtnxyRwmAoDVUbEVFkJyCVbvDj5Bga5ZlE0M8WXv18hlJnV
ltqabt7VcIoDZYepXix7zhSC6PZIuh1uwwxSsAQewMsNlLw35zRai+NEu6aOBFEewTzmNiXyUGYL
ot4VSP757bIVexxgJgqyXRmBSXt5slNYuk/+GKKIkfk8j6+I/gjtyVS5WwjOrwucuLf6mNAfSDtl
irS7f5vLT8zYUl/E2BmBeB6SoCWZ/UbxVTl79jcS8tZjYysW9nN2KuwxwXTbzqdqK86X7GX2pcEL
+BSYFj8iiunO8Jt3AetJ2pSf1RsRRvU93iuEZjL+MRJP7bZoMD7skev+QxVQk2DZ14Ld5wQUbg7+
E+tg+/IJnmm9NevS001imwjR44orDJUJYcK8yJReos5Djc3HBqQ2cnfrWIIB5rpcXPcPDAPyDDMF
fivaSxiXVp2iAlZMbeo6zKag/gcYFl4incwTamikXeogOb1WlGddF0Ou9CwtLxZvl28n2CbpZc1/
WAuZkrpCrkipaNUbL5+nA9RoLkxmDHvWCiHjNaZcLGM4nsNBObNqJgOcV9EMHUHsWQPx7qbqm10t
l+ogiltXjqTS/EUAIQLAQ0eZiZFWY+/Fp/CRO3CDvLVcAAPuErxCPvjnxkMOqFCzuC4rXvsnDtYm
8yc9DcG3oP+MLd4D+oLhciwkLZxeBjvhkYfp1BDQhxs5t3xs1i6VmSjwS/KxlPUur4UaFYy73svE
z9A0kvUSDq6Z6GbpNIcZFEa76flNgA9va3SJTAdmKHuP1NpsCfJq5WTWUR0Atpy4lxAf6rsekyfD
gWiRZOISZzNdY8puPI1hXp8jubQ9c1a/h+JJkiZsj7CfTtXw2j+Fo/Mt9adI/8qSUoIIq661nxlx
NfpOO39Diij11e2WzOJI+cJ/SGX/txQv1Mb2M/Uc5avTOJcExl3W5cSonWjRXSpQqchCw+xuepaK
tncWnp6svtR6FeeIDjGFc6BiNDo1pGBNapyuh7TFTD2uDeTWY/WDUnvb33OJ8dA91gLiYkOXeszI
2NB06rBekoWTx1ghUyRA65mrNgqNS3JvtDpjEUYszFNThduBUn4KRt1sBp2dPbRDN5jQ3L/pbEud
h/72jUnysoaoaPpfXxG5Jt+CtD6FF423e7B3Ej0RVzbL5whOL+ayA517VY4JAdcLOwxUDvaec5UK
5bq1pMCOTAptnKcCmnlgB98al/9/SdgiC8D95Nb2+Re/tIBvttCspANHJwjiX4OoNY6wV0VzwApz
mgy0gA2GXYjX2eRpnEhhk2SFB32pocsBrMRBw6yub3H1yptlwtaBvOilw00rFc7IGgjQsQCnPaaS
IfXauCgeTBGXRR73pTMOIm+1uLO9LvSABduaeTaJIXppsMk1hDlZ6rPbhJyaZlt2A77RNV//OLa+
SE3vm2ZMGAzV58YR16beWihkvfU96N9I7oJT/pCTBB4DHdAGZulguFbdVzOq9BllvO7WqvRcjv5V
b5+F6UKhchXhcNKldOGQ/2BgY4sAYiLilw9pYPChRTVSc/qOoOymIEGvkmAMlbbvnf57o8CPL0Ur
lSOjEROuQIV7KHxhFoS4ZxadsPXf7usSDuA11p3qR686YAogI3GZCgsoIT3LR1iHU/1IUTEbUL61
jNoHkcU61yzmwEfQlavDH+xPLSecoX9nUL+H6jwH1Dr9VmnNQVCjYQx4FkjE9CLt/GHz5mco6N3E
xzuSBV1qzvKNyPV8P4PbziYzhMaXpMUN0rFq0BMH86878FEYJz64Iij0i07Jb5NgXQ9eBoL4YNRI
qDKhO6hD5GxK9r/HmeRqQ9odHbKqa7Vz/disqxGGWPTgJ7YRHtr/xzl/P3GdDnOSrXOoJ6AXnOGo
lAkqG4zWxxrT3QRypabwNrH1Ctc8XduOpzp3oPgMOPIcL9/62KemWVJJ51i4G/cQ+cbrsMTa5lQN
Z/lIejvvqdu5RN8j3x0N/G5hikNo/7SDwOrNI6dpTp8BQrpri57L/dsS+yYjsFlVGZP7hqdQYFwM
TEiDCyolPKay9ttYySTvJ87FexzIkSotrloJXTbJujkk7xq3WtYDqKTSfaKgsEMhTptFlAgdo5wI
eGeLsf0H5sdB5Uvgg7uRgsXPDgDKfrP9lIqhSvfxhaOrs/TR1A6JW30DWaagZnQbs8/hlG1l8GBY
NlRG39GrpKHu7hEXnwMGMYl5iEPMPtNq+I00GV8qX366RqhpYfPxutO0gG+d2Is+SJZxgCwp3WX9
ELsJNvi9zWRp/bczUdB9EeqouS8yugCyGdkbcOmAroJVmP00WpE3rCabj9iSkndG5R0wDhbOxWHN
f4evr35cIweagG6L2C7ciYE1/HKsVqzMwa2TkF9mGITNIBWfsHCDouBa174X5YWf880btwBKsdFv
LCsr3tMf5QRsGdh2y2vxhJjICetNzGDnYO9DXoa1wH2kRkY7NX5mgjPknV5+D8rai8c/+lwmx9PF
Z/sxXF4a22xkiGQz+hDSYQmub0QHGAKZNmJl1I5tB2dtUiIT1SdAnHKM02HTnLF02W5+wBKegHww
HmPiRTrc3kmnXucsz+kHkyYzKBb+UtixP6xbMmlXycTHy5ESHZKBQlgpPk5NF0qW5aU51VWqBjKR
THXUI2n2yVF94qieDGKz9Dro9gdc9RMGZiZnYPwx7nJVwyhhqUnr43y38bcmanuY7HIjpwBLytGy
d0mfOgULGOCRSd3IaPFPPCmq9Baw1djXxjTuQRkSLTshn3PtgHCpx84swC2+RJgVew7hlr8ySL2s
p+lMpcdD9o0d6FlDWUimeW6XNNFsaUVgu11DHyWvuikRxVNtyZftfuw3SdejwjNrBnnHpMza/niW
SGzKCCqJO4pMAuv40I/SChk+sbsJgy2583BSqdJl+CgQIcAkMbQlzV2YZCCNAgyO0OJ67mivanSQ
g4mkBUYHXCwR7KCIBVilpRVoBlXuIEJBETgC0rrn7KoVneRLZ93SAbBuT5OytSv1/SJkZ63esslT
Qf7V4SjUsk4LmEOwHu+niq9VpOMZma+YNtuIlZrhdSiPG6xnNEQ2I0NzqXNShnphgcHtjxFydtre
vQ7U5oMmF6GbV+NhcRvuFPDneRXW4VDIDxHPR6Xeb2eUNV9yvn1f/bY0IaRztUQZeqxo/IGGSdq1
wZKc0QtYswPvbcoEgr2w7ZnZovbWK4y3s8GM33jAoRH9I7nCT9+75PTvCdTCkwVsWxfYjdDnyEMr
YGNXa+wB7yasWZcaonYkn3hZq8o3A7EBTq15a6IdoL5iajtBR33tb5V7iPxAhDypkmBcq9y/owJz
aGrKFLiU3hYh3IYCGYnhHQP3gdn75uyESM7SXVtLZ+gjpKTpY/45YCmTgZVQxoA7MPnvvrHZvC1d
vfWFRR/xsBPaCAVzpwcN5pJ96QJDFkeqbiXg0AEqEcsCZdfaKPQekua9MfyLfpOT3xcMsL1YUpBr
NlH3SU4wSMB7vsGeU5YtrFqEiQlSintyoIAaq7NfckjP+YtMBsd7zhuKVtk/Oc1BK/He5YFObyPh
BCwyXHGKq3+5WEizG5SjRfLEUoYcbFgNcg/vjRftc8dOCqD3TobCzvSN7TxQqR/erLUzgYikdW5U
m8aUnxdea6FepJ0OdqsD/SOJM+fblySvd8r59vrh3pCEnbaIt4sYUOGBFUvFktqc0Sl2vlWwgkdC
7gpqruP/+Os3NXGR+HWv5f5GVY7/tifD9qy6bFNSZQX0eQ8hhRndw9vC5Ji+qFPahFGsMcjq8Twf
jEHihYjEPGiZg+aCm4l6SFMeYNSG1apXxZn02Mh8NNwqzI8/0jPU0uf8CcORGBPO6cSvSXgfX1XC
FVwha2TPbdQXQxTdsC+nR3qd2mCE0sTqVglfA4jfg99XFLtxjMyq9ssoGAJkfk2tHXGoSoViKIoB
2UMqeejV4WMtyHwu/mTh+6/MHKWgwMG3AAmM3s0OjbcNsr68xwDqHOOnw6fN/79C3va1bQHGTTlM
F6ykQNu+ZvtyDb20STOB3WsQGFXf2UmH8iP5NtF7+OdKI7n/3OS6LgDontL9hcrbfj75evkIlsQF
uusPHHtSzdLmCYVx+qF4tdMaF4GgVOVmXqeFubla6fvFb1yqT9qRtGpEs6t1vVBXll8J+e6SCRKu
QBLB3ogRmIhPFVgfAnuE50RtyGSjFk89GSXCOG69H6kck6Bo++T5bADiNhzfvwVNSZ99GolWCVfP
T9Jp9EyLrw9F/gwkd2Zbm01Hhz+g2FcOnXLgG6X2Mp0Nrd3KY52xoddS+cy3yIf17p0N/zz4IR2J
4wZcQjBawQdS/OSgyWsspykUrlha5uHabP1sc5t8IiVtboFo+LVn9j3cX22dZT9pN6eF91eykXaa
6+8QpIvK2IZJS/NxQ8Sn4CUnUekhyxmo5QWnEFa7eH5i5MoIpN17U0XUfE1JB6ElBbhug7NYVJAq
LJxlk6UfH6suHhvEZf8k2jazh9mDTLqP80HH9DJpiK67NFky7SWV7go8F9A6GlIekNn8LL+tVmJh
ZpryR3EV+Q+7W6VUh3SSoF8EsFh/vxxjIAvx9d01l8OuJwNmFkQAHL8E3HwnbFCb65ILW96OuYux
lRJtzm08APGkaGiPwuvC+eLxtpCLvCIPU4H+sm0T7AwODDbKgdjJ8LD8w+a8JIcVWXhRKw6eWxU+
zw+yt03+fTqE1UT0N5iqGYrK7i9TjB1bMd5IE4zeIRHoMhhF+wZ+2sLM0KjHh44HSonEd7+hblsB
KDf3bg3gB6nfPHnoUq2qOixKZwhdiI4W+9PwBEgYCvruTMEz3xDpRG/3249cpsH9yOGv1jUGxd7T
DUhCgso4cleWELFucVVCL2Lnq2Z3HpRJkTvj5eXKXpkbibjpJpwHEL6KaMUAn/81zdi0nL3FXrmB
FWu0b5hA4GGmmiOHArWKi+eoFmFYxmb75xKjNZOGDT1+hf2xgerqLPqYxQGn8h6q6rIhFpc+Faf9
O2vXOJywY0WWuSTEWsCdSa9+cOT2TloDPE5aDGHbk/XYgHL/cdVv+/BCJQXZO2HdY0LumK/DAG9x
b6G6RipLv5ghTSwL7GmI7hQzbt0Wtkns+jwAySLcaRymKdIZQ8ZmgCfM9R5Rmq5qPy5tM1JN9mix
0Buf4xQmYsqCq7JTdVLqFbiBo7BvToZLBCCJbVrfWxIBusAuKPZe4vOc/WR2sxoMfTe3Dk6BpLiO
gGtghLY90eLALBoGUYULa4RB250L4/3rHNgm9eKPgR7uBvZeWgaw79nwXsP/g6nb7s2IbCPz8MZd
cNZLYEcpAqkg1m5YKBGgNhtsmIFmL241E9il1xUJzyJeBlJTiCOf8nr37xl9UYLVr2oD6m1z/7Pw
w8UeLu3ImvcPZZ5KkKNC7gcYaK9UA/QDFi7QUOiuv1D0P1ld628S9hb5Aui94lBRHC1OJYSzmO+R
HGZW3dhmssjeQa/UhZMGMGpBQiGbWBPjQZWpTFvcG3FkxzX7MKJFVp/g7UszmeqCIpP3LNdZBe4V
/pD4LKVnga8mmT/TH2pqob9m3RYtsP3duF9nxHrdXfmocqlXH4p/85POdeeZTBBKS+G1DdOOCTxX
OI9SCOE1dn8BMrmUmomQy84NKEns1act0vAXgcPsINH1Ig098IExu0TYlBsSWeAlC4wRSBd0rfUD
qL/QDES59F3fxHmEImTIy7//Tmk6GIaQmbFyqJyYQ3/dSeHDn9HdCPElp5vDHonpX3bpBSB0SCN7
HdzM0Iu8a+UXPVYOrUCeLVEtpy/l7NA0bFyhNJQ01IcgWvOCpKuMytbN2uu+AjdAuBId/rhzrYRz
VTnVVdmHwPTcJGp8/QiJ4HpPcdqmKPaRr5Q05MrDeRbW0HrHZtZaa225sShh6hYLJtqX16eYVooa
OAxvFqMoSXwGgh/d58kt3LDmtZLOsyGTWoQpLhHJma+BLfHIZ/Thtxhxf21XxnbXpT1DWxgpkYRy
6Et1cfS3XZ1kRQDFCOutvquxHkLq9M34ycW8W5ScqgRAsF7gamlzeW3vHv1ScP5QeJrXmCuCDH8C
Zm2aCpBVQmlT8IiUJ4z+jEsRTjCqXV//VkJblAXVMEOKW3ich0FF2o88EGJjUI50ZXrynUHN2EVM
FIwOYp8fD9hveQRiTXQcLqvd8aoAN2soQPlsmHa9fVJaiyDES4nhbTzYgt7XdmbrEzgMzs/uaPSk
CzDZy9H90jgdEq1fU7wx23osHetcoaSyH77lDd8Bj/1RVzi6cJ/5U60PGlQNUR5Wdppj0os+aAtT
dC/W7M0NGO2Z9ErvlkY1hO8OdF2vzXFKehFZQPS7X2xr9Y+PC6LhirQ4CgE2GXrdNQMDA66mxkk9
fEUne6zucZi/t32jF7mmQLITgTRjFMtfoJS5SgBV0jyJLJ+Vp4pkF//2N0K0u9OB8cM45Fo/rbZ8
3RW4pigK5FkUqiQwNImTH01FCC6I1Y2gZx/T/klTvQfJM1qtSrFxZXQX6+6sP8hEg17Nm7cYCB2J
CyEFF2ePIIzVh+d4YtRWxRZZ7fHHpqaOpKpGzjUdaVeIRCnwjLMbpr8NbvTTm/PPTEv6ynHH9m5o
/sm8K0L2QSIYXi5GbDdX/WTcxxPPHVEe4gGai/IMM87zRDjbvL9rYPBiGXvrOgDbvdLJMYP5Sn2e
AJYLFYOpaRCL6WZopUC4QYJO3u0sfrrdbNR1qN3WXtbf76NQOPRNhX3NG2d+XitM9RsKLeYwhxJs
1wJ51AfZOt4uiQfOmTKid4C7F4M++ZulISzW40UzlsuQBs3rh0uqMq1a+QaNjUAFZ5LEkbznbANY
JhOJETdRNPAMbzgVWrSj5fZeMJICvMQwAjo2gewp4ouHG0MT8g6DxBF7A8DCdANOtZGwZWEDly1w
2iiw5Slh1rvq9IJ6UAxoNiEMZuM2QFyTy51DjOuS4gudNVhXcqkrDDPBH6WTNvQkbPuNHOeXEUom
yycFrFeCYf8YBAQDTZsqa1iKqchX8YOla6sUMlvwi68ErImH9h2XnFHbq+C4S1tdfMyYy5fhdXVH
nmJicnKHkGd1hplpbq7lQmIRiMUGidDuiL3dbt6yxT9/6fjN/3kIYszHrIvREgU1pu8S/Zec9RAr
alcWniwuSMMNeX/uzbs6gf4KNAKqkjRN/E3Oh83RfII8vSEsHJDw30elncA15ZOKQsvw4uwwemjB
8B313YpPIIinjPHL+V8NhcUPL7b0rQzMHaBt+S4ie7ftAVovboS4zzY9U2v0mLaoWJ72XZMjVLDY
ruPVKXmU8aKcbtZkBOj3r0mPDFon3FlBx4L4aZ0wbJEaUxKAXe4oiujRoAn6BGFNdFeCmtnt4a0G
UIySFu6gd6RZ+NHeLftVuJ78NguKl1py6LkW/vNLbR07uLgDuQaZUgfWemi2sXicWH0Z5sJpGxtt
J/TmiPxtu4gNW37aqcgRxEAHeF5LrZxr2H9/xG+JA5679xicUdA5aU5EeldbX5ZKjEB9wp0FRFMd
Se8zozIdx3zUv9C2rmBPQOY+htS3/8Cbu8DifFV32Wg4PM3fSQgdxsk2wuXsYtiboxVHrbaVZXmW
fmwdUVLDrmQWatjpJvJsyJ32tOrltW9Zu8ysv6qWRA3mvbS6onxGd0hg2ZdE21okGgEVzu9NLmnR
loHKtSx8lUS+cdUh3NyeoyFHCsI9Qhhn4HvqJV4eE5mdhiVpxWrPYxzBnM9B9IEA/uSPurN+aynu
a/JgMUv+tljq2v9o7OjB9dyPdPEH5T0aLYyjJx2XzyvFBvOwUV4fq9ssGek67I+qcbqKm609KUqc
8A4V3uPkPIlRM4EKUfk/nK6E5tthuQXI8buKpF93k4AXsga6sJRXKax7h5p1CURMqzdPoeilYRjA
TA+CSTF+sYPiVnhybcrZkQWVQMGwRWldmF58ZGcenYeucA07vKvRUQjKt3jmUw0zoUZJr/YIbwOu
fnOiCVfzWY/fnsGtk4qvwWsEdtO6Kpqr0xF0bO7OnjOIaH9MApDgEjCzVsDs7DeAhhxOG+QjL0qe
UO8L5dOA7rdeIUcct1jIho70iTbL9mbIxRvjeldv6YowcqMN/Tjb246xJRn3Wy+rLbmuZK9TKdwu
GgTcrY1753jnHXISZNDP3w6VV+XQfbcxnrw5vcc36d/KHjz8MusR0eq/U9uK6Eqv8SgbNg6cIchR
+IPc0/jk4NaAMdqm+QX741/CBLH3CWLtcFFWrfRWJmWfyceIHcGwCtKWfHeIRLmohgOQ/ARyF4Ry
O2mgeMj1oaCZrFFwbCLqZbriVr35PhNkICXuSVTZQoXdprhShuMjZwCol3soeMt6lvBOFBATX1rT
Kh/wRyrivHNqj2QEOhBYRxx1rtaPiv0X5C9tlS383GpR94D2T53H1Kyk7Xo1WJ6qI1lhf1HmcinL
MS7rQK05kIpIJbFZWkV+Ifl+7602Yce9RhrMzkgqOc+bbCU7vEnVwOOMxsBgZXulz1ecqS5UPW5g
wnkj6yds11IU4PpFttCDAPCKI0eRV7RlqB5qJgZz8XSDLnOACYEcWRxNWgrgy14wUB0e/RXFM1sC
TwQnErU3tWxWYFiQNCX2p7v2IYO62Yo7xhbaSdMbc9bbMy5OZtgy4+OVEYPgoVGp6LPQWxPCIqTg
XMujbF8imI3nKZYb598/t/2/2oUmfshXyuOj+Obb0jf1UN70QsYwZi4Ct2n+UxTiIapBE5lMgKM+
ymnxxrPOOaFw5U8KQK1E9ba5U+IeITdTexuDqYV/AteR2mxm/Z68luu8mQIAIt3XTtImsIUimqI9
af1oexufFqOqAwwBYVbVFdg71wVy11zGdwgQx8n98bEqmBjZcUFD+73gtFdIECJKDb/bDGmzMibX
KFXWgJBF7R2kZVFLk6vmgGlCIkIeqoIUk+ZwN/RxLVzNwY2ueMSogI/CgQOMM3K4pkfL8BNuyHKH
Uqbgg8sgMpy3P/hpkLcNJCAinpIbMaD98jzbQEa7mpnnryrbPXM1SxU1qFtycHOqkdBLDJNlmjjb
ph+AOuHa6ZvJdASqVG0LyB3h8769EVrEH/ads3OB0LgQAMn7Bmw+mvM1FUZPfb17ymH1h/8HFzG5
wNN3NdrriJq929Z0bqB3XYbrggvp1b/e/a3Kq6AA3I8USYPRTyUE6/5U/bNr8Aoi+DVSMnyZNiEb
oLtrJPbLuzJL2dVOFFxM1swsMWsSdDCgceneWMNfsTKALYOazFCDAYWd455VBkyCv+YiP+IEP5qx
fA/jc61VPfpen6ZpJwkMOM5rBenDXE3DZsN63jlW7jSN6vF6RgPYxufW+udCg2jHsrbf9V1UZq+T
zwvZt2wqjPnqpTYEFJ0wHV7TW3xS1baeNxFDw8cYkiXJc8cFbJdbwUCW/E+wpBWPFZUuNqQLqUN7
g/k+3H+vOg4IJDlM1vrG+u89Lq0XbRwxFjCMHO7n7OLIDDy8p9cYnJ4kf6egGMc5sjM4uBCqEBpu
jvEVmW7LRtA8B+oM3gLpqkNsym3mUUwzJH3nqKZ/SyUWpIuaKC2GtaFU2MN0XK5avUrzX4esJ+mR
obFkZrRFzGNmHwGnOu/L5iK8CHR+bbI3IZQ/WMCOT3y03XU1GAtXzpF+RVUqjlnBJm5dMRS+k49+
XdrXfdXtDE+l24mAdlboCiq47+575ZFznoI+XtOxXbJ2clDVDQP92nbzjuzN1QJKhKeV1B//Eq9n
EdVGN/3jD4cwM7D44MzErHRDm1hZfzNmPPhr3R/coWDcZQYmlyAZlgvYMDkeQFTFxXheP3INrprr
kfYW4Pob+ec+bo4nAokBZWRhOM60J+hL9LU8iVDPvN8vZsfR9cIiMGFTUGcXy0p/CPFXy2V2Oap0
EpTmGUU97pEVVM9vuS/QT51RDbit7mgPPGSZepkaPk/GfF7NDREypYxEsv4C2EScka7oksQD8dxN
ibQWrrnspFT5tTWnpdJFZVsi8t15CkDbJVwoSU7X6EcSi1QKOGzqLT4eEo8BmC/DU+LbS/gwHQsE
C7UhP9syKA0HjucbaJhIH1lzW9sydqxivxkOxEI0GQtKU5DuNgxZQqibgh2e6jM6YsWZ0R2zcmRT
5xnIImOA7PEXHAUAZOkgIV6GD1rWWx9i5/UFKFArxGszR/FKfdIjzCYU7Z2MHFdCa+KcLgSy/+sF
/+WvsBqs9SFrAyslWbw7ApiBTz3aRNDdRjJvy3x9qYcH40X+RznBGhhjjBSB1moJGRB7q/6UCU3X
uhwiXw7H+fwZvOC3J85YayqV2ZHOrqgbcN32St89kAvzDhcMsMS3YPifMLe0JPAXenqGieYOO+OV
igCF141BMj18I7KpqSGcLhgfJywYpVFzLR+topoYshIkyDcS9BBARtRpGm0FEolLetj7prKPV4A2
U7SYXRSiEhNwD/AS95LoKc088VsXj7SQ39iATkcI6IRSv5he+M/IrlV39b656XYw+eNBiutb+AEV
2DQtHwf89ZuSn5xWw+aKAz5i3/ox3TYBhoqTD2V/GmqMJKKb/1gSNCAev+2Ss+jlRxBcu9kRARrk
ULgqyv4NN9uajgVTmqDVQP44PFyOGtMF5VopZPYAS1vAYVtsD50lLDbZGOfICPO7oesi1UDoFp0n
WAPEzdMcEVh4lDS2i3/G9a0temM+Bk3vo1fIq4sqZnFcJSrGtN9sWGP8663oFI5OXdC2lQofIXt1
IdmwC/XAaEKqPjWH3LMqYXqCT32Q5DZ0i27wQyvJwSyBLw/vkMW+/nNIzzZTduxmQHrt1yCBSDD8
AswYGtPTB6nQ3xy2T+cvf+tUxOQBdvdzdpauq1W6crQ35heO46hKa8qLpENke49Pwz+P3IUWwTT6
JByJLfY4F+cQ2DNNj/qUq/u1SfVKQ555Ajm8ovvPtSMjlgH4RfbRJtZl16Bhp5+olVPm7ozI0S0o
pZbhm1Dp47MjE9v8tm2ME7LmlZOSMA6TYfx47Uqu8If5npOxrAE//j1Z97r8yWapVozqvJjS6qKn
BVGApqoMVzlhr1CYTnmvr+D1epCe6kVRhot8omFjibJDz2TrviPVVZklEmPvSopOxl7hQLXfTeAD
PXSCCf2HOPhA8PxT4fM0UpWzD3i3OoWeV9jvFSjJ0W3CL+SVmETi73Zmzl5IDPkG5fUUeIjyVzQR
R0X7MynZ6A5szIhc0/pBHI0eOowyd7KVQkNi1yxCTKJY1NodrjxkPf+mvNJoc/v9HVVAg9sNtDHO
LqBSnIiZ7iq+zBdq9cvtI2teDuKVefZfr00x6wdtK9n+Wb3JxRayG1vBm50Go4TDeBxZZhchxSLG
OuKEkViNhtny0JOszc8zNkAcGO/9QwlWB3zcIPsLhrEsOvDzEcCL4cjyqdrOy6lChwD4GDhlsr3Y
ViN/2ng2mG/LULvEXdxQeWVDzzsHQtnAWUq0CwLHehplAJtWDdSGHjA6RN26biEjcbChU331GN6C
7tRDB11acGHIe8PKjf/Oc9DlBfEmX8SQWgXkIyXtrKFDexnVSkv/nTQph4ewqmWe+CyXsZl+RJhz
5eqG7tyCGbbHaHnRYAXxxk86qLbwNZG1cDF+GqkMIZ2u9zcM/VP/dmDzOgGI7T95zCnnyGMD1aSQ
3WWYulpn/2+kk7QMnC4ivVMAZWXy2RnFH5S0xs+QXjwpd+TsWUv3Uno51uC3tJToawXZrhb9qhye
uE3/8ZeFtK6Ec8tRj35iqqL9fe0raLlxfAyJESUbZx++khYkrIJ2FVJs0kjdJOAgZUt+LKJ5tDQ9
9kZpS08d7PcUQkN/WlR12Zdbzfl2XkEuVBcm3Mmf0e1LzUe97QJQ8ftpCN5mIP+O6PAqwCqbsYUe
t1tNPjNUhGwMhPgoIB6W2AscNAKZGV7FsoqqBXG0LkzXj4KR1dqiVhSejTP+aM1Va7NuoHk8wiB1
Y0tz8hC1bT16VAugl9wQ09YblF35oqqgFt4xaNAxTnVOOosweeP7LQd7eIH0ghE8RmARWNYUgxrc
BdNnHBzLv8rhPn2HzCxY5GTfXGuk/LXPcTf8+/W9RjHmnja2ktAxMl4AldCgsBWFu0cZvorW5/S3
c/XPPOOC51svGkc7Rlgz8MRIopM+tN24qxbJ5o7UxTrHi80RVznV5Mmm2RWdPHunJcLgzIDKPVYn
4+8QF0QPUGpXLXeM//kQaDuuKO4CFyXhObeQ66NluRtDLG0frVvLzREHEovzscXeLEzC9g8SO7T5
/pk1MCBut2OXbADRK/xDl1GqQB4DZAbaalq7KCCkyfwNXsqyvTSBxFHYSlBt3de64Y7OLVOzhM43
9eDY3R4dXOS/OvHzDPVgXOkcGMlnYF45awpgtlhLGZR1O+NEfMQ6JOxpz98p5zuvtO/eFz9g2MDj
n7vifHNlztix65EAuZar5tRkFnpxzBiwbbsdGuJqJaTgD5XiHhP4BYQ2Nl085JTXWmajKXeWZRFE
krYyAd/pJEP2tvGweF9j3laSQxYdQtPtPnY4r+a9gn+FyzySEmtuC3yrbnyRn6by9pSfQKVQ5/t3
kFTMSdrgySPD1PqtDs/dCnKKtLGxnzdHY9EbNhmkomp07c/TCRrQqYUfK5rij4pNVtpGBewgQnc9
i48zFH7QvPOMKKeRmxS1sXqHJSeUalyOdvVhL3lPo+4/SiOqJG0BKJ/xweBVVfTbkIzd5a4Kvt8n
tZQpvO7azM4HvR6TJP/sApuEr861ru3lqvA1YtweDALMtY+FWfxsw+u0ClrxWphLhU/cCbecidMU
wVUlnEZgQMcFai3l5glE/sVhcNYFEbQT4kycJgMpf5LG8CL0FI5jqa3ByQyLX9S0cNRskwcRrlHI
OuVNnIfvPBHZVl6Z41a8t2xh85KjkukTkNYFtR1w6OqZ4lYM/C2Kw3C9vT7mC8b17BIW2MVVSipT
h7UM6T7ug+/DxrPzHJ0DWUsUvNeFj0mGV6JJ31D+f05ypNFv6dAZt2Cfi3uwzO9C08GZ/NJ9UCnv
1kI6bZ9WARByyHI9LqZ4tg5zC7D/BGAnHWN4BwvLkbXyEOfYpEcsbIB0PhdkKhV+SVpDXO4OSxwM
5lIHzkUO9E7DnQXsUpWFJ+vrM3w+51ARPmjrXfu22a1frTW88NRQFrwL7zIlkg2nONLdNKEbemsl
2cJnnuZc8/jcAdlirRb9LFFp3lXHa2UF5csBKrqLSwovNJyfTGt5hYB1dX8CrKewUKJYmWdArSJB
cyEBAQtFltOhNMm5p1JyysbQt8QmQR+p6x3g/eIyQb8F4Au4NsVSwZPJoQPUQ0JAz5qpLP3FI9+u
q8wq7TGrvkxRyReCehgQ0lbT2dpMmH8+P0vYRfJiJsqPKBuod++lPPYjJgSDcmyz6lFzP6RFtJW6
arN7nsMj8avEZEn9wJ5RhH6vgU2KIGo7KnE7Fi1/dCtWu1CEq7V9CnP5vyun0twO0LyBfhUE+Zct
fMZgVYNKPZQBXsFiOiosrTpep7jpZlOed+p32ZPYvvmHOBDx72AdPApYgNGsN2fI8hEJbkuY2tKM
Idc3MvvVgPVy3wfDDYnsKSOsnUFxvjKkpRsBMy2C09uoLY7yH7/nVnX0jVz/TN/HcubugcLqurhX
kW5gb4ddKf6LjKOa2xuyvFCv7xEQoIKRiCsgLKHKUIpharWgtPa4SanTCSVQB92FdHpjHNCorOxp
qE7Q6JUuu7ZeaI+T7WQ3ZAKDdsdf/MEtxVTgSlW5moq5hSGLlxXP4/CxAz95tqh3JOQcpw1Uujh8
OJx/2UJyWX0bICtswoDC9MNP440UeG3xxxTRCLu+oTo8ByW8E8S1qtfBaiKkH80Bpxt7r9JzppVC
xa3Tz64jT3KkMv/fHK+WyCLMkbQ8RV2grhlnXfGZmuGFmHD3bpP4DrQwCBSnfhWbf/ai0m0wC2Av
x+RTztjuen0O3qz+bnO2fyppW1k5MbPhvHpitQDUDcLsDaB61f6XzA1qPLTqOe4uaO97GWgv0pcw
u7Lz3DnPETGx9KILp1fh3Us9kIyYMmlWROlAnEOqh6/FoIyLxvtDIYqXwKnmZ7wauq8BKElR/yXe
oyvSg1KgsxxpMH84gibUlQ8AyUOL0YStSTRt9bT3jey7uJWDbLkm73YNYlc5u5qI0R4iolrdHXye
IA0xYLa0gATD5Pa/qF+1sA9tCZdy5IudO3wjK52tFfvQbtgXTvd/ESyQU2Rz7MOoGXY8NDJIUy6i
XBut+O2IS5coqfYDSgr0G6OBjgxfmMuPh3MJp53elTRMgwZOCIQQxtlHsQGUa0ATlIOjggAvmcDg
Kp1Gv1bflc6ay+fCvXZo23E7EyJ+IV+gm3aX1oYOGUXpgNRvdahbJm+pPOUgesqq1p8AeXymPEtP
jieyCfH1udt8IArfZONiVdE5SgEWfEY+0j0o71LD6d+1HqGvjgfhSD1LUza7x53INlfZoZxgVsWi
h3iQ4gSqoQoJFmkjAMQNgGXq15mIEi/yuE5LQmcRHHzGcwb0d0WPMil50AluBq8e2DGK8gYZF2TA
u1PkdNAxwYnlT7fOjZtApUgxpxzBEvxXwbI9DGEQaRrLImfckgmYk2h5qvR0YWop6Op4KZQewIwB
LRSHmn7p0hZeWDYMmofTWUW80V+baFAl8pjBpYMy0MFw37NUc7L9Nv2X6oCW973iwQPl1uHH0Kb8
mu3CP/gEXjJ7KOpAOxR4Gt/FkSRtFfdv1a3n6n554QshR8n0HuZJrHJRvhVC6H0iW0V3sOg7rhMd
Si7reXpL0nYmXM8aiCh2mDLoVo32A3m8PeTZ/P68JsbF48tb+KWa7rJrV8PpdV6wi5ZDXBgffY1R
dUVgmgGyZ9dys4MQcb9cQQM4lNmcQspd8xEMaGIRf6v6jGdgUvOxlNUirZDVLrHxhUSnetreFMMI
BSH2Gj2mgnyY1dJpQD95IluJGkbcCJBtUEhV53Wc/Smgx3ScDXDgaUhN0ki7CjLattMa+LETLWaa
uBx0yVKbIJCMeiGhsFf4zvNGQHSZWwsYOB9eQ8ZPEQyAuSkummEWabrM4rKVDRcwFoFBC/vu5QNq
mEnGL3/pU/QCqeriy+4w6DW08/vItvb/YFamSj7HNoQMVP2puY5oKjCPiPUe9AsLQgIvYIyMVdlt
1acQ651mJrY6/BG9Der7Rmk2yvdxz524PVd1cYwZoMNfQATDowDNg04RXZZBvHhkCr7qvtYk3DQL
9m4R/zutEtNok+eAQ4qL/L62sRZlUjZWAuiMQyVNClhNmmVu576cxFU8rRMpRzkIiq3sUnrGH0fI
ZduLFDE/bOgcxdMf+YtKHvAoaYwJ69gtdUCoI6KYw9oZw9Zk4q085cIdoVWu5M5l3tksG2EiFuq+
4fIz17UM6iTsekgJ4q9dUKgcXL0WoxIyGb+n/jufa6CeIS1kIFwg1wkdBsqr9dqYtsjdknduELuk
NroEnrN1BRXX9aGKYvJouIci7IAN2Vpx6SdnfeGauFHYfVQA2jEhjD22V85WBfznGbwqD+zzcUQK
baNpb9QFvWRzBSXa1cNyeY5G32rGaU2pMF9LjfuIHtN2VRBLdBc0yWAVjL3HZPHpBH1/BluCDGOU
owFkCP3dlYbuXNZdONQdtS9gdr1cRfpnEEpwzWeGGnp+9muW3gcYRCZVln/ShP815H6OMOVtgoW5
/9iO/BAvlhT9xTcVdu+2kJ9x7P6mwyUa9YGlqpukcY7KxBiVcqojKzfTIf9oAQOZSHc8HM9/Iura
z/OEtujwVrsXZM6mgQbRkd72BTXQoNyvA2a1pFJGjQ4HCZ76hhpPvQK8UGn6AASh/rDuzH3XG23F
8L7JMxku3f1tKxdAvA1nKNbbr8BiWUyuwGGKQ0B5fE4KqSNZuREDAVYw4v8SL71p1g3aLM2TDIrY
0ISMm9Qyaxv7S5accKf/OSb/S7zoSqEil6adDqhCuwEv2THSOl/z24GEDLbLi6327XKFZjx1vsAH
c5nabe80J/RwByG9Cifa1qiuvPtTKSil9c38ICHN5/Mm3MOAgyBmDqLrllMJRfDXB1WTUgjmg+PD
o38aEI95Wjq7OnvCxIywFatx/oRgy7Lxf1La/F2MdOh5crlRrbfOpM/SfjtEuBZhvQ9y+Xbn6oxy
QApS2C8pQJM8eQ/FhaDg9JYgojv5bYu/PYQqdBnVITYCGFYd4rZZlGsTNeYwf3BMzjMwjEeAD9/O
RqyCOfb+5Ccv4kwM75AEq+TKjAi7M4KiWmVa+UxClcgsN/9rWcHkyUrTLUQ9xibWbyxY9Iox+WOT
57ZRuasdqLYQy/c4bkLpVPCaJedkzEfdlzqzy0NHDkC22JnJKf7J3prE0NaL6ZsuET8wdz3MHwVa
po1Q337SLc2+YQWlv/Q6cvN5r+n92osGOIYApxbRCr29bQGoccbUx3MzVGBea3WBEOkh41in20g7
EOu1eh0CX0AMfdkCr+cpGzG96d9AuHVI7cbM9q4TC4boBESl2b+hFlU9d+UbLg1DsbvFFYn57zMu
n8qBHYVt2Ym/twG7u/Le9iLhN5ByjY9oQw0qnECo9XbmGh5ug+i06rUhVULgi2307kZTYBiFdNNY
ZNfvGtzVI9bXxAvYl8x5aZiVD2yzxiYKXXGMu8XrMQu4yZNMKUdrOLWh6umQXzOQXjBMNacWe7T/
eWyObPc+tMI6khTn12GVRgOaLn/nuVwdRox2n9NyJ5snc0YUa48cNvh/Iwf4NvNnjWLVeGWP6nj0
pFE9mBi0/qNZqsGtNmC4dmQr0/5IapLOhoGisG5bdIVGbNy0b+cmyY6aGww4BLMtWr+fEHLGCjvO
TinxV05Pi1zinGcS1ECSQXnosNvCWVTCJO/0LCT3qtBXgwzpJMkFSqx5xyk0VIIQIIhDuL8YLq4T
ZL4f/115z+wwPgScc++P8KsaldnMGUC7hQlHJD4ZavEOnN/wiP4vxaCWvbcp55HhJq1JJ57jHspN
8IwJYjGPW/vpbalp3uYyAvPBssxH0x2Kn7JotlNZKn8VB05p5DYPNlqzNYuWYFRYS3aXqIpSCeZi
Ek/Pj5RhvrWfaZHcdei6pWtNTmCdblM3oFH5H42gGHITnOvRLnV6LUbrv9e0jDq5412ZWfeyY0Yx
9oZgtwcKDwIQtZFS/NFAospXQEp98ruBCTiVY+T3JPby4pzHZrqSqpDp9FoONT9oVhUrNorzQbNJ
q3CUxV/k7VkXa26Z3GXaxCH+JY5pEsTaEOG6/ROcyONyqnvrTSQ7jT3ZVv0iXjBdevfs8GoGnOzy
1ptaJwx/UM2sUFw3C/ck+1Vl+NOM11uAlrCnsvlerw6ayRKaxigYNyVQZq/gA3INL301kAOC3CsO
3/ijdA68gWzFxl4lcfu4LxKQyvmDqsZSZZL4iMW9OXcsNoYAXmsozypX6K0Q5Nm5Dq4M3AFnOmhO
Q8kO3hpa9BlRrzbi/lFnqVVbWiVc9svi/KQjxIY/bI+piuT6KwVdtZ07kT/A5mu5wtcZ9sgNO97N
tUHU8DqaGzGE7KuM0ppMxS6ixlTj8UO+rMY8tUMcEtV4FM+m1NnNdkC82MA9XOHyfnopHTqb/AVZ
bduesbzHEeMhhzE3tn8jKf6HGz3LdBRA8gLEAZ850abysRdxoIahyYR1q7MHXmmXStfsG87+8oeY
eZtEyFLgi5AtQAMlPtCltuy9rOq8CnqsIvEGH4wpKkipVjOxnWxbZw3rEIBvRabfZRPvSK7DlNSV
PYThdJhQLiRIkCnpClshLIkZK0QxdAuvKZpEuYcO5G/NAcWdz8u4V59SF6yaw074V/3TFvuOXQNG
uLHsNtb5rz3JDghszvbRvDffnbDdwfZh6RTezkduk+z/fP88IlmGNPR+9mPlxMU1jRwhuzjmKt6e
PsEAHGJEAzM5aIIOzka/QRVaULssfpNAs2rtcAz7jB2sTHSwTBzWleZ4Ic18g1JCQS8+NagAfj27
AN8Omewo3w8cZcKmA3DDUPTzBpERI7mrX2R2UxUA1QQSrt9sPZun7QCNpeunnDvUTR5XE9MTnuEa
mnM6p55OVgXFcRvsrs4nVbDddW+Z+uiduBY2cQv/l+uTJnJBP/dVe5CgPv1jbEqp1raDQcBM/lwY
yl7IYJvOTmsHNSULK280QKCvw9HtZAD0CZOKSigTPbZOflFAiLVlS05Fqj/VtitMJAWM9+yITTn6
JEoJuCWqmDfqMhJxcH5I3AJVGCCwyjLw51B3T5zYtltdWL8yhkEDW1SLsBh7WsSvt4IMwVZvySyu
o4u0M6WzbdCLJBhw05mPXQsNW5U+2nPlvu+Qigadq9wKoyHwbpeyaikR654JAwAK3UefH0EqLHxU
clt4X4PZM5GE22CahurmTDZaRk9XEWBKzbIBzc4THsj5/4o4lgbn3yOUC456q3a4SJDxNf/oK6RN
okN5Ub1V/5KVACBJrT72Ti0HWKj5P1MZwWYH+gH8HILY3+7izgVAuvbUX1DRi5yHFD2SuWQtd1g7
ReNSszGl9Ry7WTJ8ujIiRHSPRTdUWP0oKiXn0ZNh/Tff8xVBgIaiAcI1GrADPo1mcINYik5Cs5oO
ne6bQT3aSezrczAsktPrGDZzT93/QoSgXluOgyBtLkAqdiNsC4BpSp7TBnejs+k6dai6ME0oypF/
y+elxZdklLtmsfIoZQPqOPV+7feRfhQIle9/FEk2YchfM0Xff+TrEHPBkmy28OxPqxNFHHzqDzxj
0y2CyPCqVw739BMUZDa7FuLPs57pKo61hHACnA8kaanmCLOlKIHHerXPE96pqOESuRgu8CaIx2OB
GRlkhLIVJZXrJl11PAscPD7BwSM5Hjn2oTXomczlS14oLLRsyfRkdIMI3dEnxkKBBKekb9r8uJoL
jxPyxHj2YqTTCcebppTJVuG+V0Are6/iHb1+9eA+ksE6j7LulRYGuOCOa4dshnKn8OzCKuG3Sv55
9DSCDz0IW4P7R0jhywSu7ik90FK6etmDAvFxUJX88v+3Sb0uRr25xx0EXagqA9ba95N6j+M6/mb+
2tnicoj2mAezmqbX9BcIfUPXOHRvlIDDK3s25TIffYJK05gtGkP3OG45HS7fwTI6wZSTbg59JGVl
yAjhHpOjKo5kn2f0vkK5w2Fcw++4ZT3kDW8TZF1Si2xZTEIdq5TQ5qi5OoDfO0k18/KgRFrD84y9
FZOFuMX2iyC4ITuGn7s30TxqnXFshVwWcer7zTrEPsYjc2pzmLsswwixSHb9CUYHqi8gpV3GJ33v
e4ZBz3folDDNMphMr+3wVbqehJcUnbrc6eNq8IqYVzOkFTq1s0bQfnW6IN0Q1LnvNG7RnEheayOb
XFN55i/qFrN3V1PmHwf6EVxTEzFbAwwbELwBag1qe2eU75s/jip8x4C4ojZE2kYR1oJs0ldcXvEw
s7rdkGafskJxrCpc1DiVJXvICE21Cwg49MYUI73cgmtFAbjGFbHZO3cXbv1xCwuXdmvD3NKq60Yy
zxVdx54iwZMGg7SkkSC1jvgOTPnk2g0eHzSuarkH8oYc0OnXJMrYTWI3WhEAIxpOTgMIO2Af6jeZ
4iciY+XY5x0zpvKVQmA/beChct8OEgbRw8+7aMwNVA/p2QVPONVREshmopmqgUWNJ0K7PtlSMfG/
zuWEOf5rFPKXHfzQrreZ1evOnahwGW0364xCtu7AcxrfyyZntvjO0vrdMYFyhPLjWuRXPWlyuHhg
VkgnOHQF2xeapmdSnCQ0APXzD3WilY3wEzMS1+G5v195pnCsGR1qgReeDXfpBEXOuma3zzy9bGqU
5kCQ2Wn4MH79uIMon5ssU4G1M8zi9017ATVBT7yL0UnYpmVlodQHb6lkVhmKNeaDLWJ8E7bM12HY
UMP9vokzLm917TZiW86DWC20RHu19OqRMq9i2LDcfr+DdgHVI0TuwHT7CrW17/xlSWx/RBvXynKC
fqClg7bb9I5moUl+0v34tApQhBScOebO22YKD+1nyr16JbYw5B1I7rmyiuVlZMoMx7E8uovMwldH
55a4Po4YDfjnUMrPqsG7NfnbgfptBpG6yv89imDBFJrG22DoKRosSZm7nRBB6M6wDsPOTyP8qL96
PZ/5q5maov0c61RdSnuAunfUSMAFLAX33SDVh0W2rh6X7X54G9ypbZtjKmVUU5vrvOJTiD16UFBW
pXVPoL2vQ11WYtDUmYQNXhsug++/tTraJG//c5qA7+QnFBIJ6R+UxYmdN0Wdiu4lfm2vZxysqaTy
K2jYH3ZlGLHng6iTLvom8/V5n595tsBFnoKTJDfe1Y8WibQoxnM+jNTISZAxEA8VHHwX9s20dW2O
T+WSNsLRvsPsd8ulPEpPppYZchYNUUhrc0HfQXBFtzZCDIQBaBxE0sT4NEuHUHRZuIdlhaUEv81P
2RGE09flCI0rpUb8o/2el9VHC/T8TBz0YjpB3VJg0luoj3q5yc1Eed11cA6mxfJipxiRX0vY84e1
Np2lOh6kZN8mk01MjieJ6h5/UkcrULjg+F0uAj2gAUqY1dxOHQCaFaEPjkjsh/6hJBRniJx4twEt
L8vRhW0cpM9wX1axitpn3TLROiGsKlMO2CF1eHBEGadIXE+Fzy74hFzwe4hWHhO+c7QGe+8huO2Z
11eu9kLsh83y4UUHwD2sXydX6Ae4oN9KXJo2ZPXgb3VrlnZ3F6eGsUKSrWyLgjIUJRa5tgy/sPI2
jBmtwl6JQkc40fb1Q5nhuz4VBGuqw5A8VXcxc9YZ0TOY8UT+5KFEWz9+rPbtcvJ1GMx9xlyBOSnx
sJQoMpDgLa1in4NUd94nVITHyTlA08jV8GobXTrxQY8T/mvGd3f2//9EAucDJGtPLnNn3WEqxP4R
tK1bAKVFKZykhCyOG/b7XFRgeEQcv8tocpNC2GKp1HLSw/4RwGfLfKmsyAx0jOlAt1xFUoHBtvzD
5bUecNFz4RzkFx5utMbjpEF5VvhHhRHjJ5gsrHVvyA4aY/RVnZ/4yb2RIhA5z2iE6y3sQEZWkbvA
yckN39LTHNXyievU5Ra55p6IdibhjPLZgMN5JOEX9uYxR/5zy5ak9sd2r0A/xrum6d+XUhSDiwJy
U+NxfesNVKHRqiN2U0TD+rj34mDI4gJvKRXuEPZOFJSpfLqTMToGtt1e3RjRURaqETeTMBkrJO3o
3K7hODftKy//rd66z734CId0xEJ0SJQNZCmQIXXEVmbN5TKAQuCFjzB2G05HfosYuVfaWOLm1VEb
ZmqbGVZ3Btns5E4KlhJyC8EyzWntpmCxpftptG7TPZn9XxYshR2t3WA5cADIVK87dJJSE/61uRw3
Z9af4QdTNkVQ1q3GHbWaWN1/eMxP0NgLMXabaU5C0hLs4g2yLJ8ZeaJ56exYGNb2Ym+aHu3iVJjz
2jdOJYuldg0kZ8rmAC3671lDm4TX0h7Oyv6JpUMEUTyE0D0RW9b/S04uYRq3f4wUYfuXBre8HjJj
GvD7j9nelg6uIPzOos1yRvd+b6kMqcu/EQo1mc2jZe8xMUg7I/0KDJJ5jJjUkd3Zwc820GkCjDz2
3X1VQJyHiBmAI4SMVSSgz+JbXypV9dRh43tS0Z61ITVOoqacMJ1sqeqNwVa91dUdjQvHrXvUctcR
zyexaSCq+oDL0TRXh7OW55lQh3k7sP3nMExyku5FTnfa3IaZ/hJb/WCZULDMNncxMQy8MxZTzjIO
piNW4aKdiYqoJPGnu8i+3p8zSmVM4HgJ/a0NVnW5sDKBz7dTDMRefUFF8DykXGBIOT3P1GR4xoOs
zqWPbvTZBT4knuQw8i2PtxI0mPB+ALsdexcimS861rWVGPlsYY9PGWCOEf2dBKAz6xTBjBB2/6oR
GQynSNsLTLylqrR8rUf8U9zH7Q4oMp3k6uU1LAwstzm2wZVbMUWQbtWi0RG08uit7THL9Yewwnyf
faakG/xjoD5qJE/39XxeBzuhgxajz1le++msYYYMUgAORgQRYvV7GaBo+2yj6Dy4A0v4fnn2YQOq
BtBuIxioD2/O1C6ywy8Hpf/nqkT6vXaZMvUGEITqh8VwPzmKdJVIowdvvlGHBLUzJQGCs+uDEbGL
OaCu0k03p1rZ2fmzjQR1Cmq9zTeznM5gPzCP2y7t167+WLXNnmZN32CCxJPEnfnk5Iisdbfv5dI/
gxT7e5Ywd6Tbpmg0nE3C0aEAgRyND5ep/0niN/hy/3GsJTPlgayus4FS0ugISYeR1xJ7u1TDXsGf
l9PnIzrszv2Ry0Cu/jCtxeBmYtGwdnebUIei6/bPN1p50xJP8Qs7gXFH6j6VlGuFnK3mgo5ILQ0L
xobWKVIJFuYXLRsMKmAN61wtyOyuA+pVfbqX0ocGgfEkAkvhxcbTlNlT9X0rjTDSi0mA1p9DUf/6
W4djo0ujlM0XHVuECYUp5IJZoPDZTaJQ0P5YDLAJ390A0DqMWVL0yO2/UwSA+J4urJlThb/jrTDS
PyAyBJR3k4o5RLnK3wt3BrKBBBff5cDU8QiREWEh+OYORQwRNI5taWlydD8OK2GB6gnw9YQgjJeM
a16KqVw6HqSJCF2KWS2bPIDnesUfuk5X8qqVYJZKE0tvNW03O9n1srm/4tj06RqCN6pWaW2a94xS
P0RcV/nEymtJNBss3sd0hoFx3ca/h3MPlBlak6AakV6Ef7XlZDYaOAIybHVkJnoRFskC2dctTbF9
MPEqYUFooy2HykyqlLHTOX+pUHR9LCxs2hjZakc60u0vuNMCBCS5Y2RxZQacmUWmyWyrWU8qV+rA
ysMpQJ3/Byv6PWQjFqxtl1FUkd+bam0DX2EsYolGLwZ297A8ZgdQI6Bz188eQxi0dAxqs6rclMGk
lCjiD+P1qAe/NwnzBJnZIGB7JU/265HIOBXCJP0k+e67RRL5loCNIA3+iN3w5L6eLCKemVQLTeQV
zKIbnwpLbkFWp4L7l/q3wglS5ruQvFHhugxE/qWyKrxCVhp4NC2720Wmv0U2pPTQ/gUQvRDFEwox
sdkwtBTH83fEENUOIdwz2Wf1K9nq0vkz9WQtVPiaATQ5dMjpZzODVWs5rKrpn55OXpLE9W32VHzW
Q235KX9GqsIVBF94tJ7YsiSBhkY/1QyJjeasg11O5/z2UhFWqhptR1pS0D3o97eAQ1hBBsEbQl/H
WS+EcKmP56L5arI2bhdgAjOvqzDLpykl2Lq7DW+QeF2Lvpugrd0wnkzcN9YDmR+6Rrx18LBydYpj
+Jo+pgEAKKGhXqurnbq3Ioy6btd75/eVwEOjKodTAAhttMxqcOpfGcCRTk2ru4MxFOQdjYEF4KC3
9Zn7i/6V8dVAIjtC58pzkdTh6Y90+xnoT7wT9RoZ7XI/YdLneOffxwt+pYDk13L3JpJhjyeVzBPL
FWidVLXTuiyAM/Mk6r0+uvTBLTSWLpMUlKGpnzn27unTzzBOJKzDp+PUdE2ElmizLcKro3do9xiF
WYzPCPz3qr+/tbDU/LY44Qfz/fUf19vaqNOH0Ni9EGk+vgGNj+VWSi36i/GI4BZ+KfZo1uofTE2Q
A6t9twzX6f9sYLN2ipIvdcRgfeMN3RE1xnZdvRoEEZmOyiLSvPxXlB+yZEKrLYB+bLJVf/ZON/6Z
fpoBUzTTf1GSPEZVJ7jw4VIcBrFccP3uVOVt1VaDuBOGefQQlGrCEq1spX7JKkAE3uXjPfuSUcvL
W6STwMPMR1MLykIq5RM0oTdEbMSGCDZwjxnU5AuG6eEWr4NljpK4aUuYYLjShsoJe4Ya090Jw860
OrjxMe1CUo9zqQE/zsH1U780LDDmb0OXGSPgNl2ayxGzQZh9tcYXQIGeKibnnuNS+H4bjJHsfeO0
E8a1Tj2Kx921px9LkRJa4fbzMZvcCfCRFNhdjAVZ9L43TXo4Ynz5lYzw42l68V6b+jTaNa2kYlSp
ih4AkEVzJSts0yvgwEVOS4Wp2G58plSs7lLVuPVxjq3GNjEXEuVggvH4pixx1sYQ+n/eWU7CgOaC
Mg9+s08kZIpN+9R+3+BGEkgmb3dLYa//bdD7Vs9TtgvS66YOLOXg+PPidBwHaLfPm2fPFUrLyLT3
nNjwNy91dUrXbTvlMVKsxDCi8TMG326rXvkipXXgiqbaEgAXljXSxuLGE73cO/hUKpB9axpNO/ZM
loLPeET+RJlzxAbQaSNALYf8LyKZj8X72MtH6F2CNRrjHSRdWPeoh4yFa4SpheVGcx2AlyIJaNDh
BjkJS/0QQNrr0G+SBsZgbPO4toez3MgIwGMtMo+TJl2OBNNQ/c4xmjB9EEihqGSZxBpIY6qEX7XZ
4RDOge5yQnFY6jdpdw+q85yfe3+FyOeRlI29qE7ZUivy4InUvrlyyBPp/+vu0QGcbZp6r62F83zE
XHP80fQnb2lJG2uYXVH+H/KbtBg2VCoahkAFi0zhcVDc6X7+JnMBbCxVbCVUj98xpK/It/oklqvr
pU+RHWXa6x6G7vlwJL02YkPRPJoU7ZEie/mPPW4RdMHLBjEL8zPQ26lZ24GN3zWjN7j3xRDdFaxN
i3IWtdP8yFjILdrPqjspmrRkd4AXNbq+3M7UxnSFegBvo+GzsKSrwrU1JrHbdz05BGjKSKK8ci6s
9R6IZso+iWiPXIt29BQDcKn/5TK0ngeHok/r2MMkLGZmj2fxA+oNkwLfMunW21xI8nmsNbP6UciU
UczqR9AFFG/1Rn3jeTp5Sa1Mx7LyRQKeIQ2n/7+J4DSlAFostr9t12kD0uLkXPOcRs5ESQxrBHxX
GqYtLTtgs3kdG2WkmXWKzIjgUA/syXKvlnG+QWxpTEA+7gdXseg4c93YWqJvHeFLOcvA40PQ0SsC
W6BVpeZwRH0CJjTj2sSjnQ0eePz5aldAB6FnyV8a1oL3BEt6RlMHQtn2xAAykNDd4DVGtwoTIVfh
5t04zkZXBgTw2AoySwq2Tfc8StekudERVyU+BU5DbxJ53tD9SvJFsnf4tI24xJ0mnFoIM76D+bLR
xD8Wu7lSifcPrnb52MdAliUL9KGKeYzLzwybxesGlMk0rjViKJ7aAhYtDyiODTD1+SfoBlb59N29
WqF2SgZvD9LsuMGG+8gt2/k7/o4YJJUvt29SRFdPpK4ekAWcLPPiQBSBbqanVQNw5vF0yhgFHPFA
wefAEwxFEfFJ7kw9K/Z70j+jSrLeHTPKsN5yuAvq3IYEMU0QLMZ72dH6oLRBLxLmE3wNJFSVOdpW
FLncFg82Wb0Na2PmC+waK4xhk7uv9i4o5dH3FFtxD86ciePW8W3DdkO0+9ZCZIpiH1SQpyVt/xW6
PbxKqa31MxH37Pj3duYvOOTGKdmvWfxfGbwo9cuT08dVR5+HcsgQoCqKxJzM94LXaocpJwx6Qv+X
fGI0C6dAuiHRuflqcYi0Xji3TCjpuFFeacZvYNtcz6kT00MabMB5dhbdeunGYH8kXtiguqhq+23V
4GmVEForQ39BOqoh1xt2XMAs85XL7a2LosUVd7NQ7WxehqAoRhyio+c++ATx+OCp6du51lF50m0w
INGiJz2Ti++cu8hHP/QM7yDMI/wQDLHc9Gs7BwEWSycbWC0syDOfAxRKGhw6yQ9TODSnDa3gx2Xy
CtIsOaW8SJhmkVn9ZyNNQzrSEBY58ns8x1Kc6nN9JaEWb44u1c4au9hsr1kEIaoOkSHpJV4RC9sK
KIxzTVH8BgrZoGk/MOjoj/SSGhZ6Z5QOxcXj3eLY0XhQDIQgYWOAlh2+dYm/ldW49C5R9a7SwKn6
cMTjKhv2oAIiBhUDmv0VYUuTeewNMY5+xp28Qv6/Vs+zAmJ8gkIsD81NirIVQWvKySHXRNblX2t9
EnBRr0v5N7QVgcAuw0Fc7cm8X2KUhvwvcK4QHrGQDUT1pSxeiEN29k+2VnYL97RGmpVBDeV/Qyx5
FPkSMyTEUvqX6uOxOgSsxI45QvFzcPQQoH50faB4B1Vf6D62ptez4Wj1QliM3SFNDpt0VpcTpshx
H+qTyy+vXPIelrjPQQMyMuHSxwcF41E05hguwyHdY9I5avBXRTdU3KQP00KKDeBsVzkNpDFrErCt
NflXm1hRrYAWnxu9xnqmJHZtJCi5ECQ6kJnQOtADjcLhd8Kg88oBzTHcByXIU+opmlxdsJkcIVBu
eHGJDsGIPafDGG8MTYtUEBHKV5/nm3hi2mwbRcJFVlHrshSfYaF5uE8BVQFcMuyEF/TFcuDW9gUL
erayPzt5xaewjVqLi/fZcxOsxE0d/JVlV56ltPjA91ggiAN1QVTUYR9I1nmIYf783K7TriEGJa9N
dik4b7ixHvDrEER2hpwRCyWLAppzToYh9HKwEBNAq0PbxStP1cKpeGq85ObSEC5/UOA6xzGHQgZt
EWXaMcF1pT4A1QHZzL6lETzMu70aJOFF8FEzwD+RqfQsGAq2NKoiTlld2EUtjvDT1VSv9NTzeSE2
1iOxGcr6TXI6pM4gPhrfgw0Upb765RrDiiCXTgOvpZdjb8T3z1TnXtQlVQBziePlmmZCatvAY3bL
6rQE7yzkHPMbC0OsfiUnQXkELPqhQtLBXWC3dOW1ac9o/D+4KTf5XGHUpgrhUHM3IryjgYgCQT6x
b1PMaEjnQqcrFoRT8BzJTeTtk3Pl/vi7BkuXwbtCnOS6jANBXD1BbMTYNxDcbd3s/kwRmFp30sNF
KK4/7Gqcf/Qh6NRLQkK3f05IkaNO7Li4mGUA2YwIVY7eldKVC/IdDTYEnAu39XeSocJIYao0wGm3
A9J9eB1vs4s0JyEmG4ABkV6cH6MXPKs7g30HnmG+XkUyFmgYB18dXLEU6WKhc4tOZaCR5nyzBGsx
GdT1WNy3HScSvE+hKqdTod8kpZdUu5j+Rz/Ap78JlAmNlMlQV1SDOOq6YT7Ub8ChEXoY++ftKi33
Db//w6H83jKy1H0n6453LUKwB6BugQCS2Bx4AHKwC/+A4kDHhbInWE3Efzoq+KKqDhRfuor1NK8/
r4pgI92yLSwrx49RDVhWAHsKT6/jEdaNpIrkEBgpH4Kh2FPdxjkfBfETLRjkO5PxrqHHOchf1Ds/
32isLEYGIGhKl8u42o6Tpy7v4GPUrbtCmE2WTzXh7g3qC4RDcleLqs/sfgugPxhYp3wdpk8y0Q4X
MBc+7Vc4UAUG7yj3DiWCP/Wk0EYzfnu99rKtGajsKrEahENv6TbQEQgZCH8mNHTrgTpGQ/dATV5g
+OWpkETaVkH9SbbPnR1rKWNfjiTvAGflb2Zygmm5VtMxdk9Rq72son8LAbl0fUiZzZPyA6+ujPcL
QT1KxGhel5NmOm03UOA8AW3V6VRUq82C13jYkXm7/wqA0UHWIULHfuOZLAOpZfiXD+e1TYudRY8u
VMF3dJLtEedfyAI3vB0p2r3LpuajuSw44s+n83HweKCZfhUW6ijcLDTF66gUREUNub9REu1Yi5sV
fGhoGa0AlG15q+rW7lTLv1fS7YGDkWJ0ZFMelQPhrHrsL0XkCNmHiesOj2005i1h8eeS7QgTBcK8
c2IkceT5b4XML94UNdngSJ2q79d1zGUiEhDwmjZ+qdThOV82njVehnOXwqhvhSGyAcXuB5N7Y7wI
l2qZESKIvG8jtVVHib8OaklswzBKNJa0kJxhPTrGG3K4He7LF47JapXdZC8cphuNAT7YvlTe9gdy
PFJar9yc8YuRHK5XjE0BnzAqOtELtin9F4P7qemLd6QDhCdz4qWGYbBr13DH56pDdUCdKyGCSlok
EAL0yQfp9Kq6gM9QO1JK9ryRYghTSlrc3ElxRk5YGUTtMiJfM0Km6s5s3aPSpov04L10vMA1de1/
YYAmk4FOt44qba3rEA+UXkRD4K7s02ERrqZbK9mB5kidUB6O4Qgb13YPqeNiNBPNvaqodaSTJYO2
e1mBrISDX/+n2KEcekbWZU9HED0Vk6dv3Dplh4Z2xmlF8HjfqhLM7e+U2J64sv4c4MdkRgPqWG9Z
6ODEyM4M+YFy8QXqgeGCh1HpK2yF+Cy1SEprxdG4KM8LKjGdnxRZIohv0GJYCD8n6V1l584gBSw/
bkZpE9u0IaCawcetPIudZKdWnczpjaO0VnR2ZLhMEOpJOFYmYzGKdpauVJdbdUwxqry9MS1WB7rZ
muayHDGW0UeNGfYNdAR/7W7RQvvE1fK6ZONFY53Oy9Mey3CAHIxz490v+o/idTnDR++y1NMXdoGZ
84E39pJYueAywwMkepZ/NLaNbeKf3VQSBt7B4WK32S1P6HBSYiwAiu2T0RlBo+vYodHKbEuR+9Re
NniCDXDpFnLp3RBkupGRW8o8hmNnaPKAsyddQAqUFGomXjoEoHyDkT7aucROKKgFi96sEvme5xxn
RK0Owh6PkHW1jCeLpAxi3pOF/4O6tqdRVkbeGVFo/nmNgeF1BXIpkumBGnXiLlKOZoJjE2rSfi59
lvEERNeNzQ1c8ihkc0NVlTKXwgYA7QHmfJX4iBiQ4Tq7dcMflAZsJdsK1Z0736EAn9nOtjOVB5N0
kpZQ9E8sQTMvl39d+fjZaByCSB5MPgnScDbbdyHdpy3svpX1qb9aqUCF9Vul6LJzWLQhrUjufjPy
m+tgbVsNuEzglNdoEKZEQFcEQokRAr8XSNNdMu1WWmIgrVPetC8IfsayOPW9IQtJW0wbaM4cb1xK
CH32QwVjQXbvR2hOPun7PW0094WJzSxCMyfomwtlmMRW9aMW7oiR9OvV8lTp1dWo3m3IzdUcNxMf
ZmWfWdjl+9BolnnyjBETzrPLO2SoOef8gdBuB1QQZ60UuYmaToUgNs6OCZEgc2NLEjvECUOIOWrV
4JubiAhIIPzN+xzfvmpyPIrwqnt2u7ch0I+CdSDk4PvIlgo/91VvgBAJa7Esv4lxKXzrXBhGktUy
M0p7qDG2HeX93QhNmo7zBZhWvkqfIKmWOP+JjYSvHf8rew4gVfoB823APRY1QuvcWpTnJpk3nsj0
gxjmIpQvrbuHz2i6vTu5OM22V5/RCTxyb8/SOIKG5wHpGI187ezEZ5CKTNhUIHOzdAsufxaeHHuG
BBtfdCs5GYp1ags7Cwke4mVH1kBub2u3FWJ7bxTU7FRr8nCmmnNYVF6ih9akmwx+nfyg/9W0Ar0M
fqfHfILxb1EcgM7bBq4tANy80n2RaI7fT1OItt1TgUU5UZF4NRwMud0vYwfD+DAm32N3U+LfXi64
gv8g4qPJpTv10/WBVXCapVcCmOdwNcSCm2lfCBcLOewVxsuszxq+xmAO2iwDLm9Hs5ecFDpVHRds
aHjsUu540pm5g6XWm4sJltqm2QgxYn+Lp9Rkk5G8KNStc/JNnwZg5Q7716Ce28Bez7AsW1Do1VUn
Ve1HLmFvSIEQNvMcxjKMyAJLyn1Jdoim0RRMhG9dY17NPV6fV1GoSeM7SRW9xlDXDVhxnELHUI+I
2Mr8R8abzjHfD2/U+6LtuSjLuSyCChVnZlrGg4/XevSoGIV2xpnTg44w6snOkUAwgXDx7R9RoYnB
eeop2muPnEhePpjse8ktV3zYRdd1P3/Q+UWbsqyQIFJ3i7xI6wKSK7e0pPqop+yUAi79uco+6AoC
y6vFFwL8YRyUPqAud+2bjN3LzirhG0TY/9DuJEPFIv+dagJ8zG/lGWAfgqYBFU2uxnDO/98MbQXx
HH7zFKo9lXJn9omVuym+/VjOpo3A9AL4hyeKFz53kJqzc9RyMNyfMy9I1pSjQQaxaWqgvsynbOvA
0WgdTpA1PWz5gaYFdFPTipIy/SIZ4HoMgHUpyzKY0kY/JO9uqmBPofHEUBcqUfOXt/PqWhXT2Cp2
hDMsjBAJ09tBMwPMPiXn1bWHIvs8UXzLKL4iMn4d7V29eQFKsl693mIUKO3bqxFtywpC3VLKMono
Bmh1RlccDKvc4td2rtO2zwx0FkT8qbpdbsX7B6Tm2mCqXgfet2cwxrErKADmh7HXJofsEJggtdu7
wLgYGtYfJwgffCJ1sAtizP6zfeXUj3wqcVrlfeWH21YpOeiEivMW+HxeAfihRtFoUMePamgmuXDL
3RVTwKjokkI0827BOAfPvmaqcclLUnX/TpiUEmpM4VkDCRZDxu/Y2xQoLKmoD7ZuMeDbT8923esH
adjNWzxKKljHW1hAlehnVH60xWU9rjPrtCnk0yBoViaMweA6WO3uAerE0NLktWVBUwp6uWzPAQEP
pWB9Nd1W/vCejg033oh8ajRJoeNJUCPk521/BO8GBl+N6snr5N45UW0oELQhsJSc+TlulOoQWUVA
twL87rrm6B4YvSZwd0yHFyliiTVD92hc+7xgVYjOAK33TirLe1mJLWOgXfYnXZdEcfmu9o4f3Bs0
4AAstAqBpbBnhI0WrMO2gZ0ZNcB5/naZY4JGMHntHAP8hFtRxCiTZj5HmFDUo7sDZOsHX8ML2KqE
/WhqpWMJgD3xm2Ly42AB81L+ekwQG392F7cKo9zYCSr89K98tW38U/uz4ugc0jssJUkmYYmYgD/t
z9ouYaZV5MN8LV0vQYiAz1aVbmy9Pzzv9++u2KQFBraeXrwMaMcFGiZOW3qM0Exa6meIt6s5+jrI
Fgx2cnYzE0ewkla8HbFqXfOs5ZyT+vT1kq6T/3Mq/Wmku1s9Qck5arlRfMHGp3JjADIr5qI4BtCE
ca+GNaNDCXHsknkIuAq0y8RV1SYOgyPR/uDxjDZx0zhZ2aADE/oVEreENV29rnHs1T+Pltla1ubd
sV91TQJ+M9xAzJc9HL47aiYCVcgpIT/I3osDSbHRB8xcVZjbveTSH9vLytQIyvp2d45fKhah4ABJ
GOzsmRpz59lLiHLk1Q7wuoGVnZSjm9nTqbKeiFccTrrAj2Ce0T6AtaQQhTnOZHDi6b2GAv9o7P//
+6C23rtS99VTJCIvzFxyZl9UzTawKzN0ZL3DWr9vQ/NSGrqXtWjSyN5HD0yg1I2z7OQj2iv5O6tG
JDVgaVQGBoMXzHKVsKMv+l2WVKPyELzgD02BTeP7veHoAKxl7yne303B3b+T4dCOY+E7ChUjpI3V
2oy+Ul3TcXbE/QlSFw5rCG9bs7Qr5sTCC5yneE+CyCQENp2Tw07FEh9nDiKfKdWepPi8buLf/CR9
/gLSngTfWoI94ALyzkOfV831P34JnLsb/NcD1bG7TBv+MAjZfpO3pUFJX5SsKHhguXpPJZfXZcdj
c2lD2jkePES7psMKfMVDPxbwoqKpU5Gm97wIY7GP8DVnt9xpPYVmSYPPiFZR2ZOO7ltOviPjDiIe
STf3aYmXaucRLMgkNLxh3QttuFrLdYqhOkZ6Ju3f+CADIrgTaUPEvPIdIXflNHERLTV3Eh3FTkeY
S9RaH0GjXMF6fKuB5/8O/67MHV1IA8GNyE+NjeqmCjqkUeMT2+j/4fWgmiQyECJpCFa4F63ei2rJ
9MdcfSuAuHhnspAOZk9bkVK3VQR3j0M0r/AG2Qy4qR7xsmZusxISKarYZExrF7LnO6TR0tcOMK5K
hMtlhKF6Bw14QrgokkJPUUa7qAxcl5/20Zg9S3gE8irA+YIRJPRA2ihzP4cMRT7EOLoDUKUAwErC
pGGN1KaA1n3wHd27gGx1cci+fi1Ax+hjK4rmWY0AlYqKpRnqaZeiksmrBHECQlqHcPUF+WuiOZSy
UJKi9DYCXFo+FaNkmYQXWoDQnfi54//oFHQ/CmHrkSTjrxg6HE4Ad/9OHCKDzQUGQhiTK6Lmkqg5
ssiLw72EBdNU0o/v+hPhxySWgM8/OTxq8+QM0hnyrRXfzd5BTulP4yjbLeBYyMskFbSTZLVKSxk7
2bN88XEM34chxWPbscs6kmfZcidDo2A3DA4fqh1YaEPjN+3wNTZz3co0HlcTKhtI82tSJRTkhq8f
oZp4HyCSHHLb4LA0zEjoyG2pVcLkiruz0zvwZQWG4HwFIganrTc1P6U7ilB2+nW+UXrQUSHKRPgN
FQMNy7WlkaZX34NX1lD0Dio6feyV9ay65Hbw8hF2/zVXCW4XlLPh9zV3InqzlaHnF/4VTBZbrN/V
F0sD2zsi6uhNDHypJrm+X4sIoYFfMWW8VhIIi1MvwdGxHo34cm+ZblDGE3/j4QKuuDzCl3Q/SvBW
I9MzpSjiVVyaL8uwyiVkQyNN2lgz0zFiCZrDKUUCPwsLudc62yJn5zXXHeIsQYOjQi8GHPYlsyT7
uxet3d/f0e533izq8DBkkM/Cwav0tfiPVbq/cziJ1wES9fnU0t/6O0ujDm6LmfhOKERZaus1k+og
pk3TgDSe2nQpzf4K4YcbJ3xtYMwI0swVoM4Wty7hFJD7yGDXdMflIGBHP3wJ9waHlfcFvUE0txaN
RIqIGZ5S7Vk3tIq3vxdR24xBWO3ixt3RWUM768PfiLtOwkR+his1TxDvTma4zW9OU+RH35PTt4nk
Ghhy4hJh/axJTj3yxi29QL4HbtozjEvlIr+s1lVt+GKwflTzvG0Ku3/LGYuOEqCJmu3++I0z9VCK
4igc20XprTejo/OzX9JP0Nd5uosoVa5tDlL5hcsOOoYaFZBa16aQREq0KSq90BZsJhE1fKD+LLsE
yFuXyeShTLEaA5QjoHcB0GMs/gWE1ufCfmQRA7QrLnmiUQDj+dJbU6gSPe5yrp9nQGrGJ65807SV
7uTCg+QRRnpNtQP/fHE8T8yMyUxUIJx91ZRegxPknMHcKUnyVJfU65EmuLj5e3pW0Lk1WCtg11IH
NskHv+DBKl2p7fRgmnryJVFcLx2a2U56oRg+a6e1N8N3xwYpXC+H6Ycak+5Gfr2+XKdzkC+qAPbv
UYy06uyRE3FgBulm6OXCv6X8Xx0rTiNYsitbgoK9V077nsiCSRD9//Nvy56czTMnxMo/s3+TquRg
HOBUu+pPVSCtv2sWtYfhG+aQ7CPmaw2H6qxDnUUn91f8PJOMkWtWcDmufllQ1E2Rqo1tzY7cjQgn
93wdPTW2FYfN8vGXiuwaX2HJy7P76dWLbSNy5Bs9vo4zOp5FKv3kzdNb8NAA0FNZy5T2zx6LKk8q
SGl3HRbz8LeZ2J7mcTwO5NFiKof/N2iRw27bCQ2cdzeb5/uBpRIFoR+nMXH6+mc+hbK4GTKu6aoa
lE15Kgjl5YAQPcYJfkD1ilOopkLo2qA/J2NWlgTAfFPjo+Oee4bpKPfAwy2R4kcc4svbgnrr4qx+
WTNdhZsa7KJJEObxhZlaC7WyRJHnfGF9hnYWRwEVoZflY4GkqE8xxGAcVdMKbv5iK64BDK2TugIG
PF5zC5dwNe0/5/4M5Lkjf5DV8Mx/hz9pcg82u7AgEuK/2Wc981dM2IhfJvS0cXdO1MA+ImkzAfhF
nSi8Ab4b5Ew+IOu4QOGO/ysnRE7OhpAp3JVkPwUll1v7MHMVt/IjdTQKn49CgIwb8oLWVuMdDJC1
pTSqfvx6C36wupVqrNJMZZGrJldBxtbyjT7h9Zal+HEnSY7d+snEq8RAjCU/mWicAhtTi2cPzoGf
z6fqURF30ul8ukLInzjjckiw07D7J5UG+1VkKFC8NmqOGrZF6HC3fCYIuFSk8PhRreZsPFsHnzS0
mCmmHK51Vrd4nI0NrovBuPd13kglthQ905hwqR3TgY2mslZQDfRODkl6a6IJ2l82IOedhFI7koJ0
pLXThxymV15eIkIOE9E1Ex6iMIxAeY4NH6Go3kJ3VRreDCfgRk3mUBDfdOGExLEFVg4ZCIz+hh+X
OxLBWGMgEv3D4tS+/nXcAgHbXg8WT0Fx2noSJ39ZtQCEVRHN5h/VmIkBtnr/OKc4JblAF1qlgdo/
M1fn2x8x4EpOd0BTbblalpfsaX/ouXt5J94Zz26UZvCO+Mft1YIa/4Ye++6BKwua0VA//qpfE6lt
fnvRYmFBfZQBWTiIMu+cZpQLi/QrfdOXqEZtVe6whVRBb09r3F81sRVu+GwtlILc2C8tkHzOc2mS
hXiHYLGeoMmhBSOyk6L5314IHg/e+Akz3zG0U1+l5Rn2XX32EN46mLTM17J97KmxTD+lJ51SC46B
0vCnvmqjZhII7BTOs6TFl8uZCf6y+bsKfJIdgMxdOrFWOQZxpUdf8tDXsYyRd6u0EQWQ5g2zHasw
kgLM0SM8iUW0WFbulx01mQB+ay3PCfAVZM/JM358GBUknk2K+vTXKxp+9KfwzLMlP7ojoMJMlVyR
ISl8XH4FW2MOMSrB9dP2YD6kRnbLyuPfGEAf2UswRa1Y8v+iKFWuviFROYM6j9MLkL40OkIyvHC/
NwvTHigb/bg5hyzCd1154PRHZBZk2p+6LlszTA5/kY2tO2KQS7NOTEM6pXCixSDFXdw5R/ZVqjcE
6C9DO5yYVMcPPfoK1JBtEF0dBKYVtOdFgWJcUIEah5ilDuyqpEeWKsozCzg3Ybi6RWEQy9hUs+sz
GhFBI/RupzKsMdOAhzx/8ZRtMYKggKjH76pfVQ2noF/tcehH6qdsWL5BN7qukFQrLqB9hznSXxEH
ipPCwV+pJqBCEj36s3BMY+OI5ch+1r3bSmC/hPH67tsd8ZFE88D75GpPTU84YPNa3S7anyGyTHoY
YYV+LdgXyf9ewHMMNK2QR/bbDBmQ0tFxYLpwKQZTRr0DcOUQMadJoxAO94zjV5hTbsN37UHgYC9c
XxEUJHScmqQ/wIDaLsw7Gt9pI72ce49bnqGCanjDv9NjcIBDJIIeDQJ4imops/CZvbX/xZ4Kuubz
F3nhtpO2f2v/YApaKu4Ft9/7m4C6wc8CnZR4IkVbqEsivtFMDE8q/ELlmZG5wtYp/A33QT1Bnx62
ZNTGvFCKmO4u8Ze2jVwt3w8Gr0WLjhJ5F19xKaS2vRpuT1fNNqXtNtQY+ZatR2umQdmitYhoNakc
AVXZ6E7JJL7T3l52larMKaW8dDNjP1AdOhne+0JIkXWQlHrquueGvj6eHlTFpR2dN/eN+150/M52
BsVxM1qTd9Jav8OTpknMMukAhA1gilxQxdeFqexGhC3+dHhFkqvr6byZ0MfTA3eqxzw4+6VPaMEF
8qKlfkxGrdJLxxD8LzPOOcAc66C9Zpn55LpWv+ZcCF2izSxrFTvmmZD77WoerlcbR2cfp+fxGLcM
g+A+QpxxA4ciybp7kd1qhKUyNSCfWI21M7QQD3RFc0KYMijC88LNcskFJmf5PamU5LkTiNSchlp/
XfS+wmPdJYhJQWbilDrBoI9rckwVpQNcOYZ8Pm4PFFKkLAfcRh/uH5U5f4xxllDLdVK2rVbTf5eo
omkmf3SCdbpoeu60D1ZMEBJPOZ8RStr5lENEIDc8iJgBbJUX1U0zpS2uL9dq3sDcfHwdxY+RRlpj
g3K1PAGbuzZtnYtfS839Z5lYbRnrP5gyHZheZDm22vxWq+ZSYXuAKMQVW5AHFxlVKR24JGDUruBg
RvkGKSqzRSrJH7OhJPMZrWezLU+Lu52xygY1M9DwEtP31fEKVmyM0AnKdzk6fRhjDaV4scibjph6
wV5pUjs4JtEpgeiLHdzQypBYT7yDV6uwOwUqtCbu0ZHhFvBtkMGDL8YjYVHzBEl6bJoaMaMtGWfD
+0PrmT6O3zLG4FvtKIH/4getAsKeFk/oG36jxGt1bx2qi5vStqQmMaVPD0g3RJ/zwT0nyNfdrKpQ
h4xhxJpUm9wRxcjDkM9RpIBT4ThBkMKmEVldbSLhnxgVi9EwwwtVrQVojcTqtEh/PfPB8u68T7Df
s8miB/vb6erRomrzmJtW2NqduTgpfnnbm4f0D3gsjkRbkFrILZqZMxqjEkeqqUGLhBEiGsco0tWo
ttrflTPp8q3yBJnoTVFgGdmyYCFFv+W0MsnYx20B5hPH6QTlDhOMN70SVtbWyTIVnQMiCheTJV93
eUw2qqwb7iVM6yNv84fo8vrAgTD8QsoYavepjPbymdJFQoNNcz5lEjsotrWVcRH+pvbH+8JNTZnl
i6Cdvts9p5V967vEPP45DUn2cmGZq2cEcWcjw4CL6Carj+FfDWy9m2ZEeJEDhyIg0yHO1KEAMpp5
Mck2jVMH2nQ0LIEjJp5IVLNuF/VcJ54nevqX+FJcg1KfysK5nGZvfGvrz7K7ycH95LFx+KAUSw/G
lwEcSv4C9OE1InON6xGaQLo82Z8I6tka3dA/rXldj2294VBNfVuLV3NsI9poBT2rEchqeetrs3xK
4ADUGdChyAIHykn150YOWT2lKEhGucjn7zG3pv5X/NJm8DjYi9KmsW3TLEUxLAJKU0H0yiHsRYt9
35vPUcUaNdlom+6P/e/lfXmfULFLwCUmZ60OxDOtysxJGqO7CMGKERL3/hEHdsoFIC2SWiHXnWg7
6WUBHtmLQ73QuE1/e922io3YC/4z7r2S+qTF2fadppTwXSyqQ7A8yvosn9WdFmLtu/Ydw7O9Q99r
rxbk/dmCsWLsfr3mj2bor4bzpvRhM20yNu1V/QA+cEq471RgMCmHzLpa2y7wIlGnNVWjzXm2NjXt
DKPrClRWR7Tr6Ez+1A+jAhHAXhT+HhgUzsZZCjdzJIy+lkg6HFqUqn4+Mjqikkrtp+0Cgsfjn0js
r95Mohz8OsIVjSXzMG+J76p3Pi7G7s9q4QLFvQUur02rNqwiQL3E59Ukmn2SixW5BSA5hy1yVPO2
Bd/QK62RBIuiysMrokXbZJ4ie+Nk4OlGvUsQXmEYBLr8YZsrb4FXCiHJazQwTf8fiG/fTAIEv7Hu
zJb2V/btxZwT1+EGX1fuS2iDk2IviC/8PZYFYQb0uhLX6PzGNji9YN7Ty2Pu1IYPJThBkPn91o8+
GXEeKWQcZ3xwM0ArgVqST5hnMSN/nILx9ejGDvoj/KFDXARyzrWTqdYKQcaIR6deu6TDsZ7e1Z+h
mThRQO3Ewiq1nymzogCt6bbYqD+nmI5+s18YZQkTiPX5a/mj0uSq20qSy6s1m7S6uMfcoZBd4Gid
mLZmhv2Wa1H9ujZ/D/IMo20fl1ebEOGrVN9fHT24W42A/KVN9TSwRZv4ZoyTMRmxs5wyiNrrciDA
qZjEFkaoR2F9jpguaS60CHNXUdYfodDLb0TMuX4yOotJ7/3FlamfqPkSFkAlbXPxfI9pWU4HfDyF
2CHbJFXZhh1gXYrf9+MiCd26P+b5XlZjpxaGQo3NeS+PkjpScIFLTzoRW0llkLiCxJ/sE4ut6yRn
8VemtaHOG3AeHikz0znyI7Mimq5pKjQaziFnY/p8fhx1qujmd/xHLfNlkcsvj1HU/xj1327KyJfo
odv/PBM8TvkNCvx2tkYFxycOEbJGxfxQiVTzPjQ1rh3YdsjVL1SCSAPvY2vbBj48lnLlpABzgKgq
LPQOhQD3CcJo+R5/eSQFnF1ZyvgR8OePfK4cxOK/d3ySo/wJX+JPIunA2H4jwf5tNrLr/CyUjnEL
FlGuRrFzcV98UDo94QV+qg0Jm9cRnqE9f9V8AJNBj0Lrp2TpSIC30upqqrAvA7TA+UJBKOpBjRha
T0oV0g0tF8wHAD0y5GoygLS0WD5wQxdz6dB+g2Xeq13vyqagMk93WUuKCq1b5z6CsrbxXjRZNm1J
Fgu9GZPg5mIfSDCxSNoG8suHJcS4bRdzoyONhK+nOwMJSgZtq/Zni5manDoZ8/xDgD5/MX0jtLHl
LW6eZO9/9uNxlSIQy0pee2qC9ccwQ+MLQgIyhJba1PhUxTztdeYrax+LnKajN1I0ZxfYn1J2KONd
uifx8vPr1IQ76wxlQzr0oqtZ2R2AzhoiQqlthYtLSsmx/JKeLDOQdCLbdxyW8o4rsqS87S/v+6Gv
+qpfQmQATxN9i2sKAV6EvdDpOIr0AbMO2iGXFdIeFoT+WmXIYTgUrZpBB2IDK+5sVccfxuwqtCrg
ipQYIA7O7yM1pGVKvTSODFf8Lxm8Sn6ymkRs0CFaVJ8FslYiiF/lL4ZP9pu69oyGyA/v19XJMiRR
/s/Vf3QLJKi5V5tneCkjja8YuY9v5dqKRlkpKgh6NIy39PZzCj9h9Sxtm4gdEiEr1G2xp1E4L9J5
ZPWl2FUjsHx2WU/8Ud4YYCDetZqMSVMv4nwaSaqY21VnQ6v/3f+GQUOKqqqBnpxFX25xADBVpW3S
BU6B6VMNMV7yNpvwnN5H4GuqW1+tRTEut9efCStETR+vBkaRB2qClaGERBDvQRq3VNSTEQ5XjHzM
Wv/3lFh/pGWr1iI0vqjkfpa62xW35abMyo1ovgtR9Yy7k7DZ9YvHCYWEzqeGwvxVQYm1/Afnhr4k
j2XPzsvvjISq9EP8Qqd1ELSDaBddxCQGGJXln2Fn+qGGY5Ar+WTDBo7o/BRN5wVuNVfm1SqT0YMN
1qTv/JNbtp+qcgMucKqwcYfqvQKIIx395bta8FW5+7rxU3tyv2iN65pD/vCD9fFzh/57gAaLmcZ2
q5GGEZeiPAqvNnTJw2NHFVQCnv/NvTupHvJi1EqE4WrV4ZypZH7GHbq+4BTt/BQMawJxEfsQpseB
z4zFvilgmNJtRIYHFGZ7hTgwETC1874EDytB6F2syN+TivzDVBzlON2OAwwVNOPQOGmc9qSgoEOH
OzhsbKJdIu3Sev4aWGu7WvyDxyc8G5USrFWsKyA89qSptOcFvRciHGYFEmP1BWBOJ7KsJmvxYyry
VC53L57x2jFWXRQV52hGEFOzj6YOBEok5ZcRBJZivYuxaG9kIGBnQ7/0RBJOAsiyuWSi5hNJgaT7
AdpfwgBbf5VsBZ+vjeDBLwuOXHqmJh5DlKz689o0nCzQOOpTSin1y8ZZmuRxA+TEfchnFJWnZlA3
YKAFsKp0LUdDDzuJPkMb/w0RLtXiMWZrqmRB8t6KRl9ATI20cABrkjc+9MIGM7jHa4eLv15RxmPx
NxHQiShe4E9Px5W6kFyef6HSGavqKbtLw+EGWXCdUSL/WB2LwXED9GHVHG+0tkPSNcP62iJKpvSN
EMP2ht/xSHiCSw0SN6E6GLY/iNIvFlLfByFEdJ1vU4bmzrubDtUK+Llh9OQfyq1hr7XFm2xfCtlm
f7a+gwJkftM3Fht5MgmIsVwxRsPiDI18p1I9I3kK0vnzsNN8vnjSQRvoCK7WYOoG+z5w3nzs9xIq
+K9ILfAYGqIukYs1kL9m/xZZ8pQ1Anin120+6bRvgIjDA05vhYnxX7TcBWrPHHnvwLH5rb4Yaptx
VviNJdWEYLXjERd4xxdg97BzuIIgJGw5fyA+Qy/iKhrKZuRgdUsUXXWORgM1Q1aJeHtWF68jrKXe
1eeFZB5qOg1UVqcDfudVyn2u2vmu3Axp9R/JZxKAbGaFcQ8O80qtI3szlXsvZ/s2ziZsWnU6C4ze
YsIFlOHBG26oXG+9OjWGRZ6SfHkcZiTrmSlG1kYDTJAlTgoX1PRA1yjYceeTc1LfCvWRPF0o1aaS
7xBW2O6Gg0kGAKQQWxJmGgcxCGRegOlIJhXCKbVZY/sEtKB0U133rZIBTdqDPfV5JYotll4SjxSM
P772AxZomI/zM806VTBXhlSNzgN/1hAqoYU28mThNPKRG/sdFt9eKFvMjk0TOYC6WjDPTT/tosQw
OdAztIxGWx+NnUHTzSuw5/DPXIh5B1A6BS0yTWFUQ+hDeqJf4B8pJdZRLhfJH3r/9b0pRo2/0Tac
yijNENUQO2UrnT4gqTQLvxeVhwT53LsFDYaDVKDLoMJrvT/OwTs4hwUaALwxC82ecYjiQXZV0iST
K6+rW+phUoezYi+EF5w4iqrc98rc9nIYFyIqoOb8OHm2nPJHlwnMcFYehNKY7usetzuFqsYIdZEY
9alSl4N1e1KKJR7CvTG9pvEZ1j5PT64ynBkqblkqTNMVFBBm7RNJPUstjmmw7nluqSq+WYDKwXyy
0Zv6EQ+MjfNdrOF2QQeE7SwB0GlJE8kmaO+CWILwKW3Rhi3gZ8fAQJ99Pszx0fxFSaeRIDkXq6vr
vxdsluLUS5ss3kPFOHTr4QlY+vfEO/4OFF9x3pf+ihtZBP7AyCC9cA+ZU6TfgvLpM1Uta41X8Mx4
lHQjIchXngNISEmgLCaVQoTorhfsPqiavfUUrXsvE0S2blN8lLLAeczaaJ9IS37QY9coVOw0/Bk/
S1KQN+0H8Y6NhvrZxwZaoGJ5R9vIk1NjLihxAvzlI06ddOf2S6++Z93mBO96Yx+qDRJp0889VgSc
jHM5VH9NFtTm6eF8bOmC9+UvtYFOOIG4jvy2kBOBu7ubdbHMV+gJePN3AxWIlE9GcDIg8P0b5hMl
VE4bWdq8WoxlYVffgp0RuiEhtQDB5ntQPiPWdOKCkpb+eSJ3eDuCiOeUmskGqR61OLdZlAxDCCM8
hxnkL6qFJOqv4cUIpjgmkEf+MhXeOs4haR7ELMsKh+sYRPpRNaWDbZlydEtTG2YakC/bpr+YZ0wj
BYQePyYXaw6Mu+2xmg7T5do5lTqK3PEUWsWat7dwOseXCmvvfZYiZ/uCnoATHrj7wKspFkWonYLg
xi38T6MFyEEuSXA20q6OBO+YXk5/cq5hMudYh9w1GP4edDX7g+wE72EyZtKhxJG/Y/DD6uB3crEa
EiKorpwUwmqnJ1hobVByuJAwrdohUWlC3vGw+5byCJ21tlAeqp6BsJGp4vAnF9S7jDU9XtJtXkRf
YwFNqJWjzmx1M5R4/sCETiK3VMN+UiPTY5xQ2zYiyajzp40opBJQJrqmYuoG6wlk0AmH4PnGX8Bf
49JE/7hnU7r3n0ahjaBYTnQ6T5PdTDDvCmyEKCt0JQO3IrH9ZQN58lD+mtRtEWCAE6iiHE/PA+n6
zTwS005dhr8t21LIGo9YzKy6WpMqVO5uKV93su2kIdUO0Rl9BAnouKUGeZ2scfWGH6W7c4xDcyPK
NEXjAgrRmA51OCH+TYBZ7Ql2i63oGU6EK6uOSSQCj9bQiUdBH9WB/hAev91TfBwnCSCCFAeMjZ+A
EYVrexZgl6J9j9bBEZjhMQMNueeEbUI3LcwL/Q1+NvIdpGYVYYopAywJFrmTN/hsXMGiLfOhpUtC
9OHRFCQx5fgfwk3qax+y97wZ30hzMn6HzjIHTn7rTA2udtGZ7QRJSV27V4k3Wje0THdkBUyNg/yl
t0n4BSnLfFupkC08hAOV0ih7qUFpLX6g86MeOZhxAj65Zi2gNMJti3D5FnB2MKUHairaHoTLYZ4h
9Dyd3b47gsLLJxZHogH7olCiWKJ57QwMNPH2xK2mx6HLkVCBzNWphhB1wsCMLTg4yhlyuPhrhpP9
JCK5iC5LJZ+/YiCdVYd/s9PhkPzqouDJ7Od8A+4PQNaoZoNOasyGrGLZ0HQAGFUoQjAnDR3GB5Wi
jmvblPdSU2c7dTnzaAGZQSdHWSbO7p2HrP2kCfgnimEcxK7KtZim7WTkK3pQIMQZm34Y8JDktqRP
PEicV6CuELYjW1eN3KNkMjAH5Iro/C9MDrN2goU10tG0xMASOHopgJ1r6dbZp6ydbH/GgJ3s9244
8FdUsFmzZa4zkeomuR6lsiXA3TSrUdZq0wiW4ek4ruSCs4tAX4Ihfz7pESh103zANd/jgzl2wkMC
gR+UvRoiaKb6djzB9vWzWr/YmrzOua6RnZs9KmBa5bu02E3VHFnbY9BqjXG2g5XoMWXA68VhywsJ
Z0nXC07nOan0z/SXTBS8VYo3It0qVoEVqvgpkARpLuY5eQM2GMyTujVrdvef1mCuDUoYvCMLCYeQ
l/J1SHjbKLJGTa3wCKJ7VvG34sxcFvbjMUjPneZWWR4s8+qXQ4VKADnpWhWaqtYO41e4C+yT6+Qq
/MgHh86qyToari/KcQD++ZJoTt8w13x2SBP5obezmKy1+pS2ww5jHLQv4AUfCm/0/ZXjrqgjsS1i
1VOtRY4E2NQAf0DVbtqwUvUddjs+DMDNTF2o1PlFWzjYBqf3ZaX3/vPhnQ/JuyyDgecakU9nSWWJ
EZve1LS7sC1XpCtR3glUOBtw/54Mhgu0bOUPQOxLijh7hJTY41XVHA9NevNC1JEoTjpEFqDHTH5N
6molaXPT0uY9pYtMB4nUSy59QOCnpe9OUx0nt1pgRSLq0P1sskr4oos3dofPb9/vxgkRZvXm0AqU
PzhnEH0rXM1w1jx15N8O1TDyPslNKYJ4t4shO5fccHA9JwIcV+b8FF5P/ctQ4oRM69zWv6W7NhAb
1jtuTd8qB4VUtLhzpSJ+8U074r3zVlK1n5tiJMU/sa8fcbjqNqwaMcTjHY32zH1kXwvKhUR/Pz7Y
sobAd16CpgZX+0eXrUTEDW3TtUU96wsAHtM/xViIvmmXnJHBdBoaHS/XNVVDJyh424kdU2x/D1H4
HdWSE//XJco0SbHDkFjMYOuRCVrbvJ44+SFeXTkQ4zJoap/Vz8dUdf9PCI5l2KulsI/oUH6KKrV0
/tdpLmfDbHF+T0g5Amv7pK8wLc8u2QXvV4L1AH3tb4RS2QJOflM8YHw25XBsVsaMIQrjoFX3rjPD
lapQ5aOWcLJ2wrsNpa1RU+GKu+VS5GuFjg8qheiGz1sb4zJahiEgVK/m/DRxS0zm08AnJmN1Hj97
AOS72iqCkBw2Ag5Zze819meGCOlWzpCzHKZvRi/EGAEGkOeWFfkvcXFDTeb261xfsMHGsd3KEtjO
569TWvy0fUzJ5NuGY0adMZE686Ir9+xtd2wEb2gbFwhN5AfJiWFYSS09aJ3g7+TGqWF3EHPLYB5+
H2uTY+kCuofatftDriuNgIJIaIhGB9a5zuqD1gy9eJOmA4/hMAxNSCwugWodjRhFSDUB0IhYemKK
KepNqQLcO7MUoZlKeGROOKijOU7I0uowd5CZ4+MQx0s4rFzMziSc34qwg+D9YF6B9XPIAZcVRqje
FmCJTJLSMLZOnxCo5x1eHuEn+6RN3FQRxqBoUpdE+atsp5ZRv1cyp5kp07kKyR6IHTlKZoxK7d4j
/waZ+ELqIpwnx0oerqSuSvZwpSrqeaDig/DoQbtaMlm+3eX+veZoBIuoJvhlzN+ItengANMv9Ygb
khxoJ3/WSHjw0ayxeeSY2SmyPxKeCCi6bdPCulckla6+u6l/VRCRAQyy7DFXr3Ytc3H+lx6Ae0kD
q/kUTyZ/aXAbsVPbZIfkcVrJJuRnEvmuFlQ1rAPQDogJ3ZM/NRmPdE6mRtOmTj5CqwcTDWY59NYw
Kj2p6UqJMxIUeLIN2X1MqyxlZ96gHtkGk0uJ95dP1PfE7rSmkFV6t5VjccIoK++ZZWJPsDbnqWEN
CjZD2V+cC4Ds1NaGVoTLiy+fe8u4P8kLh6imKZM04aaZMAMk7GNKctP/a0H0BFtLCYiQeWALS0iI
0ncMTKx6bS88v2XrlnI1bx83DRGzo2G/pvL7YWU8MFuJADIKGcq7QjeyRg97GMOXmRUiTW5p6rAm
QExC6KJ56n+zQKpx0zvNZ0Fq7DWc1tr7MnNwZPzUV3uixTuP/3fXBfEVXc9kHt2+6ED7bS8EzSYQ
4PrSkC1BFBWbCFfx+MXEAyCQHK1XJZybjXBnZ4Gv3gs0BUgY7ir3QjLebwNFkcZ1IoUyk0E2tnrZ
LLCpMbdaFdoquELetH60QNAMrfnW+BcoSvO+/Jayc3tb+5rt123KcOASoVCrjwmMraxvjBoQN4NQ
nz7Fk3Hu2d0Cgo1MXFBeJCphHFXCT89hHOnl9OfHPzvDlsvZFUx1ZAg7PqNq3RMib2rtn2mLCNHk
zd/+I2h8cZhmzs621RtXY7xLbh9dUb/qLPwKxacV0O/rDx6F8fakmikFG4L3WSf/gaWfxOvA8X6k
6MSdfYQOvfBs6Q403HFTvGUM60ARJAQGai0A4b7TbvSelG/LvkwCJ9lFQtxcWpzYFqrh0D+DmC8x
7rlfVyyuMtLHJYEwWr+bqZvWzYB0jtH0KE8xs9FKfz9a1ejDmFzPcKrqiknoNCeN/Tntu78o+7Th
4Azu+cSeHae+xiNVxQ/adKeOYHvcS3SkPfgQKDVOcf4nOLuLnwnyWHe0aYBwPDkiWaOiv0b4/8jZ
VmAf2FUmYljGZvMC2s2VYrhOOFA/UBpLLxJ/5HxaQv0pQEpJf6mVFqgea1USG1YMQtlwtQQEQ13t
BoiJNdxJwIIarQX8VEr/Oy7jfv3jJeIjx9MfSDsxB7YcnuXgpuEGi2uwIQgYcZm4+YnhgNAR1DMd
l+AqsbJMIoPrRmJQWT3qGzOvIGfSdU07rDWhqzjLnDTkum4jrWv+/i7fK37MCvUziAaMupjA3h71
J11f4IAqZbe5qAEdWaGQSTjUu5SCloT18+MNrqH9iotXjoY6m5Jgq/++33dt1MuEHH1fYhmAA70X
uJ3TuEHxBTVI4rjatxTdBf5XqVPUNR+m7dGSUDyjGB5qQB9bO+BIcSzMYtWikpNky+LHxQTgPm28
IRjgZR8GKvuHqBeNPXA+ktae1IBpMS1fYXIvewzSjuKJyYHOlASYYzX4oZ+TYpELtlyqLdU0VGyN
iytH20RcP04NGq0Gc18hkmWVcAsVFArjwGAa99iUCAjquDS77r3MxaHVIv0sqqHfSscv8FDZkj45
afjFL7vd798D151GidJmS58qnRV2XAnhr8Hm6yIjqWMBiljeYi+iNUa0mf+qB/TVnyPjjyR5WERI
lesYYtNziK5k5MDQKfddtrF0+pZ77ZrPG8p/K+YElqvo/umsTGVwZ64k2KsTb1bOq5xSS0wQHAon
KbKrDnyxaQTDTDvzp/6n9mAJwhWyx6Aox+UJ8bOOKcPiFm8hY9EViFd3kBqC9Sc/AvSILt5OH4SY
P4/7sr76iKthbyDfjis4eR9oguLWzaI2fuOiViDubz1eaH2xuR/DAQTqqh0CnDWQkl9rZNd55E9/
De0V1x/N3imSS32YJhFLKkN3u/GGof+X1l3H5oyJR/zgGjtD8FBEzRQ3ShRIg+xLPa74iUylHFYU
2qPHg0Uc9c2ApCnqCWopKhyjMQvgJ/3fs5SCMuxO3yN1k5K5vCQ6qvmuE7VLTDg9mXFOLVfDFmk/
nh0tvYVrw8MDULHWDkBA26FkG4jn2+STC2sCxIlJxoeoJSuKg4+qdBhMbxXkdEuqJVXig43LjpYw
sWp1XkgZgBqu+kiBVyV7ZBpewqtRLPD9aj4LpevV/FTAhNBdDxjzSeXSUoV6GBEqgfc3ct8Is2JX
QJoad6NCxjX5b/g6q0WN+ZZiRjdHbiwIaC8GYk/PKnVzMcEFG3+x6ijzEX9PKl9hsX3PObwBynGS
UFWgYgT8u8mezhCUsCP3lq2kGuug79uBuLcTlYfzlaLSZQeAfUGz+61dGCsvpy1CUHV5yHg9+eST
Sv3viXvdT0tV3IM6O5bKGdG2+CdqtcNtaol2eFaOi0OejXXV7EGvUh8UauKk6/vMDpXsd2cBTtrN
ERsG3hcfuWczIT2pUvPUUrx/h+i/lNzmlOZ8D11IvD5kfM20uCVHRb6JTzd00+oarG6qfSZtHafY
8EOZ5u12jt/mRhwaZJ5KzVgBOME8IcZTKiw4ceOsQor9mJBsq4SWduKNFn3fEYHz1ej4jaLL8Ek/
A+fJDOY+WM1SvNlQceiyUdbxtJu0/2c0g+Qkoj+DZTy6+jx8XtGD9gKJr1cRdbPUGmZ3tdV8+3/h
6PjN5W0H9fNc2rWDi3CxKFkGmbLfg4nX4aci+8vI+YntNrVDBMjDROw9ejJSyisc1IEz2r0Ey4/d
SaSmSABnN6GqL4mjORZNwhloojf3/AR1mC9TQuAZUYPplVXcwUhv+M61wfcq539NbtS6XiPCAOdK
zOstt01RRo8ZHu6D/LdfxnmRPHSp15kYvJYSy6DwNBMduWqZaQIl80kQc6n6GK02A21nChbpT97s
SqRdT91+7bPGPWm/xOyBHbGFkRfBD6YFXxsO6pB3wpBoEi8yXkkQdnbxiuDbLOn5gOWV3Yyns8UD
4BqDF5WY3GNn/Yg8Y2JYVhDCv5C11gAwvlAUggvf3aWcB4J8WvK6x7hvQf3z98BdpT0xXhTEGy2q
TnhY73sCnsLLQuCekgCoaBBhFXJIB84BohD5vPszo4ytckx2SWCg1lSo50bw6k+0UFUzTGaWqscy
NOg/PTMrV1ycK299w6i4qdCdbOmWZn1c52JaxFpjVdPE6UfRETqIktE5ekL6153g1S+7/H60Rss7
fuCbOIsmBR2QtGoOBTRPygPQEqB+T325KDE73UnIlvEvCiOqeTezDCVY4vvZM4eNDBbWMQX7AmUg
eByx1mfnf+I2jDrvmrXZeQSM+s9Osv785VXC8XywOgNWk69jRYuNQ84BS/+7dVVLwae4wyN+/bmr
QS139B9iaxvtc/YiVxBB3HhzGgpfuFSPX/XctVDLNqMqCKjZ2hQuADihrdV4lSc8UyDwrduSFr2k
wSP41lh+waTmykcGPBwpa8OhliBxiOHJ0B2IhB5OaWHN1gvW+x2Y2tygDnQHyhBE+UZTbitNlFhQ
JmOwk3NHCvV4x8EK3hZ9RaWGNTlUQVgIuqI8T1ID63YNszpfSYHNIzuSVolYwOxZKj1uAwwMC2f3
wEILAWjYah1p+FPPPwi9Pvbsrrw46d0xFZ+CRFjUq4vebEKxsROmrNOQ0BwAAMwv/cMvovnSSarI
t83ylY0nOpFRjlKLMXgExI4EGVW7DhMWUdXJJvYNIrOH8Csvf2+dzkA/JEPjoE9/j8oxSmKMS+g8
HC4KSW1YkyMakpbST+eRuv2M1vUBtEXfYZC3fE/mYCfU/wopOFRoNnlWHvCZxtMZ045IKLxzMf0s
U7dCU/lylSlI0w7v1TUbN08TkYBlcfRgO3gZey2qSlswC3zOwqOqqS5Y2Op83w0/nvvPxq/iIUoL
8bDjk2ISP3tC0XYFWkTNqN5zMOlJloXdmkPW4NDduFc9MWC5OH6HiZ6ZCA1FpAGfocoutWpDCPPT
OSNZRvgZQIDqyZ/BKuYXGVP/mksaVuGd9RnGEktBvGpzHMaGGSsjkIe5IaGA2w3caRio5e9958v0
de/R4P/BDiSyM3Sf5vjk5agm54X3dZO3MC++gBNt2L6tfMWWhB8oeLzbqdWKPRRN9A0HecotJyYb
xU8gfazLSoYYDCEkWsB+66JzbHXVPZC8yL8l7/JNCJtAfkmYvsU7gqW7I/vKlHSZiqYEpzjTgHHU
VN5h0OGBaoedwArzk2Q7134o+l5ExIP/h07iOvQxCg2yUCE9amqu4kgFX5sR1w1d3WshsTlOY31e
GTv1aPIpgMKykIwy1HBKJNl02aDoSOOutms03ILIFtdVW0YKYVjE1f8zRfENXRIUH7HLqhSXzM3J
d+HW3HHWmxGiFRqHgZHjdnUesTaZZ5ScpzP5USSqDVEkRBrZG0EPp/9N2M9wcRVwhOcwIX902miv
gb3bDs+Ax8nW3S6HtndUYIsPtsCH2q1bLsVhYfNJte6gyCaRx764NshLaHJ44FyPQucIcyDoddU8
Gj5lcNdOP0G1HrQ4yevqOa367zsArX37bWPsDzFzgRHk/BwZtVUXPVqguyPh/6hN8QUoy2mBtDBP
Poa7OWAQUUMXgmMxdjtUKFXr5VxoY2+aMnG2MRbPoQD/mcVF8Wz9RdnTC9nGyz1dWhdK5Yc6BZcR
2o1tFsPlvwM2cob73GcThX46iTs8Yx9+5ZdrkRJGKso87iZVXtSNNDVbhj3UhT30o8oJwq1pjQhI
OKowSPSfiZNy2Mm0EcmiXMPLiVzoE4mKrafkHQ+xxPjDAuFkFOG6khCJo3eDJAjHpBo4GRViKESh
RjD98uvR61Z4yUY39CpuW0ghRbzFCaRBNLz1gVyLnCGse4AH99dBRbfOYy6CDK0bLysBnN2UZCDS
pk/UGlpL7W1P/ECA3+BUHMjLqjXhqTV9ZVbj8RqI+tCbjpW515nnKGZKs+DupDODu14bX/cGKLAf
SG/GCMSlOBpu2308qIa0m2ddTtS8jbc1tPbC8gdcbNGuqXzNsyhwmAZr37DN5g6CxgA/gut3Pyld
Rr6Z5dn6hfAFQmxjH/nbecEfc9j6YpRSFDK3BENJi4Evzw0hBAiXw00WCWm50hOTUrJyAp7V5ReT
xWeYyiHVNhvzKHKJ4t92/L0qCnFhWqJD+KOe27I5tfIN5xsNtFNv+rrLOW8KXPeCZ9HBumNlZh2K
9cWK+cUjv/F2r+J8/6OcL5dabi3fpRRBNiL39Bh/s3erUpzeJut0wPiqpVwvPk4QVnoqcZK/neos
OUwhEzXd2+y0WPYPOziC19cx+jBM+1uyrRb4oqXSzGu9BvxOpHo1BXfvOYSET/DBvc4Z+B3sp707
mN5jrVFqO8QxL5Q8iPTN0oBI/H2ZpdKzUCJTNPyDtP1Bqf8zmZ4FvuoaqnS9dhz4h5X7eFoCUV7d
flYDbZgMhVARB3AxWupdwouPET+nCH9GZMFf0pKegnj4K84QB3NAQI/EJrG50bv0Bvz0C756eHMC
wzi7c0FaPyD1vqgn+kqa0GHa1NkND+AfmJ4Z5ibqF0EtpGn/McEhlRM4LzqYL0+YF/Yei8CxyyH5
1CTzrwybij7vheiD+VMz6twtbkBYle3FvwLhBSKBjMbqWq8OomscuapQWkqoDF1pMfZ1kqHV5v80
yMhwPXu+AhRKI8aInkQ18W2nJh/MveQD2J6ui8HGq/J0ttM/4ovQV7s63Z5jXd5JgekRwcY3uxLu
wMrZPAPkgIVsyNYklgUkG2jjXhJYAqMcSMjgKPT8cR1yszHLx0oT1v5XifBTyCYxwtendQI6yy3b
bpq5vUcBh1krFIVFluFn2dLGZ4djx7v2v2kVHZNVjWx7KWifVV7Taw6tXcxIgcs+1gR6+nG4h1cZ
6pQR+ba2fKsqg3/6PKrMG9p1Y64ZG9mNlCp5OqqyBJR/ZoPG0Tc5Cs5IMxlrFycTLVc7/DUFBDqJ
AwLma7CLBrja8aIQED7pMnKhDEOz7ES1nf+MGJ+mgUrF1kvXKS68fboUB39MBjGm3QcJIe0iOXpo
5OoTSVBbJ9MFSphLcPIszQBeXlLYxiqi7focWtTDOWjBW219ylZ3r78S5n1Uxr1iI3qYTW6CezHT
IA8+rRtZjX1BqpPlN/qo8T8fYrlFwLyLSARGM0rn6sF+wVCTmbGbCW5hwHHkdYcBrvFQNzLPfnIy
riVjKA23hI7Hy8JC1tFzRDdjc/QOlbODkygAyyNdVAAGR4AAxny9YI86/o19Ca9RoXxIVQUnz8Zc
4ugTBPYZgXQDEF6GTVgEMkAMcv1FmZPuK9ozT3QiCpmAMvQ6XP+OZuOiVIgqzduolCMJiZ+WChTH
UPDzn7EVL8192zdbtFkwnPRntpvnKy5lcEEKr3V/JZPjuqpz/lWjn58z3rEFu/SS+dPa2MkPRk9X
4tUUbtIgU3k9emv+J0zoRVsJy0VYBinR9CPfuxI8MwX1G2h2zZ/Da4BYVp24Hj5EcBbZQLZgLZSE
oQ9QCa8D/okIzazGk7jOHOTDHSzj096pwxWY57o9BB8J5u1DhoXAshPJdVJsZmCN7qiI8zdRdqXs
MIYTBd5xuYc3XyF0QRNlua3QlAh+7wJ62bm+4Hd/+4hp9DfKEXx6V58Dyl2NdfuWbhxesmu7a2U9
ZLubTYqURFdVb4a8yQePdL+zGEDZhPkUFLZSH8HUVgBaXUBt9Ldle/oPLJbbgdgQLs7PI8XCKjdX
hrVuvidGkBn/2rUFURdl+KGKI5HKrDLUduCpebCVPlt7XL7hcp07FTdLCLlVKpoGOTltOgE6cFr3
bzJlRDDlDMj2xyRDskSdzDTIFiXnWokXZKKbQqey6TfcD4RotPon9G/CZZwWQsYf2IpsWxZipdzL
hJA7M8J3rE5w+gYJuxt4WGkliqX5cjCT9/NqVFBAvHVW4xEptVBiuNYUYhbck8ZHtA1LvZntAiRq
XKdXuW6esO83OvKioW3MSpIVIuGZ59VQ9K/SF+mVWGVR0ageVVfzcwHEBEjXppPfTO02QQNzY7An
/d2zt662FiskqU+Hem2xzl+YVwg5tOL0RQRAv3Z+dvRxnAKe65lqz1R700pjsqnzmc+5LpVG4lvB
qpEBY8CjV2P+Au5FHiNiP7an4tdLm5FgdRCcEsbP3Ud92UeKLzMeK7NbQhuPYlKoovN1slcCI1Av
BbvZO4Il9wOf/950wbIxfwIzCXmzhqe+fXyXsLnwibBnTAl5uVZYist7V+bwpRs5mOInxTXnt9dr
IYVIRIFemDxvxa/R4C1MDiLOpQWl71oTJqCrckdJOfLAnrjQtsPXKA7fEg5G/mAXqAMVH24qF3wN
WEtfd1ajGkSHZl86ZikTR1ghGbliREeSuNQt/6G+MyLWEcP+AAWbiBqefezTVitF7kB5fy6cjlzF
FDTeKrL1AWxxBylt7a42LT3yZSYPVBtjCa3wwYHCN7Oq1z9Nc6cxlqUUvVnID27+z12G9+5CeUU7
cU+zcCESjg5fbIcXhJaT+sxqlcYNodtlojCZK08S6JPqIJX4lCAkq0TNYXF0Pr9YlagHtJcx795q
KCqMBl4zaTt3Oq2fWqTHbwm4o04qWl9DbtS5q7jKYi6WdwyIzHS3hubk3Tn/Ez1RtdeDHuz+xO0w
7EhKAME8y608ORw5l1iT1wIJXZ0pPydpOHsXLRDXJ1xdDgFQYJBireS3t+oegOS6CKssuWVivUIt
f+Zom+zFl+VvgQ23IDd2PFkv5EK6BnpWv8Vnf45iGmnfSvHNIiKx7ngsRsiMH4TBzx9Ulei6+gnE
tJrnVEyhue4DUU3P5t418KCMAczy2TBmOmat585b3TTorVC8BZemaX723ihPzpIwC4E2TaatCSI3
xCN/2P8xXVQklTKYsnLpW9M9/2CImPTwbQoZtRYRzGL8SPt83x3HvYPOi9QkJ07QkJyKYWiDpfXW
r/9vze1mOdlPfZQFFL2ENPBMNmz/4Z7ojszq3REAWlpXvDksaQ/J4SXR2Ufefu5pfPV6TMqZ1MZX
HmuMJbRQk2tE82uZ0DOAWs5RfG7B9KVyrnmHGk53y9ZFnPZ0rqhjerkhq+AX4cyyeRh+w/00suHI
rllZalJKsIcLDU/gOiQMqAv3dhJPNzYFpOPUoFGhyvDCsP/MGQURyXOn/Tr2hg3RaAZeBvkx3pvi
NuIBmcmfzt9jb4D6h6OaAJ0Ejtea016p9c53cF6e7D7KFh7pfQd5xJX9YVg2K3zkhFXcE6pjlcsK
3pAtgp7CAM3s3P8FcsuRdrrySYtb0cSHTlutuIFgzmOZoCp2wdqmKEAQnm8ohXXtRRHPMUpm2OlV
QHXy6FpHqj3b9Peil9R2DmLKT0EoPs+x54uoj2VBNtmmFSIUVBxHi/Nki1+CPJocxbKdxGnGxbsh
3uHqPgzF6F72At2oNZv10bJh/VULIz8nYGa7+q2Q/6HyC0dTDMCxe+xDfhvk85lGnuazE9GKw/mX
F2+A3vHhCbOEXdDlmqQMdgzQyf4Zs4HrUyVxgm1FFpeTAQn5UtWqPi/BC9No9m11mSI7tYG0+Pmt
GFzbsc3ZOazyiTP1APwBl3yScwHh8s8WgBG0gIAGRsJfSY6Xud1BEgjgvZIaEq7TIvgGzfboWJWf
/Eh/Ln+oa8F+qnKdXTO5dbdJIgRs2B9ZcHIgeLeRX8G6G+6Xd+MBcNmr67jRxhhBnUClgVmHPj3v
UGjeZ60k2VJq6zd5T93Mtz2I04yC1lntzSchWzFFiy8cf6vyVqN6TSsQy/AMeB+z97hDgIHaaZbN
7kxLKeX4No+IKpz2J0kcyHIxc5cPA4C3f5VDXOce1QrexZaQwdQ9DBUF37gExUUgfUJ3BZ+t/nrm
srZ0vimt+lX3rDQvS4dRtiHxbcmbIL2cBBr+lrF0XxL8lpd5/AIiRfExPEQ9LPDJ8M7K2Bd/lfPm
miVeXHKSiJMRPg/BwWPSIi6/tpH9urumlurb+Utf6JWW0iV2XT8k/2r4Ar3+YiFF1bIvk5DHVY3Z
SU/TZ6cHFJSkslVLVmkAw8CepzxIGP5mfkicRHKtD/K9XVrBgHuqBhMLKGdJ/cy7jVF6IzMf2lSr
9O77jyYEK17V+iz5ZoW8wOMuGvLHYvJbwxJ2UcPTUOlZn3oOd8l/RlB3mAat8KZl/8N0HedUW1wa
EwwX4xnrMkZrJ9cehfJNdmYsGXWiYS7Ymteb6czW17yA1K23r3OMc/zu2e4QyTsJBh6FhZLYuco6
LoC0ibQSzVChGBm955hBtwtk81E4gYV1egKmeWMr/eY1/QE5HQv2jsAl0957VVnk2ne2qVOYBWcl
QeVIfBqRo0ikfOUS3ZHfj0ewSPNVq4L/zEglPHf64ekcxoDfDakBDeqAYHUpvlEb2efa+aDaGagn
ihsWvq2hgObD4bjyCYR2Sj3PYyOSjCLzKVN+70RpfX1EYuUixne4VT3xzNDBLBNVS2QPw8oKii14
MnmHNAJ74CadLRXfjJN/B8ODWmiL4+2daARoN+VMbws/rDwwKT5hRxChXfyW/nS58oOYpe11Fhs8
gTUY+OzaNVmMQkB8nQvOdRtalAinNejyzKn57aUSewW245yAAbd7mGz++SY/QaKW5HMGPQe33exV
o8NZ/7/j89RG6vAGHNDYEH/DX90JtyrNh9iTKOxdWJHuPQcmd4/QLMI3k5NL7w7wL6LCaI6/Ld5x
sQi8nNOmTVPvaRIbHwY7fKsKSnU2m2Iey/BEkbTu0N9y2rTUL71D+IhPD8cUSftq2gOIn5Sl5veq
IKDYZMt1qTpyn55dPbXtUg6XCYd/uGeLk8LJf6NeKKIQYLZyadPWRLepGBsQ4Nddezw/E6Tf3vyh
zly9PusAE70ECyEs9VKPIit/s0WDHHWuB1ifKbgPEmqqwl7xZ42dfUraeu1dxq6p0i06G1gJU8qA
r95V6HjNnuXy04KLnzCsrCkrxZ/M2jaZ5dAzT7OLNAa1xEibOiYDGrI+fxLlzjAWAKv9TAFahRa2
OE7yP/dY9Qbv9e02paS7CA6OpCsoeFNqDtNekRwY9iXBLlTRUqiIFdUrgJASt/7add52q49aTSBQ
5iEEvL5FBx42dV2BJe0ylb2EG8L4QAXsQjB1u8kqPApP6yyXVpaMIjZusSjZsZ0UzDj53hnmK0py
Ol21ve0j6tzJnqwnfcSfSAbMPyK6AZdZnuYpslDM4Vx2oYYlgr+IGqt4/1oNhRXEExaQEGV+DAe7
ExJ75ftR+aRMmZsUVuOmWhJFQGTQ477eNrVrptqsu3nUAhiH4ELgzlDkuNp92Ohky38UEIhyY8Ls
SY4gUllehdSMhsgo5IoCa7U2ZLjSBo5DhLmmDfPCCfUidM7KLym01+JJ+0gE4+9zfGYr2qNlkkuB
wDa0ZcRUxu8ojqt3OiLbh/uMfGyOtsPRVbRJOHFa0ufNfgSHyOrNHijRvOaR1bP9IJXsd4fHs48I
DJt8IHuxPlVpRbKOacpl0yESN1EpSlrGU5gVTkqwj9lNLciE6VEJv2jVgLi7zz5plID1AQvj3vpP
/V0yhscnf26SLUR0LB+ubdJ5gretgJuIHYwZP2V5h/Vh3iMx4iZNTaasrxtl4xJ8yNiC4aWSv1oR
9kuDsR5ODasi35MkrrOVadmC6hanZbrIljkV2YVa7Q6oQqFRam9B4/3Y7Gchg4pcMXH8VGYGDC55
KdrQ/f3x3TJS9rqV4eHbfzsskUwpJU1Dao/3nxbEvq1/Ytto06O2kxk7+BeCbZd43K0ozE4S9aWd
bqcLggZkJAA++rLEJwPf2R4DI5/gUOpnSElGnOP/Toz62s9fuQz1u8j3PTex5Z42rPpaYniFz47O
qj3/iDkRC6P7gzJdQtbtAgJ6UyBxkGYA+LOdOIGP+Pa3wgkfmBXtA9os7vJrO5T1kPvxXWQgLUM0
hWKGiRSt4oUg4iwgXrjmgd0Lc9f46ic52v5iW1Wy12PEzYRwLh5a3r2cJKDaRwpci5H+fsUFBcJe
CKO254c8I2ztGbXkaiyLu+AmYMjWDpT2nCz6V606WkSGmNzzkBAp16Men1GeQqCo7Mfq+ztrlbPx
TMUBIbBhWI+HBrT5WYp9FH/7+z2VDo/ffHMyWG+o6hQpD8jIoQhPoG+GIN7y8Wz4x7fzilpHVZ6/
wELPVaYneVoa+auJyTGsAGWV5F9+LPGnAqgiprSOuYZNw4x+e38NpLy1n7IrzfZi73AzrQYGvrjz
PyxSogHETqRdyz3GdW7BqbD2gqwhc7AeyNf7QZ+pdDzmGHvyY5cqXBmBzsEhFLWrKOudHxNk19Ox
+4HcMBxKfXmT3maDfX9dzAxg1680xKqv/u3XSiibqI11z4D3AuxNqi3VJEN2fP/LuoAdS36xTiyQ
dn2zgdWyQSEwiwSURMbd/xSIgxUtqrKtzmFcwJRvkbFuAiJMo7oxJhEexjMSqdMR+6cxwpjKiGVM
sh+rHFfBBDeAGVPyi9OSIkUOsm+3MPYwNywntyNUU4GZEerqHG+U+UVV1gbKJf18J3QLVYLoTyBU
wRVdGutlNxwkDgaamTPnCPOmnObyWbbS7NY8POVyfurjRsFx6HomPCjt6leevlBhMmeh5k6wxgzS
izxZSdXTyTsePpk1rpgjbtKSWD9lzTWISTIAEws8PDgnfFIuFGVNS57FUVpO17Mb7W7Nkv7o82M0
BtSfUaO2OK+jHON/nRvDt6clYwHuK3x4scox9ziDHDsVusBZNqlwXUb8b/5zJYHUmyj68vehL6Iz
kIee5ryLUF1e0ZgbXzkDwbM/tEtQHAWkIoqAsBnkTecMzXkNsm6btzvSov7NFRyF4dI+MwGzFELR
00lJpkbfT8VFG2w40HOAaCgG+Qs2eq/jHpU3+UAtFf2Dcz69SrFi5+jZjKfH66thzBH+95dIxJMK
pfffW0GFBk1HbEJXYA8c7VoO3yn0Heptli6aIswvWSuaJn94YcOFErjYlaJRIgTo6wZFsKK8gZt5
0tRaKYVjAxNdHi+U0kvxS2/8GMypS/V6Wcam8Wvn//bN0M+pp+VKuE0pWZPyLPLxBSnLZKwuW3ke
JJC7yNG0Ct/OCaCj91AiUOU5Vxk47eqX90FmKNs/ex6B8ksQS7tYF9pi/FxwIT8KEUAFpVmrJnUD
Cne/pQY+GyaxTPwEdhzjDeUWBj06lz2qezYZRJVVhHU8NJHinnQGBgCMZkNl6wRFgf9Sb4Vpjahp
59jHZnsrTPKxnZjO5oSlsWly6TPYPr8gRuWrZ2pDWqG8av5XoTrJvrYOYX0FNmnJdwlPd7DQtc1P
VfXA7ftwVhMqJjKZ0REguzP3INLDWLtgtDa/E01ZQzysyk0fS040Wa+rZWmn+V2RiQ+bAVBPDnbz
0xxt2Xrt86RXV/QjHdfAYnEZMfqYJLU+7LcV6n6cCkDauBj5x2JIrPCcZiYNqM6JFFbJ7JyupQXn
LEqwZoFibuWFIENK3H6fQj1UAsuKFRyM3v8OMojLXAR1u2R3dMbdDd2cOce4hgCi2eRhz9crNwz9
ZvUuEoDuIo3nJkpYCwQRsaLx/QhAHNsyMIZNdCJ+j9LKkoDJ9zPSkmhU+u1swl8YLEmzuhmEj3pH
5Vhq8hcpbgf6d05MYI2WkpLaO+zulxLbaCkzBwir+KCaDv19wI3rE540CaLrT1wXK+JfJabmvu0+
ruOp8xUJFVZHuSJkpGCVMiQfRTIK01IqKKFBs1479Wc5NWIpBhNPFDwBt+ahTAMF9LJsLrMIqG1r
FpRv35J75R9xuj4ogUI+XGHS8erx2cTWu0OuDFnKEH2Dk0OE0ZodGE3NOdC3M1IWLw4MShbWKDu0
sZcx8/fUlvph3KzWTscwKiSt1ykLbq3h6Dr5atcaUOU6Qj/3Mfq+Z+zThNqhfRl8d3tPjY3uLt/W
jxC+W4NZDR+W0yoS6dXwhz/pzpUXp1vCoCg8MrhtCcnP0cC4KkEMdNuVxaiWT5htZxZpPuLtZPro
uU3WMqXnC5/PE4BuvLSnDKJOmasbymM3+HuaenhiK9e8ic6dgwoPN6oTQODZU1Ofr+yUtB0hsKUs
3o+MnxfELT2BVsVACb+jIe4lZZzeZr6iig5j3Q7iXGngzz6bQESgnQGBZ0ZSXJoZPm4aqJK2jVHC
+uDBGadbmkKt+i5vNqy0jKOrXDtesvtTe1J1f3wI47y6X6HllP+4Qt1ScDi8g3ptOCWXIDhZnJFg
m746TrSXzkzvE+rI3TJ7NuibuaeXFJevzlv7iy3o4sVbPIubbASL4uW8LglbY0K9tBkIKvrzGiqW
xqTLn+wt692PfEarogP8YuVyxeuXT2IqPBmCP424ZnNmLLqtWuSiN8wAww8eDXLTViZJynVawVsR
RzlIuTd83r0CQ3ohpVBtVqG5ROY3TPx4kPOOiACD+bVQ2TSiN3jHFuYjvftefXIsv1zehnanh9Qb
6NtZB6bMQDsQuCirCAjIIE/pty7/mDmy0+azHzCN+DYYDelTaxP9cG3SpOznUBq8LT8z4NnTlGc+
7ZdAJ33eW/Fn4utIOFUmYXDTnn9V9LejOsELkLWMT8yanEmsHqm21DNcGGveqiP0kK0Bjcn5Z7cH
N/6cmp2xVl2a8uGuzunerEBTyjgM8i8fWucsQFOTD8r1D9NtlEwq3LzVPckXEiY9RHJKbmARPAAE
5f/RHDL68Vzgb8Pj73m1rmnD0Hul/g7EMiNJpnqFBLxQlLti358YiyoHbzpKXzWi+dBm8m0Pyaik
WuscSW0SwYuKmOIbGEPFQ55yK0ZRprQCMnFu61kuBhA+iBBURyf/3YKlvstWzrWltmF2qBAY+kIz
nBEmzrYrRs+E9t99LWzfzOZXSHf0QMKJGMVJoRENzwemK0EmHJ46ElNJwzDga9PMzaWM+vB5671F
XCkNmSPyYYkNSoz0gTXvBlSaf/tcUwNO1DV8tgxjV7MqGruAAEUUQK7Rj4CUrCv8/LhKuHtE/PJx
1OarUI3zVn5RCmOiL2+JO4OkivwVOXnEiXcvrIwoOiKyo07rYKtRB0QeLjN1q+zYVjlX9w3z5/iw
MDFy3sTKVOD2qXuofhLExs01GPgomTN2qjyOuU0jF4NugJqvilLOR8e5OPs/q2kEatseUbCYOcL2
qZn9XCBX4bJ0iXqqx7/F0ytflU11g8H8VIWLrDgLpgrXHAC9WFA1Wqio2otAIioh1DtaBp+EXzS+
NUDBXVBPoZEYEmoqd+VZxsbHgRiYHPeyMvwaRqEaSXLgr4bXaW/LA9JTX39qyAIs1LoB6Cc9bMLN
Z6/vJjvrfIytRPnejzhN31R8Peti0UsRMrqXHv9dG46LgyCEVHUrVBxTsS1pSTBxpKlUvGIV6t0p
0cFlGJ3vZzyGlOGqxz14ACjGlzX3+UzYS49O+zmabPcLd3gPF+294hMdEwZpK0pairfFNR6z8K7K
ixd8Z7gMXLWx3glJqh4YdkHrBBu7h7gTwiiuINWMbh3rJQgofRyWgJiAm/T5AU/YLukgC/PHXO99
zSiCCnJVrM4BvOBGADabF1EdWssS20pn4doDBZjZMftxWi6YpNA/sqKxIMTHujDNgDmQu6r9ONPR
dXtT0fAlYSCiqy+jF/V582JjIW+Pq+XmC/gpBWh2ofhnlXfkgCdAq9HlXc5ieLaToP1/50E0ryyf
aGNf4AsnlGVpJEzxfvXOYnA2DbUOS6wzrEgY9kXFgCQNwxjbmBPznZhb3tJALGrIamZWWHKoxcYS
zL5kkqNo/hLSXLvToE2TUWNZKLg8yAC7yrRUEsXsVv/Hv6sfeSzHZFoqU1/bt85gUCQ67S2QnaAQ
Yla+S1IjREhMUyT/HjF0Jy399JB5m1oQ1UpxB/wWRnabVIimH9G+3Y1BezqBPQ9jkUiHez2ikAMU
C3jLSRbFhhS+01KJnyfaIsYRG4d03WrWs5w/jUB3hGdqRFMW1akJInlyyCub40o3noXNYOFxSWS0
YTEXuWZSkUl7udoS+jdgiDG0aUOWTzaFPOv48PTy+bja6nWrb+g+9QRHGr3rRSSJPSR3z6pwrZys
uby4ZxHD+KELmtfH9H2V//Tf0HD5rj5lIH6/i4zRvlXdJ+d0+3y6uSp4eJVTclVyCG2kuq2x7mc5
TrUA+s1/Q+lf5r2jqcoD8O8yQ7LO3DYZdub1K2GnZJn3HPAilN/UGaxetqZGEd6iuvemFS60a7dt
Nu202asAG7DG1K6xTx5wtPyzpoLExZEth431bZ5EMidi5Ltxam5K3iqN/m05UOiaKrLUbSuN9dbE
Fp9PkOOWxGgVVzCJHYoXHgTHh+82AgK+NM06FX6T3Ah9ANEYe1004toHjuFhLBrXWQS6CP7aT1tg
VdKzWM8HJQqZvKJvYdP6ek/xXy1t89irqxkScdwSwQQLVNTxCGinN9A773zLX1JtsUmfXo4bVfUJ
fyGA1xPWePRP+GafCgrVfBbqjFj/dYDhImGA5qfAdfaLo7J0j58pTR2e6m0lUiF50gXf4ggzAHZS
Qhq/JTRAGww9j+53G1GUgpjbOimL6H1MY6lB0zTFsWzwPIyx2dQFjAwexGdB4y1MP2TC5cePMDPh
XOXuyBZjuNeLnTF8RqpN9iVxHaIrCT4uqCeupldQrPY8T3a5wKycqLDNk6FoYDTJ3u6PSeUnajRh
nSBxWTY9VXj34seNECIfKzOhgvdKdqPT3CRb0jFl9Y3iP/bTwwXaisQI4gvC275/cHMpxY2aEop6
7OmlG4Mo531XPA8Idw/P0uqRpJFtgVzjZPCIwhYBBmf8sfTokNR0z6216ZUYEWcXn1KyMvmLMEtP
d6vQ+f01UV5gMeWATpLBVqVXov/+B/K6IyAutbU6/Q+lg855W6NVIrlnIP/eGSLgtOQL97F4I17f
4fNI2e+0a3qjUMt1Y9lDnRouX74P1msl53LIIAxDJ4C63iBsmwxYRe1WNykBnwVJTTRr/xoku4VU
x5piBDzpCqg2WGgQErpLZinrJ6FMQBS3T3ssb6yrmsHjar8CtuJJjr6n1QYx07vXRbB7fTcc1jC/
MHfD8LP14Za+NFAlOGHu/oEeGHq3VmF9gF+9UMglJx7Cqpt3zVx83UdhqqyiL3tCk5x9P4/2jsug
lnn/zuLtAQ/Qb/w73OWZ442XHWaAAUdexPis2fx8RDyzG+74sX7ieuAvRlvcXtWSztuo+8kJRhto
nGvI42f33u0+iFX+SK/DZxfJmAnQwWxlj1g2plrYxc9zfBXUgmgArwMUwiEn19GBID9Rk4Ob8d1r
BWA4AgoOEt1Bb3mOGMVvrNDdRU36pwKFxOsuGFKUYB2dha4XveIHYk8uFWobQaFCdHzUG7dMQk75
EDpyhMQb25AjG8O+LAliUL7toBgitIdtv3TpPfrVmzEmCsz/vbJjLJD2gQGg0okhTh3wUgBHOzqv
kld9UmFknhBsmagIfZnOYnOIZRAiuteKzmYXzVB9AZ0qKFeYP2TxULL8UgABq/4Q+VUY10XKXOii
pU0exSlp1bK6SchDIno7/IoNYwb9Co+Gb3NoQV0RQWq170a8haLGGVNKDekj6Ndpn8N3ZvIG5N5l
pvd4EWK0y8kAPeqij06AJEJr+rHefAnaJTKs129Sh2seg/HZ5hEAdDdXwLmAvD9kjYlHm/TK0wm5
SwaY8Kns//Ww9dk8GZ/ZpjnRdY4MXTDVVmP97hi04AzpzZ0yGWkoCDgikCUtzbW7J1oUZwMMkAkx
+DcT52b5ru3u0FQtwpoXoDhcVJLUbIVG55iwbq7rLUB+JbiT4CvAIFnIoxQD/VWPapqav99z8tTD
T1XBg9V4FgMhGaOYDVCxy7Ld/uj82HP+FilQeJaKJhYrbDJTAjE0VUMhsE8KupmqRiWBt8h9Ir7b
ctGzmC/M5zYpgiHgpXexIIzgs/B11Zb1jPZJNks5MzWJ88nzzu4k+ua1IEMSF5wtcwtNDyu0Ao3y
KDRMqpzE8YmCD1/5b0oD7zKJcX2y/Hfbf/XhiPyxASNx5iSXkYP8egU1COPVff+7ssHXiq/ftGfz
HO6OHOaLuySL49pD/U7putgmPWwHKIlkyaitV7O3tIj1sf50KgCX6Z7rLcVv1/tH7nepLhHV5MX1
RWOHIy4E/qCvtpHysdqbdWYZv5SdAJNAP+VXugshajVHokLCyQq7BX/Ta19AGDh6xCgwgEwnrICT
+AMSjcD7YyqyaeVY8fwQHl/mi+vJT5fyqxUhSdXN9LheWZ53h4EwzuayafJeoMQbYmdsExazqnUl
vGPtRgZMWE65xW+ATiYiaw3Ionfll5Xb+AB41chfftNA5rAKL2mTtxmGiavAO+irFc6nn2YSNifx
7MmHh+m0kJniWYg0qshZiOYB75Y7iBc+u5nDW5mm3zDy/XSgIYPI0rCTnSwvQW0LS6t/8BR7L6oL
80Oyf3U8XmGRn9rt1Kqb0o46BrYWb5vpXVNYiRRHrL0UuEE7oqkqrbW4WNdM1cn2hH66WmW4tVYo
Zueao83O6IbK59icZQ9nTJf00sYcOMjCgwH1II8Jdu3p0L4ccSPLG5fZkyqngv7h/Csx76zkSlTk
GtP+MqNjX2Kd13gTrqGktxQ0gg1/X+sIqjQFvVT9Fnd3ZzYSXo8EFuTGeEIBLGmc+YxU/Z+Y9AcT
/PPQ2bHYYzCLS1UpiVwVa/04BpzxJODMNZC7Qs4cimL3duZAJggCr5lFlBx+zQLe9Y0RnUzJe8xp
LlayUQ0bqWakgTui+1T6CIcH7Weasod8YmmT8ChrxLMv5EC7SoOB0EeYs4hk2PAWkfwqL0D12uJ5
rVGE78lm3uDgzG3i4asEtggynVlpSglQ4coYgeJw5f6W0yWqp71CgRVHCoRmQ3N3hlULQgiHH6rl
fnWtvNBkWTr4vK75jT3ARHwvpCCrOwcQHnB01QIHkXxQgthUebDmr3uZtBPuOMBbjNL0fgku3dIp
rinCTD3WwR6B7MK5Bal1s7Yyx7rIgqFunImOZbtD3tckCM5AFqHTRqzuBCbWaoNOmjuO4pjU86ow
y7osT2NoHD1/iCIcLXsR7kXtL4+GuH/xMZZnkkm0bK31l4S/sjoZAQppi+XSXCePxU+hEzKWr9Hx
ygfns8YF/lM2G7R3bxJduxfWf/SYBh2hyRCnmJ/Ka1yRANehzdz0cgoup26W02LT7/SdIxb0eVlc
f6THf9n+tuO+fFfqcu1UeAfaYQ4If0lXWgTUuQHwggpyFLbVwSm69WklTccRrUHRLn00biUIu56w
py7Oaa+haJf7pR8fI4EZsUsFuOsyfaDAFG2EWchYITDDByvyGPmz4roQGAR2cYHdr726rggmcViw
PxW3ZFbHL+cKbkscO6xTRcQ+JWJ5Z0TQc22EmGrEJ3BHPv599r2u9A3iGwBNCxsZ2HK389XKCO4p
63nyKxX9eabcDREZyj5lkjYrTiYJnH0Y4ch6z6fTVDftMMBoUOgldeIlBx0spZC17lOrVPGOpzl2
EEf7nL0e8d1iy/0y2a5Wx8xYVDHyUvc+qIav3M8ijokePHKG3AelDfu2msRTwQw70IIbqpJwoPfx
kRA7eTU82AoY0/Of1w3eWhMpiCKuW6wYPtd4ArEevr6KE58Ti0dJmrWh1WYGJ0H4TngatE1OLCsO
tkEHHn7TrXPHdIjeGcwDjO/rjvcuLa61eHOWn5lC2esG6N8SInQIalcbQM2mfioWth/3vWNf48Cp
ZXMVJhe03gep2VWPDt2r/ccNBRqzFRU7pKvScMVIa/ic3nF0+36RvL+2exu5hueQcBllvGWZJz8c
hUT7b76XT+nu8IVJ2NvJZoDmFyPCZQirSPYFuavnb5TRoHTOz8WVIrBFCFWSEg9UZTXKv1rwCqFX
U0beRWj+hvneC5AbHoCZ31uByXxkehMBsZ4PRxsYsbPkrDO6wDyWDXuOaTsesNL41wNHFwR/kMiV
eGSExtlboTDmjolnKERya3cUBjKvWYVtGSQ3blMhNc1o00xL2rgvXejiwtnE5jiAff//EmqOe8in
JUYtBU7WfmJAXl5euKYh7ZXDpFlbbjc/6QrOD1GbCKsdX1sZF+LHopHdE/54LM8SCJN/p6ZIvBAi
s4OIjhZ8NMwzB4a3dVPmzCbMEhvCMIjqcWFQgL2mSOuOhr0UfQDJYO72gRltzLFTkfr3jLmJxBay
Rvj4IrvPpnVpbsC0MSdWmQdpBMXu3wuW6Us0/svkxsQ1luGLF6EDTsfeA8yztYxyDLjL425BrSNQ
wHXwOjsgJeKnV0KH11OmLVSMtJ3hgMZMo5nrwRhZ2u9NQhPnIE9VbXMh9+Ptzutb6WJPWx9devph
x7Z+ldhBk+VobpKrtJQcowxump1x7tYLqwKayMuRqIzV9APmtpOOSqHDEzJnL3c6cSAThnIR0D6L
w+viAra/+fFGMOGe4UI0ZGsiUh69Gj565vdgOYER1yETY+dJdt+y63SKGE0r2IwuKPcsxEBBGXPl
MdNXJXf4f8i6unZaJSz+ZtbpmeouS1N0DgJcPerdTEExRgO3raWt+RqiWgaalotGCkNF88bXzFRo
3xKLr2YULinxrw+D5rl+gZi85TFx4aEkm/IhOag65mZyHNwXorLEBNBLn//qMLHiLTNnd0Ob5gP6
jQsVvu8GM/4Ue3ZwQcHq7SUZmwEeV/yA/ecf3qgGY1r/7qKr2YAqCnZiweIJX4vbzGn/4gHaFR9R
gvYlpOu7l1PvluSKAal4I8t6O8CY+9QNEU94WuMDKx2woOTKpZF65c1ZXcPW1Yyf/vgw665Unlol
xThKdL/h7rfH4Ciec2eX3oLr8u/fXNL09hIjsh/r9GsHCXiBpjJisAn94897WNBH8cFrwgP1r9LL
2XRZtAojX+IjsgQkjFQBD8bAywN+RgvPTpa0phSlkFgyE5XqCfLgkOsFohh3Ylg7NJ2cox8+7jsr
ReNsZRxcNeUiXXFlEHOBjxSica2FCQiFP/5v+Xp+blK3541fCQMNK/SPch1smmRv7gavOQ3mIjDN
qfBiy9CMr0rPOMTVZaP/YGDA//pmJl8m8HX0tkT+KwfjIOKoPpfknjA6DJfLeLt9giJU9Df1zApQ
uX4DbB+q/qCg8JC/2+gR8jl9uA8pjC4f7okN34tlr1p83ey3Lv1cLIPur25QjxGdkcOL5CfIQlc1
CexECKTHP3wkq4h1CPGy2tNyTS3OX7K1SKCo8A+Fk1x7xhyxnGz9IvY02WdAkyfwZUBNeDfJax8i
DqNDjoH9KbReFFg5u5DDZMMpIbZOru6XCEtQhLtLnP+PRhSYvatCSVLegUDIQpnVEnB/IHsSy4nO
jI6MI75OUpG+6JERmplxHnI4411KOxV1V1hbg9CPAPWLR3W2aFDt8+h35LApn1ko0gp9cehSEQBV
0vysqKOAGt5MsPa9wQEtqR2J+hkztN88lnreRUvsYa8F80PrLxIIfnMji8DJKeVrxJZcxNWyIWS1
AwdS7EEVnGNWn/VIZpngRjc12z5CCqp4FPsPdPEz13DVQOYZnKbDimzAV7D0oTNfZMfmPRNz+Aip
FbYDxKjx6xn17D+U6r4Emxa/zPEAnUcaUyBG0CRRnvNPHDYIGkiHpiaZ/9rK8wDa/UiTVwqdqBOV
3VyW9Lu7KcDRsCHdj7gcIhG/wTKDl4qkgBPGNv7n5Kd0WSWyYaOFn8klh1GB4WSVvVXiN1CasDDa
n2tZLFaRGL2UWdNYqlyqegFkuW9fFWNfUDOgm6T1RUna7+sN2Z0YdYz7E4zFlQ1j6mO2xaVe/Dfx
882ExKWxHvRPYtzLTatr8gMIm/WGCUk9Yg8D7YzasF6x09qFMbLGtzBOzDaiL3oJZJTtn4KzvRs1
ZsOG32o+791YYnKkUp+q36ljG4Y6HAPb5ueBdqEv3HgEoHD/Q0heKdTe+WpLcb+cd4fa/IFYvUjf
22Bz46d7NMR5LCEWhVvJRK9488guAblxcq8V57k6ueAjsmUTiXzKZWEzZXhOV5mBs4FmBqtm7wsM
YY6Hzu9ck2A5ymNaVGPB40yI6gU7QuMza0dOgazEMPxd/d7sVuJ9oeTpezYSd7WhpewKZ5BwLdi+
IN0LeLwiSY9zed+O8Yb5+ZlqdQu8zgpMN1Ce4JIZPlF0ZhmKOzuPv/djWnMgui90o6j45NH0yP8P
jlDMDpNrxhDCJbRkYzsKEa0gRPE0aWlOhF7gSXIlbbGowCtMut8oZsdH7PK476tyGD5GHAngKGN3
IJpRyZ/JXy2j2mLwJIz1MDdS2cMbGCkDJ79krBALYgECMvn//dzxad64HgTP+cV1eEg1U4A9QUKp
Qxe+/Gm/JQi9qqkKjjp6ela1xf5/FisObvujAgvpgOsmSczgKDHaEgt726UNTzmGYAJKtUKnL/Ea
4TJXU7iQedY77qQZ35T6hDFrDMw38hUvTF7wUO5mNISbA1+5OM87VtEGD+nnc9dzxJ69a/QkQ+X0
d5herOOtiOeUAsLp9BzruJVgVWaLx3Z+pP1XIh6jp3cJGxdqSM13ezdggsteiC/0wNLFowP2A705
3/1TJnsK5V9Dc05+LVbbldo+nzSZdHS2l1j9NkT4AYLUDpx/JRy5agmhgX9WLFvsohEzHfvX738O
HrIq2ybRpzzHG8AYu/gv2orZaeTrALaGEnbddOPGFkyT7MTkB5RwXX62wum5MwRENLqgcL7lGSmg
2XyYFWyk9tg+Gg16wWF7huCvarbqtCzlNoPJDjXTaLeuEgDx1jot+641Vm3VYfXoh0gKJIots+Eg
MowCdepSuv23MtTnVo+YfpCFGW/WKnElQOfVEHA8HdgLHiiiQ+AJM5sigFqzUBljzH6gcYf3QD3J
Z3BUP+ZOOQV6T77vBU1+g7Vj+qLZQEo9KEG5OfRSs2t2Vt5BhmGT2VHfU5UgilFpKoeKB6hXsZ5M
Itvj9m21HregIfsAMILF3o+RrU4BN7m0FORRQXSMvp83lHIWx6so+S3iH87ezrw9l0brMTnP0o43
9/azEes98Hm7dcjyWfWHmutNJj/gIAv5cViNfR0+yOhqdM/TxMTeYTpNjidPIYbU9iPHnfrhH0kt
xG0CF7/5wbU3wtyia0TWpOFqazpuE7qo7joM4RJypBBMfepLd/jXyQnRfT5fWdD+Nt2dz9A8jpmi
YEFpavHdgEpgbDQTUEIAdGKjHV2exieQQa0HP8ITtjPs//4unxf7rz5ax7l2MU6dX2pg98LXYQ7M
DinDKpYZb/U8jdWolsGSaqkNdKkefGz7uKG/RlCiaYubbVbiCRU0WUglL7eBbubZyfNG6R+P/2bA
KeuHwXbnvsbRDJ3uBECK+8+81+N2+hazeEU2831rPVjManRL0wQQ87E20/O2FUCgH97Wy+zm3vrM
pyRKNNV4mbDc3Qs1gViLh9c0IUI2Rs+WLdIekFRGpMA+/BeBq6JIS63G4ZnLYhwfROwZ8lfZ+uA9
DrWgqYWQamY+xlEHvEHhs6vIs1CxiubJe2uDQDlcxe2ef+CssYhqpMkjlwfE9w8NHpbfKidYq9vw
u7EPdOi1iy3Oz99f50aXqAwmHF4EoD3k4YFjQ1LuexQSncqnjf9NJPqXXCcD6DQPdMuwSbCwLQiq
+wW+OgwtzzhM0HKWdX6W4vGl/cDPE5Y6OxhUL2tmHOd0ybAxPalGS8IbLxc51AgwehF2hPCYuYii
UxKPPtmI//1U+Fl3b5LI6aSKNvLeq7bl0ZhbgRHEPm6Re5gzcE7hIY7lXGbyAO+QqVh1BMn5grTD
o3COeI3LH3CGNnbeJNJ99Nkx/423u2+QNeOY/J2LI2a66jAUJE5zoD17Tz6KUbojUWweqwLbo1n0
vI6BnCX0dXr14GNgbH/pu32KGzL0srlSv5n37vjHCKCSXNYA/drYzwCuJmEqAQ7gx1qJM21+BN46
M2k+kV9dI8bf+KUVEWaNmPGN8+jeWaKR5KU0uXrkzWQlBIR14e0OwdFLfM73/1abC31g1+1vGdLO
I29hnBXroA6kxg4Fhlv9jX/bi3VrT4LSg+W5vlWzojGHh0UiKNisABquNo6V9ETpZxDHwuu8pwbo
qFTVCcgYtlH9nA6bCKlRjKXrtNfe48p7W1fKqvg/ael0tSgcTLStZlcCkG3Mx7vuE2NjYzG/vxNQ
1koWHIc+i8x90zxcVPsmo0U9RyYe6X9/FreCCaj2mcMZZiLhKhweouRRLIo1xb5sSWTma0qlNXvR
PkINYh1f+eePMrMUZua7LF6W1hc5CMTP6VIm8i+TYPsWDMFjtqhZblMSr9tB6xF5AmQrTx4MZk6n
CE/F4VNnrt4GF6ZaDMF5BMFMcU1cc9jhoSIAGQkVS26vFH8yDDf3j4ZcA6f4GU95M7jzMAISQ8gQ
EdImn9gsXH2mBnLpYPtFnX0OvUra7O5ku1S7Y1uBiw0ej0qsykympcZ5vjL8K4sA5/7VzkBZnR2Z
xYOqn0NKL48E0HAm9eUFgcb0WdPgpbIcfVM6wGPW1kJYc4jDz42Gx9PNOVieOZcAyLWZvPVVTejF
D/WxYAuTYiSujVMWFgGLbOVLQArgdVWee2UAmOvo+ufWR0Z1TMFxViWz0Lh2LHvPzuKJI8mkHhXH
BqGb/c/VcThh9NSCguWk79ZkPV8cZn4NyuCX4ZLKXpUwmjTFwaR0JakR0rNuegVoOklQNzte0yzL
pBAXJkul10cnqu/HQTaxEDjD1gsTT0qTcBhQV68P+c9Tr6Gm3sTySVerNLs6qvd4yRSI4GNJ1dha
zfUw4GmUU19RTpw8EmFS44Hj4fMtyWTR4IqGOkS04fhcZdfOfnLi6Quuz8mm0kMlx6SpuYUTPAuw
WTDC6/Uy38Ohui8RlaISpdyWc/MejgzpYonCzkQc6ZwEUPxbkdx0UJb/Zd1C9zQ3h5CtMMG83dKo
V3Ky26jxa0bymxj9Vyh5hGNsKMrUGJWfogv8cx/LC/YMJp9S0r0Dov19EqZU4Vf3nZypEzultfBo
YfMEu5E9+tcINdDfx/QBnttPTbTcFwukSYceOjsco/vlHlLwbVsdIQzfpl5tb7ji0VywPdCfoWvW
FA2RgVqtu85bLpf+fJwLSgPuO3b2bCYxjXqmpQ+RihMxoCXw5aRaQJ7zbgvJWdsM6nV7KK7nh3Dx
f9xh6MePSlkdoi0GewDQM6WEhL7ImxND1qzQMB22ssBR7UYz5xENyPNthyoAAOiOiplc71gMj1zK
3ZFI42NoegLC9/21W9J9boDQQo1Rd3N0bfVy7bRz8h9StmVYjCa221pD/RUG+9e8iUKW7+LhaAIj
mgXe9uf8Q97FbVg4/DqXJA3f935EO95KYnWKGM6XXsPlwiV/3TuWCLTu7eRlAr7BnbUxt/SImIaW
V9FYaB9n4TbbaI8M88kGDlQbzxP3SK6Em4Hf6y8wLrtPntCNNf8rWJ4mIgG3fZuk5QDdS3u3xjI5
UIWBS790mCJRty51C1ioT7r9mmu/XAy1y4jb2UAEr2pGb8xV2gFpaQ+KBPsE0BAF8R45wNKc6TXl
7uFk7lHcvwPfX6Xl28BVnX5Tys/wADAhJFLQ730TglAKvzNgnwzPXM+VpBqClq9sdl8+Ma9NSAf6
czuJeoRKSrDQTTYwlNZk5n5dSLKgt8DPRNLrZCy32zB476htWSEqadI8bQxBNU0Ux4JVO/0wa2oG
b7CWQqahXrhAQscfU8I82ark/fyWncCU21kF36E4qAVIwDdPXqCea3gAq0FPVFc4mEZeJOGAYK+E
mMDqXUS9owHA1QY7YvKNd1dyv0PSg1Atc1aASLxdrEyWmWbwv5ChDwnfOQV9BOv2IiaGPoL8VpPE
TRQaJrHdDxL2kS03kXU2EB53O6De0fNfw2aUWHG0W5xDZJap0g/1PeAPNuYD2uJzHIIn4LHwdf7n
/O2tYmjrwSAaaJxLrAqMiCem9Pg9xD1I75GAafDtx5Kl2DPwbIw7vGzGqFrDSPd9DrLWFw9NLrBf
h4cBQ1V0FKUUfPCNTmitTR2WunCQ2twrWpOnoxZA2Fi6wp4CghY/OgQE5svofP+tTCHvp2bjvLiv
SA5sCy5keuQWAA0Q5f0X/DSFOdY+tlV4/wlVKNCKFhWS0p52TZhRFftfhOaYP1OLWRAlsqBEeyVY
eAcjxfQLIGjI/hkb0bgYgB4g+/cJQCBwRdQa6hMnG3oOtvDVLzK5FVkbLRRYijIrVxhfeNO+89MV
kgyV/NxD3Vd856Rji5a6Gyix7l3/9GnftseizvmLEw1svPtmqvQpXI+/NPIJP+2vd8e9UvtBHQ03
pQtFbtEEGzaIErn4l8+2Rg3iOBtjvU5ZAUXymMvGqu7B0yHGw/tiOq61Eh2luGPnFMiPc0rJO9gV
UK9QbVp4is1ZtBB+RISgOlrCS37s5iTJbvN3NI/czf4B2vu/ELf+yCU8VX5pD3J1tk6nFotsALRW
6J5+3MiW/Lm5uugrhW5dIoOwxYr2yf7Ot+/kYvF3rjH20ZYaOcOrdZZu9nOQJfsJ0NGijJgFUonC
pcpIW3J1GeA+tas/BD4rg5zB8kvcLzP79xJ6Wy8fH5TMAOeXuaBRJIsz8FXHHtyhcSN4hTFp/WEg
88qaiAd/9cFSN/5SZ5XOwIEZMsdFGhAWUQ23DbGHvGYwr+RoZOYlbTtyO+rmv8gwHEZuNNZwCZ2U
J7OUPqPMn2xjre6fNJF3cYzeZS7HXQiNrrYk69k4MknXxCCgpuhDz+RFX/U9yE2HvdMAFKMMINmB
xuE2N6W1IoKgdzzMJbB2tP1gqzsSvq8NjRfBYoA2PbNtec+RVAvgChOYQO30noe+AyZ1Eo/uHqM2
GGRXYy6bF5nICdY73MmM1AdHiqPqeSrOXLcp905xnqWdR+kue6/rw0CnDXDy/8r+0dxUNhXXQJ/l
0aEcTHVPNgl05OiE5Qg2pyKnHVeYD2cxsewnNys03ds5kcHPzJk8LoipdKcrN7CfEQws3rCWqUG6
iLJc2XWaGOcqhX6heqvML2kkCusFMRKZvK7kkuNIBawmNDzm/g0rKRJfl5nsLnm5eSR9TCA20eSV
qKKya/cMF2n5YklQEcFxEOChyEkLVXwlYxwn+qD+FlR/sBc0taE2z6HY2k5H1rXFS+JHk5Irti9i
So6vvuNkukISHpcz4JAC4tHL68wwVud/k40E1rN2B1VaExKjoXg2LN9R7D/PwHqNLO6FFQC3qJPs
4fWlq6yJQ8wieGirA6rpiQC7Fke0EyBe6SLw9jNC8XsbkQ0N6eF3hlW+/3N2Mqq51qVoxy79lq4g
V8Yzct2LvB2c2oRM+LEgFkZCRQ0FxbhjOjkf27bknx7kJwxajRQuhJNKvf6Cq+y4J/k7i7VzTfYo
Z+jrrH4Wm2VCXt6OQ97bbhVutrQnqRahnsjE/GxSd7WcEheXc2PDUeneTFPfEQpr6Pnn6EpsGRHv
NFYzbRVAckraANYhEJbh52RtBeK0huc0G4sJu6/ADdm2vPFmoxlFfO3PM9XKN3k1QQ7LQq/K+NVl
oNt5bszQNDwlg9y1WEJhwHlP9JTFg7EkS6dpw9NV1nZHiFJQF5XnkSox17z1i+TvJRDmLOnqs4i9
BJ3ru2h5d3yfQW01lig01fH1qwBfFgw4G2MwgTTn/Nc5IvjpXaMr/2b2v0ZSnYsHKfCYkAjem9rK
pEfrtddNf0r0v8ERR6poEtV+vhvaXJUR0OmsHPoyLhMCGyXgkZ5YrHOE2tUS35KlA9xcciTsCpnj
smiPNNCaQ1oMUB3FqnB2x7TqasAZB9RBMGZlL6YDgP2aJB00t8QKrFrYDgYFPmswHGe1bYeqq6bv
eGIP8HcZMi0Yses5vDkeUxiGwdPZMvGXzRmbkpvUmJmAHJ85jFG5+fwKIxcDRLv1FPouyj7tCVbY
XClhP/zr8iFuU34GDJl9uX58PfG9lb5dlJFOneRy2VEVYKGnr4HfgqNAGvBcmgNVp68e1Dzyc6G/
ZCkdX63f81rShfNoEX6yfHjhA8XON54iXh202GWdMZGnk1vO2eR1epar1/w08DKvc+vWF/yqPEeZ
HoPHXZgEgf6FBKWzgJnEWK9lJ36epJb0SFOv3IB0U98wjEjhlClt+I+nixf97IbmG33QnVBnMV1A
o3nRW4TFLx8WvXRL3Qh+aXEogrH0EcaIL5vlncSBVqftvjq5abDuH+rcLdBwjGXrDquEgExxioVS
UuOa9IRyw22NMmc2V97saAPcnfM/lMSqEu5X6LcZLADUcqKzef2YQ1rCcmIJvZzNFkjjmBuBK8Xx
tEaLuoTDlFhtfngNRiYB02RyLePYtuyncgWAS2CM9MWGuMX6o5VKuNvut4xIJYCMkda47/+2Ki8c
vBBzXe6/OWg+/ygGo18gLk/ZqMt4pBmNxYaYomrQRBqSkjLaBKg1Mrdb/cf2XLAYwK+gUFzh1uj2
m5spnneYVInOz8FPiAmOswgcpjR7iVJt1xiU+PzD7tZfKZ/QUk9UGVBcp4sjQnaBdnlGYHNGwsQU
Rqd0d7R1i0XE5YLGsFZMQtp/TddyUioe+eYivb9wCvZU6RKePjQ6h8xpyjsb+2qS2jbxap8YGVt+
NSZfScqIHAubFBZsi5oA03D6Isw3jmfJvMg4o1TaDNYugWzp2aoT9pb1mQjw+TSDkD+k4tuY7efq
8trGayarUTzaPr6GPzdah6miTG3Ud8e69nQvNc1bqB/WycJbLWQX2VzLkxdGaFigf7be0TzVs+eh
YAD78fXClKDjvoIqPslqgXoBxbatLaoP6BAox+GDVcQsWQJEtKFloFntf0pHqwpTGTQkVoOjPmyb
IrcMP1IQF/YeuwdTHVuHcUI82TrcM34Wbr3ybex6OhyefeZDWE1MMi0E80asjdl8tU6QvQck6czQ
OXDU4Vlm1cBY5JD/HiWdATpeWAMYnWBUlPIldLw3wFRmhWYjtZVXt2G1ajR3GH7dgphd0nHcylpP
4wNJczIKzRbDrkIFkcMUU5IG3QcfcsP/JbGek8HPVL4sW0G6sICnbwlPc1241hKSxdr6xFOfGK5W
pQe0cSxD7cOYJa07dXrYB8VhI0/lfQPzUYg1rU7JmukHG2t0Fd7QPkISXIKUUfxNsppW8A6GwbwR
BGKc/JwZlncG0Hb7vdXPuoTbEfvD+2/UhNqfnF8jcUQolkxgRtXvNlfP2yU+76AKFvdORTTegAmO
pdQglvIK6JQC0dmsP/nDdu2A2vYGx7wsENwRlAo7srYd1v1NYxnJs3CygU2Su+HWprUc36DS7MK0
KAAtPUK2jCFfBBhpb0Npz29xUZIY8izlXY7dxefM2hr2K7nzj4DY+lgmDEhHKaUreO6QmU4AryXy
vEYFY9n9zMpKB4aXHT5vS8iB7WJ3R+BBOoC9ElEKY+mx7mgq9NOLVLsm1S8ceRP1aVRFayu/1RsU
Bn2fBex56WHEuUqcBGx01AdmX6oLv6G8dY/Nra7JztJM3TiGWBr8wrizIMnxlBxvq08uHMM9sKG7
q9anrAWtkyJa5NDUBbfZvhIe0jyV97KGaIvVgvDnN+hfDajpv6JQd0VFAo449+WXzBXEYwhiFpqx
eCNzgHWcWkjQGzvM8FVNiscnq8HJ4KjraW756p/DtfQgkVnYYVTLyfqGi31S9vEdyblx8ekSA3IS
G8Io5RefqZ9JFACQcNw3hXSz9Wt4Da3xIbzVB7YpCCik4SXaLXJoMK2OKKZyUSLvR5x8V3+Y6Qd3
ElkigwUnzRy2iB2KnDodiUF1E9V/Bo3+JvBFxkT3K+5QLm2Bbr8CEwAVogthz81Tp6a28rh3oosv
QU3L15ViGBd6v1KAwOgh1IHpy78EeKX9aUTWS8xneFK9YkUMoabpygDArRPAVei27ndSqkxQx7Ky
6vMM0NqjjNi0rmZFo4LE0jC+eNRzhDQTn9+V1cMzzntpvGfoC5prc/QhxCXDH4YNGNT/Ez8cM4dd
oxrklLJTUP0+Q06r8ygsdRK5LeDlnECNoezb+fVG53jGfZ8Cxodm+kjZ0fM5ko52Ps4FxyoGH4sQ
hrjFeu34vWCZj+BYrxNZzCmKjtlGfaVTelxUwxPEaAUc0ZKVzbYaorAq2DqhXrXSGbLSBK443iu8
SA5K1LffNqvyR4x+W1APR2pLa1QqtMpZDKKS+0G9s/smGEfAR0WMVMNMot+ejrLCaSI0KCRe1lDi
wgHXQkb5KC5bx+UGi+2gQBnSo98Hr95oG/ER78PduCkIW0Rk/Jcqi4vi6WQGeRUVGbjdYgaUYtrQ
uD8FQvE7rPjkEjwqtNO1t9j/14g1T1H+tyC+ge6oM138KR9CN0vxhf5mxK9+x6sHklLPjsVR5u1p
rX4dTCx8pFx45LY2fjsVKA1XRK4McCdm+AvRMChu8sZml6NZwB0L+VjyrZo9XLPx3tyn6/wrWSOB
CI8gHu1sK0sY+lh92m6CP5DIZtJDjfn68yv9S9R+mwgvPXNBwBLPzxUfgExcLRnfWdIiJ/rQSTe6
XgrKAxHIfI/jGun+BhyaQBdBYLtSH+gTQiS7ec9XEMwahUeSqjwXo8o828BMelXiUzlL5DuJUPbj
rZQiH6hh5vosXhHYeJaqng3eNRR7xEdm9SBSmfF+aWJK2umhsSOAzPwAYn56C/qxPuIbIBvCy/xn
nOmGRDMeK+RmzesrJeHjEcFv7sN53HfbPZIKJNzTVjSm/m1utwb7XwNnk2F2pQC79xyiT+h2vR+V
LFj0yPUuJwzMd82W9GFLdUtSFaqZDz0+BHdHcRsFFBn4GUbxWjLDzKESZybrrITTUynrNIw39fu8
v/pSgeaxENZBLqcMA6M+stGMPyXcOb2uStZt6F4snYIEK7FFnVODkEmoIM3Yr3pTtW91iuzqmcP/
lC5zJD/zavnClP4SgREFkTCxLbGaxLMGapsJJrmgE88aXYv+2REdepxtygtTqxBO444eHfN/LznA
dPGV/HS5C5yXomfxjRDzgjRiqaYbWdIesVD/+lNUU1Iy4laLSq7+Tlyjwy00Zu8r1EXPkbktUHCL
dEXjTE0CZ9KPqtoML/KXb8o9mSktUSHtCqzePZnLyZ0E2G9Squb73Cj1dJTpCZNqOthMtwSpYxHm
3+oBuov57auYO4LHu8i1dU4ACGiBUNaVMaM480MG4py9gDf6ootBALxf3SEEihcSyZ+pTyTyMdcR
XihOaNPR2iwXmSpZ5ngu0CdVqs7htv6e23q6g3gJQdeMD5eR/galrAj/BdCoNQZQr8wYe7PjFt7q
LFUwW1O4vVO1s86SfikjSst8aWVixQUIX3R3tfUXkXQhMDpeXQCJkp0iBrEQfvoVXOKBWUBwO3aG
ZR5ViJQUA52/CjBGbi6X0mpVFmvcVg4lttMTct61rOZwMyPWov1jtrd/26he2F/76dzao+R/e6O+
Ao94khoSi2JCk8hTtf8J1fEEtvC2nLALhA7d+Jz6/lLuQwnk9kv0AWqQt2JDs4FufqYE8hGr5onD
rfsvQFPUS72NBs/QrTcfZCU+7ho4qalxwtDO0j/41srz6cesllpeutxA+kxSTjy44JISdLtFWeVj
553mrW6gAJa4j3/+12WF64jWuZ/qbcy25pciXg8PSBeT1XsiPdpTxCTHrgyq/T74RRY68mjBTudT
KKS14pCF7hZU48tFAreeB4ICS+UpItR8H28jvOrsKaY3Y9p2dB1JdQuwk90vdEN6HgqrX0dcfpTf
IUdGMZVUXq3h50jToJPyvmIvhyH9+GZ/iDYM8y0gKFBkod/usPW0wsmCzyFQUzS3Gg67ScnfMAoU
V9WnU047h715TgTPZQLgGdyjPcu34gB7zoShSCj71YYoNGNfg+cGRmAhzBzDJ+UTk967F+BnqqEO
felN+Dgfk/6ijE9y+wt7/plVqhbtX30/zi6eMTftca8Sj3B6Gx6uHt37+3q2/7JIQgrsA7c9BKnu
EVfB1RxNv/7c0xlyTLH2dnHERMxBSY6ZQeCzwnjxPHMx+xTrmT+HnMeSAaw9/EUW1PaZP4NDGP19
s5e07dztb/Dz98V8XAEHBcBN21vxZNpHFs2gDDsMknvyG4ya+UReKMgYEXwKxGNBrW5/W0U4Khgx
nvhjdfJMEWmJZMj3f2rhpDtvnsYnQyGTMLLLKZtmfKOs7POGN17Y05YsU/8qBvimusFpfI7eTq1L
Bg7pND4PXUPC8o5HnZVbsPpudwCHdXYptXd1Ms5MzylY0XyPHR95D0VGioz8HjsB2FZIDrG6E/NH
C/ulAzAwaFmqiKhmLcSB/fxRVR5iPVhmcEEmSG1uvMU2/KAsfZWB7TCwO/g5hxm4BJkXB7ShEG8r
575sWoE+qMTc9x/GixEff7QYvyG2Hg3urmn867d0ZRE2B/GdgJY7cJzyYETgLXu2tUX1VphJRYrO
eFaPXC7KpK+6aVtt3QyNbL8C1mavIrokNyEuTPHeRq0Waf0Jq/bO2Q+OoapnzpZimBPVC9IiHZkx
XB1JyefzdEBOAvRBCqiS+3IaSaeSu0bkrleowpD1SRfkxUg+dPuhF+ju4jtOVOlyZD/50GH6TTGH
jhfss0gjP+vIm1rOLouxc/uhYjxTyS3gAyV5fKZBrpvOOh6aawcVmhjC3Qi2jASRSgdhRaydC9bO
G5/NyTs3sMyVI5AD9xQT8GreN/GQcheI7tL0gOUr6XnUJiAnztUOAxOczC1U3X0uIp3QQIf8AV7k
5TaxCdPToThpMtPiV3/CDpKvYNREsIRNGHXOc+WRbECjjX6l3mXD9YlukJ0dmizrU1RNiACOvvua
kOW7CQ8lZJRT8q9+uFLafuJDLj7K63mw63DYPOxvTcQ4uBiqeKOobC5IahcSWGwZzszi1McLGvFW
ZTeCbzC6V+a5WkqjhhMBA8AoDSILO+x1tdu6TcijCwNcPCMZlboHnpc6Ua2oOb2xp83AK54CQiGr
42yz2aC/weHb3cFRy4TTMoGrBmCjoMigHQYyDUVXE447EGKeZtPN4Kovq4N3BnwBP1ofJYjWyzGS
11WkZsx+FtC1iLZ5JpxhvvI4tTPc5NCa+oP16iH2PehJPM9tfCv/08Nz8yHtoEAkAKtcbHASaRwx
BWd3a7UHHprn2LjEOhCVs9tTeWGBQPC7PZRRhP9we9lYtlpKWl4mIS3uIum3r+9mlUbhg12SfveY
fG1IuN+SZz6V4TKtkvraxNljKlNNyoYvuJgf4hHztK3sVt1S1maOCPL0PwZuwPRmd6Rj93PPgmMe
oy4yRn1PtDG85u7r0E90w42iEsbWsWVbr3Z0U5ryBIEJBxsMvwgAXp4W1EycX1BbGJGgVrYliRol
SeYgaix2TMGKRLSnEJ0iYR7+8ifv8Hw6lGU4B3eRNEqLS9GO2RrjY5Q2jabkjIt+XcDVzFiOPk75
wDeSElgav7b/1+lkwumP6U868W3Yju98D3yEbzeoe5IzXv+iw5DLW2k7kJKSlqusv4/wEp17u9Kr
n3Wh3tpwSLKaXXG8ltnQonDtRsl7liO7HP7rrd4SYGZ00sk+p+UtSIlx4rSOejpr7IRwGXsGCvDy
QCswhBnDA2FQJNqzw/ag84fngNRSlyMkrMxI28QP9zOixnwfI+AcGwyistRdajw5puid1iwkD5tJ
yGiLJUUvH7Stgqcb7QW7GIYLcpT+lY5mDZIWhiRT3qtYaVlQqrKAhVWufaktW7UzF+tteTLqAI/r
lmcmaeVN/fzW79EGI7LRLjWyPU6/63eAfdVw95HCuLzm1Ps24C4xdcHw7rWvz4F7jALELdmsHv+X
7nLwWAqeBdKmg1se4Yka2gIAAP67tmBZ7CPK+KFl0Xn1jka0U899fEXFKZyfo3qmUKm5yBf1YOdU
alUJMrzJjTgUE6LA89rtkKoGCICTa6I2yrwDzYh8Ts6QOQVT0vLw7MaGtYTYdi6WdQ9f9KhMDLE6
fMyox/5+yrdVAQW3jC/8it84aAF3alQogceL47xpmHOh3suxbLmQXQoE0wOlXKSjEbzGybaF0mir
+JMTSOo9IDiI9Vi1+oVom5H+Hylz81MIJJuTS/vDddy9wHfXw7Qws9SoJCS88O1r+iPSRGaBrDYr
OpeYx/AA23y7u4HgtYx6oNHcSvLBAVj2O7EQHJwWpTpl5uqBXvhs7gatK1XaqqjFrgR+4wslz3yx
f1LeABbl4WT9RCCZGepXE1h36adGdpz5yxjBNW2cWZiDGc0xUAiK5cBlu39c4iLcLyWXfbFEhV4T
/8PNwzAYX2nBioo6kFc8oC0eGJ9vxp9M0YYo6juL5ADMy/ClZUg04K77nOHcvjxxSJWvQe0MzaNT
F04bXtifl8DWgwVneFgoBNXyYvlqraEZs2IbECly3b+4E//esF2kZRTCqOhZr5iUf0TZWu5RFXsJ
QLlUcomYmVp5CLDj+r7Fnj+bSb1FvjHhkiPki3mEGXh0REqribZVT8S04FtvtB8HGQw/Zp24qqrX
wkxziJs+8+iX9DTOaYXKq64SgUkmj2LKDqndBZ9BR/L04PWwvTNv9+rDK8mAvD/Obuk41xRT303s
sEZUP9HTjjffRvzA1wyqY0260SqYrospyeWoPm8WnYouAmjtYmXvu9HdqH1HI7ien5lH65IMpdX/
XozzyXjfc8O4tsMCyLbV6c/AfCoXfyF+alpg0sZsdtXKS8OIhDZ4tEDYwXt3vWYcazrYrol/sdd1
6w4BrkgtMc3h5unLUMmWghLUNL8FmeHjD8fnnJrtzU/wgVFoVrWPakPqY5gRp8/3wydhA9ARrkpS
fNMYCd/LSd2hlD8assPwbzB7X19k5RQ6nAJX7FeFZk3gmKkq652hkr2Qm4+IXkIZQQMnuKleHCNN
CjAUeDozTZFj3wiemuXOA+eUYm0AWnQMatY6tROKZS468GSvfShjU8d4xRAdrWW8wghpNZCXUNS1
z8XM+M7WekGm3urMh7SSmD5tQnE69axlooORq3IUL4yEyWnjlGqnjWoXRSN0DwZD69XPxvcpYK6S
jP1nreZPEBBTzyYva3R0npgpqygWIUXDkmjYOsRjC4mWtTDqcgS5QUhuzW6kJ43zHLLEBOc3cJG8
1Lo9hvkCW5Gn2wgPXcaWSHucq8qDZJwzfIzC685eUkHFefyasl33vGPTOVqgs5X6lRzkc4ece5wS
rMR9qZH+W21ZCfeCYG/9cm/fON22FeuoOXc/qXlIUQwcmO4BbSPsnqUm9lZVJExQjTYrwEIc074C
9cNKPQzcjdSnuhxlCjQJxQif7gPKTxV63NhVTga1H9Duxgl4MYGekYH+NbwhaHjLeBMFp3ffw8+N
TU318z2kPfxDUpfiUMmxJPfEsoPTryoy0R+LVdDi6KpnNOsKCC0MyN5ce2i2ckzq29vOVI3OqIQK
O+swdL5wG0yV+RN+203/YoNoKfwka7Vhqr/Q6Bi2YRoYdDuj450UHJ2OB9D4cDUXM7mKOBD32aLb
7wDe5/WFJJ1IV/xMXPel/jyNRMR+NlvenKPRy+R9MWfR0Oq5uZ3FQo2QSvi+Mhwv+530qpOyt7Kk
Y25BWxKbWIo13tdn5dqWKAvxPJ48Eo3O9UItR4150J6Us+Hkrw0A45Neh0/yNmHdpECfZZDfAWwE
5PXENlVi/IlcNzuToY335jJP+JecEuDwVSudz1DEjJUy9nteALh/5CL9/VQt54lB1C6jxX8mUBdb
esLD3erGipsipXxwmQfUyr0oFnI5vQVILTVNGUE3ryt4/bV+qSBTyHZzr2qrJWlpXLgG8eAYFtGQ
Uullzzc2oTup8ExQqaufR5K9KSgi3fu5YOkTOu1A9fXa/rw+7RYuoYSo1w2ZGKM+lcTKWlhd/noW
IabHUmzXkYpuh4KeMDtqlhxjzqW4u2VpG9txFpzewQXszP7vp2MGunJKMmikbPl6BPUZIRgZymR3
LJ9Dod2cV1bCH0CdxN1iLjEpP1NArV/x5RwfGB4C3unmkrr9dZpYY7ps7/+lXaBkuiRiXGrI6uwm
I7wv4JJSnw5n8VJvCDmM5CvezwwU0bEw08VDlnEg+JoYLkuI/zJHGdlJMIa0jsDb9xmQilEs2+kS
1f3+YntC+hOvBRhi5bb9rh1D7hSPtiryjLmhpWH/n9nkvdRYsQJ7wUMSzIw+WfHod9HskoyEP4/7
sFWDHGPiIBV7YjUWo4R+rpSUT+g47a2Hnu3HiuISl3SBeMttBCVQhVTj3Be1rpOU6+58imM0/SBm
c6d0a1y//ZYYuH1Nk21pKmctGW0NZdwazvhHdc1R7XMSvoOkxteNl/SLuaq4oQrrUF71KPWNMJfx
1sCybbrREQ4hCuBW15FzI3TG3jlGNr9TEC6rhjbtekCpfrhhPEuzSprHu3RRfixJI9SBOgZ7somn
dRhOOOPEGYBPFJGIt4wvXD3E98LVpFs6fy89cHXaRzJEJkgIx+S0lTEdEpTw1fO6bxSVwXHPumHo
Umhwro+CbTknmon0zCX9z9zrn8vswI3Nlr4ZivVfHcVgzmcq1jePFM1846fogJUHx8+8e571Po+Z
UdoeMycpwdXsie6P4HLQQIQG/TzLK73zWhNwhVjePMYnuxbSO4Ies7mi2ZFeSNw/uk6Nxtf8QAQa
nsS0G0iiuq011FCcvhOi1yExx1YaF8v/7ZXD6BPaTiGru6JAzSgrJkz+IcDDutJgaPHPF3LSfPWj
4bsR3rfyWzCfRu3n4K1nVzXk+1yZkGhCJ1VdR1h2+fEXlo6pS0+nobtnrHJ3+U/w9yrV85bru5Ax
BoFDehNYBs8P3gzHLr+7Q4JOa2wrDwGPgyzonQPAoqSxVmRTuTHcXiB9GxwjwQD+ueYwtQWxUU6O
GtWsLqzgeyiTuQUCuDum2L2imbwK46ndWg0HgmcGX4p7wE9VY7Mg528lPs1iyBVAh39LRmOyQ3Ah
mfcaRev4gGpEZu1C8eynZyQDZ4RfXwn3VKtbwLIovw2kUqUz0OW7NczqdnPM6A4Qw8YfViMnFSGo
dOFZx07cZDSH6i1qhhLAVr473ic8Cdd/5fBaed0trry4m+m+D8NW/ElljKasU9etzPL2EdDxCT71
2DdyULokdqMg7DsnjexnzXNAV/dmwc7R6RKxQzp6ANL2GQvQrZ2D3k5E1pBwHioCnWpndj4hh7kQ
UssEeyrlIjAt3BfrMNeu8djTI5Vu0XyvJRtEY2R9UR9TEGbgCVb0hX44RA5pE8YaSJw7nzaUYLQN
Qx1dvyBM75d9YgXU+CMdyuftvD2obzE2UhLrUi6+J2B9yzyJxeI/+7GcJaJthJpLNbA3xKhH5la1
Hps+fcwkTP74jessaXH6p+oElMuUy/XlFAZvCGR1iMhH/YmJyDVmZEjKvUmdf3HJa3vK3uZdDYoi
yF9SfG1GLMZqyfya+wd36ngoc+V90kkmTbGBUS88pKHYiquCzB6HN+8/VM75bgTzQCGsspgoUbw1
pc2DsQXLSx/IL1/9ajNStg7ye98tZR7vzOYEtqj/HEL+pDjsgz9m687d2RqBFLvZhwuxHcLptuge
EYEZ8SM9ZUDvDK6sh8M5h04M4F4BW8ismWCLXrvkMPNmDow9AlxlmKnA0TQkTjHlf2Rf7C1loC4+
8rYazyXKJ5gjd5rqvoJIq87mZzFHoI4yaVGONkk/ZJZ79lOZNBMBEF+3aLzZa4slPs3AfZ9J/4/i
9X+ziJ3Wt50eskusmbbikluur3RudEKvmVNoELjcBqAZRgjvO6DQBQ0Flw0qlc6RHjx0Ok2oT7pr
zmFtgzT0dQ+3HhW4sEtWACD+Yt1p3ItyblH36NlzXYWzE+1yV/U8N7OQ5n3jhrW1P26Kz6sA19OK
WwDSrnxmBFBx5SGngpq6/IWwFN0K+Yl0UucxDZkWbT6La3x3xaNInh3ZR0q5R5dx8TngSO2AKt8u
MblMf0IOedlU7lKCJW8d1amOf4dozcfBpizDNhLf5rIhUmbt2FLNdThejVLdiSyrWEf9HfSaZec/
JLBBMZjEM14tYm0ysi+INB0ttXuFVwm2fKk6CLkswR9UjLxCA9CHNZjV44WywE+/GCQwZAqGEvMd
hnf3KiDwsGP8r1zFnD5xw481LyTSoQje7eh4S904mSWQFTCGPXhIgbzcW56EotpRWPKhr/1zJrYj
5M2tsKLTRvLrzhdR3gK3yRTRPc7oRRrUbJ/rojhOOwaRS7V8uFGNu1B+aU/kIDjz8vZV6BdzvZDt
+m94/7kCoDZc8dUk9oEHw1LAYxhhWuzALnNLUUZ6dZK0dG4qfYNcXJaV575uonPt2pLKbqlLk0LB
eJdp5qGU64DVef4D48DCVwAc78FiTy3MomLi7/NkNofVcCfwbZCHA0MHiJLeYJUeDkHX+m7EPn1z
bp/lmmAzArWt+pxg6U0t8R11tmFSMEfz/TL9qtKnDis6fOn4w7fEuaup44fzVzKmfVbt3dgUT9mV
7t/03nyGBw5vOP+JeqKT00InqO2Q11Aprtr2lmOd8o8/9LO5PfVOKK233NckKht9tves7Dh/dzEs
Rix4f0xi3ekvR0IR07pmkT1t+y1Qadi8aevbdlBqnmkf51LWzmH+4Eq7PA3FqgOC+Uo2e3iSJPA+
tRmB55MTTXxvHnwwlWU9SK05ScVVHHRsV7J+SmOo+TJAr6u2ddLu0OnvOeApAh2DGcaDWWArNdU+
ZLDt+BPoM+3gtROtbPboEx0NmM2e2W+4ERQhQ3tjBHGIzGOQF8qcSZ1O5SOVPgPXQYRGXgBiOtu9
GiGP4n+ltq6voavgiq8yHXvOAoNH2mlWr6lFontaaH3BDJaobStloODECPEDvgG2ZAbpBxYt92r+
+hkYZgtoXh3yGrBopW9DyrQ43jhN4IHJ523KNcEc2NEcib6kr7JCzDYJrCHnXn+E7Q4/HuOb0rpL
6+dKl0HXOpbpxU3ulXW3NIZc2XVSS4+8s3Q3cIcyLDTIIlcO6uUvvT5YiKf5baYHw6Zv7ZsccsTJ
QJ2k7haqTanOLc0dzOrp44SDy9mUWQc6Q9BKFEbP2YX/DZWAI7AJpt8a3jNvlcOVYfzGMW1KL0jq
QG8SpozYDBwz8Ph/7tsRKi35SKSSqAKFURLJL9Qfac9vhi56M7CFRQm731wZQ016D0IsNSs4KMfr
gcaLLQ5bPfhC5HT4RosKtdSeXaf4gwq8UVfP5Zx91/QW9zEr61BI2htgiv/em18/wMhrRTNt3S5m
vK2ecbMyzfhgivgaYV2p2uFbl582slmgLFp54PYb52ppG8CF6NNVttWzD25wh4XWw577a3abPgW5
dlR7y1Vj+r5wyqPC+uVqnl22Z05rSU4J/UPqMY351bW0S04+jDbmYZNu+deq8BUsHkE3fwddY/eO
iFOrmTgoznUJtPB0k1hK4qGqw7gcuTt9a6Wmojp7j943FfYggZ/ll4+GZdNezpJB1/WlCl9HbsLM
5NXgpzH2Cxe9sn/2QCK1O4h2W+i/5ewJZC/IQ3wvbxmn0pM27Ws4/f2VSIgWoKaQfELIa995W+b4
stB0VSYQZtPaiQCm3+pnBJc2O2DYE3mHailyyBOxoD11ZLQYDBWBwAjW7njfR5EpkEucOFayeHhD
jL8VuoeJxwzSP4vhN0qxY/D0XrKiwGXx2hNxaPSr0nKCRBpYJUHOldJUIp7pEpzBMi/asy4yx9Vb
lQ3W1U+3YrZLXRnK8N0qUGieTkXmXzsM8gj+1t1149HE3bz22L7kvhz/3DT2jK9AjmYERrvgcjrt
8NzNAzfVtltRjwStCNIXpSxBnb3ZgtE2H6zEWF/zLX94g+npCPrjdpvb3weMPcQx3N2YCBP9zhDJ
lyU9B0I3QYWnAWfSAM/VCYXTPi4O4R3TPXPTm+2bg3dAU40uNeSC4IvXuPrni4NjiTlRgpVBGQls
YplGMSDBH5Pl0Fr7VIw+pfCneKqg4VcPMHFK/C0U/+VYeFT6Kfl07CgvHWqFJhZlBHLxQ+8SlIb9
suKVYaCyPuXbmEzTm5yIWIHwvcAU2wvkD5PDvVMbsFMaLGa4yU7hN6ucKY2yf1318B/Kiu5foeFe
8yykDi2baTtJgVg8yumvvysMwTU5ulqemDnVW7djWbw8cvGo0ZDOrAL75GLGeXr3KbRa/eGfsf2f
XB0bapkV41MBanJPuJwxRJ5dsCSRwymsOiuE0tkiLdsUNI/Rx1ayikX5k6B4J6VXNaHd5EIF69Mt
aoe4bEB5jC9ClHtrscSrUFKj1N3qv0xZM1ZTDm/h9HvZPJe1w1Ng/eB/pgF4xgT2ZcWdw2yprAOw
Fa1eLdemxCDvhFDSuXsefDKehxML7kW075jlQRU2Hv6/18X7K6l4OVQQ+vRJCu6gYA1sfRzaolyC
fIJta3Z4EJYLw4hHlRBtgGg74SqkeeO3+g8QsiyBLYOpA67MBG0x0QXfU4xrn7CPtiuUbZslMyFD
jdXdzd13+ULebDNFmVJbStY7YiRtkHz1+G75FAvLn2juM1vyoXyy1iTW/63TN870T5Vh7DhDMiWQ
inWsK95KwmXt8g77D8/PeHCMl/+BlAQH+6M6qMHWa8kZBGg7A/udkOtBA+pG1WuXW38qqJBj3flm
518gCDTESPfy35PGtsV8/V1t3iZO/16D04rYgbsklSzntPDNQQydVYBOGQGtFPxQWZn1VKywVJ5/
wxXBwiNolS4q+YCJoiP/h5+j87LX8EUgsIU2ppWgq+sLLm7J+GGspHc4y4p4rwkfqPbe9hfjnGt7
7xl3otCpZt3h1Ebp/v+2phoZWCxE2GtysVdUN2PXO7cksHXoDfiSmoRU11quknj1bX31hyuYGdjm
MWeFeVqwQgTDJbAC5opY49p5cADx5qv/tSepwZ5SvaMqY5CmaRc13LgucueTk5pDS1aNEWZTdpcy
TV9rIbr3wo8EiysctzDhIKCkmKiAzYJlIq4fqycBRYstKJdleYZR6RWtpO0frHE9gFak4SRYSmKL
JlvH3wVJ34pu3zlvwGQDhfgeDa9sQh0ezjIWVHumAKSmbTj52OaYgEVW4racs/kSk3+qC/S4psVg
M0MoHsMhrMlsAFUSQfMbM7zUhJytVljPq972tvdsealrT7Abz1geFEYK+4ySRyrlM2THADPdOTxj
8ZLvLac57S8F3iy9EBjyBI6cKSik+1AM/dQGs2a6seec+7LodhK2SG2akNbqZ62HAtcEtEeqJ3Fj
OHz1zZEYEgYsYmLQpKQHK7c9gKuvZ6YJjtNyWYW10bEDjJfpCXOFnv0xd/8ocSbFWfgSOt3ntgLF
8VtGUWUhox87cf7bhrEwf5R4soszzMjTczGDbDLwbQnZq0EaOnkDJwXKPh7hsqcHOn+Oy3n1Wr9P
GRXwD5oiN5xDNwpEjdqAHk8l3lOExK6xQV+bMnQm1QDTgoDZSAzdIMX7zGfUvzdPLkPgd9dS5AGj
UEkHlemnEqkBaLG3fSxuN+smEwgWowLFdAXfo2Z57mLXl/cTWksReKhFgpNvim9LLWXdeTsvvckf
SZbtdjrGUktutM5zoJwbgmQUa9ZMgkpB/b7HwYKUFV6sPSRwcn8PBjPlEi5TFw7yZSoI3hU30h6/
MU8cYljr2o/yc9gP55jLvq+xWV7lLlvNyLOeEEvKJBz25T1tiOJ3+elub5FGH3UJkv0332s6qzOs
Szo0oVwLtfRR2P1gIxL+fEkbWmemmQDS+w4SX0j51hiA0hmuuhxj3N25356smoQQJ7robVAgpTgy
PcOSOIrSDJZh30NjUAGH3NqYGyT2TaUYwHX+kH4RWVa1lzdGGkYATWqVMso6ZCNpgctww7j08gvi
P3gM1qHdzK8Jl6EF/bboiYNYW1T3Av/hVRr5Qn81Xk9jWMRcOvw3csnnXneocUyVy50jlD970hmM
F421q0veHG+G4r9udLDia1srR/Mz9v2wG4qlhgoS0ADOqBYL2aA5f551H+HasIjyxG1Ki4mH60Is
eraAGFffb8hiMU5zlMYk7HG4ePuLTvOY/EYv4oLvzHkEJUIni6+5kEomLvH6RI2akzXgyQJs9gwN
0hJa5trytbqwDtlSJfvsVwcooSJPWjhrosVFYjg2KhDFjbZvjfeb1ZUtThZ6H+hfeWCUe4W57crO
MO0U0hBZyhdJuHou88W6Pqtz41cp++TNBpv8MfMnro5c3Agtv1PP8pxLFLiCsfpC87yXARc4YPgk
gARvgrLVuhLXGau7ChAbdkgaKoqwizCA6frPkysQsQQEUnmBjvBAtcXL5qZVtrHNYeyvT7MBU2AX
rYbyB00KOx/NQkXtXBGb5An9pNnZA9lXU5k0qs8AnXGSlV/+xqE18t57+9gdXzaFKcNBwW/e/mnp
L8JtSu9QVU0C3Vg5gOzdQDfsEU8QXIqjssDk89H7bqry6IwEXNtk7PQwR+b4PNjWTwedG0HXmejE
ymZOWdztqOLUYKMAMJCFayDioIVX5b1Bi3qtTai0gKucSQRez1yyfY5575ArmCn//DNp1atSQ1rF
6zkuKjW1TL/x2js208YKXHHFY7yqNUGiqYIck2qwmeWWzlB9kgmBiDG775s5sCOJ4lgEwb0ljD+z
DC1vfakKunGAhWW56a2Xbzekfg61h5gA+nQmC9UmB2GKkXDoWBICvmd2VdqeVD5rGQn6QQm3k6wC
JUhqh/I6MCdSUVjVBYHsMcVQyW+HDhp0Qj85A6LqXPjj/9tB9waEqPiER3sySm2BPOsBwOEf0w8A
mAv13A1v1dI1sk6LgUnUAI8Y33E8kpwDiI/LuWTwtYgaR1MPklJbpYMHorcF8UCp9Zev6wb2tLi/
VVc1siLfTU49csUdRIQCCECg7Ul7BW5D7qitURqC87ItPVUSqL1dghAJUMgZioL+sQQBY83zMGcD
azRRJgiczB7LAknvMGiXutlDIh8ocBgfTcONryqBuCGTo3QDFxXbhlhdQRH+7HpVGtaIokH4bBHm
q1D47xkqkiOnqWsb7wiYVwZ9hnCx8E8WbpJ5ev01+qV+gutMc/wRbxrHW+zy3wj/+xnjVZh1ztnJ
mx2TJMnYqlHlv6vYGMpYBGSRo2R7Nf5PxRDMPhjuVeSGM6oyY5IHgZ46pRsOab8+YIKEjTUYiH7Y
DlMXjxxBJrXRdE/aXda0GyzSjR5o2HZr98OC8P8GEIy4UOXGOOnQWgRBnUjGTWdVESMPZocfZrVV
yPqdBshcOORGIOP5QCD2koWu1abZ3Hn9OO1eTWLkQB2Y/sfJO8uWnCCpg+AF5nNPBUQeOVvieY8L
rcXbVIDgoC/4zGmH456Doxeynw9h6LY/VXH+gELWGbOrUeTb72ISvu37IN66Oj4m7q+MTEDRKQYB
z9+DU2uCVS4zfYf2M1AE9Z9s9PfdwgQRT6ZLIipYp7c24DNdbQgYtOua933LyzU33NGWz+RytVkX
CTR9bKKK7vLYO+cAIXugOpAkS/35ES9GYQyHDa45Om2NpgOmVNlTNEItt/WXgQioxAQUlQP/ZQOs
aRNAXx3NfSs9luOhNCuW+WTsE6mpaEYgxFWuN7R4WRClUwf3kpWzkNeKokkAaXgK22o8nvHzdMmH
7Vgb5T1yC9VAmCTaCWpmL8um4Hy3X2JnuTI+UOFM8ZuO3s/Fcbuj86IooxJx3zTv0bh6opefWZ7l
z3m2VTy8jjBxo7HVUe6FtWSXabWBgUnDp4pWVkjK6ZquLOggA966O08GkP2U5uEPNgvneZ1cJTVp
+zr+GWsUp+pakJHzDl8PneflXWfZlOyQmS4Bh9GkCd/MLQIqqLeigg0XX62CMzTfuAx6/PW/fkfN
eoAf1Al2LUsC+fz3TX+fEApQ8fRpoqCBKv38vfwM2QZe3GfcPiaIyHQsIGYYdJzC+V8fauLBHXC4
0vsWUTWYvu+Hvz08lRNz8slZlc80J9vHi9sNSrVK6PrNMK9ZFNRsEC4DPfJ4mTOnKUi8ox4VFPHr
YvDinCbi4DswcUtUQn283+CTsqyjgGdNnzv+1IggKKKtfrhM0ty28H32h3R/1esNr8kpLkJZ2MAf
qC4pe072FfEgqw0BHlptgOpmBEbmCsDbB9277X3EHRH5Bj2uuxVqhl71D0mEhjwRlhH9Q6xyLCvX
rJhpDAnQRcKx7ohJ7XmwNXfCknwq5ocBpEtS1Alkahk1x66mRekRE642ZSs1qRH8krPHIVOFOW7b
iC3sDL/oLQNFK3W03DMdf6d0uvrOEL0+eQTM1OepMTzK5to4tJqus+bxvpWazNcbp6gkG2jaDEAd
o++fnDWNrpulT4YLzmaPCCNWG6cPVvYp/XYOkThzhzZk/zYBknvser5i/Y4B5YIksLWPjHlBstGZ
CoIeZ9weag6URlCfg/i80PNtqE2hX6XpSdIYBzV1mZCIkQyrWZm2AEJPcTNLdxgxu6UdozpKTr+e
cgphPCBb75rSaTHUrOTX9Qnths6iTKpFYT7Ge6QfL9JussJqk9kLgyKPIiYFAc3v56LMp1MGhv3b
JOXr6ewgsIWbl1tu9gNhWJEVcasqjehgsXcAmXHjhtBLVqRfM476yGs2oM3ub1AJXcRPnSUA232a
48/YcGXp6dehBvAbRpEifLSUpfeyb+bfDSSmUSk6IY22jxj7MKt+jeAf0qUtUmIrBZ/zks+LDeT8
BWNv/ZqkhcrbUT17tzKY9YlMcwamZzpJ7DmOSnBU/WQa+pNA6wN35Bt5Z8GdOalBLqbObhrdDSV1
sCqNYAUVOraQGOd/oxlkRWMI7+FxTsOYLFv3zXwBddis1oFRe692NP0C0wtL2+UDlIIiK1X/AvD5
tgoOpReo8TzdX26nSmyUcgy6U6KdGONk6rC/MHVKy5PdAOW7DWK3rfP2aNNhWZ8HfU14MEtxFAOV
qJtG5rl8Wz1w1+TFk6B+BHGbwwLwwkUrYyugPhdg3/JEub+hsWWHfZ0eSbpi6MRv2XT2ODYsPrh0
tj2rqlko+DD8PbhGXI4I4WQ0BYVfvGyGlYMozkM/4GzB+NOvmi62KMtY311Q1JMFq/rmcSWt1lk3
muQNRdfVUB172Wg2H6UXDXweiKv4mMamgcrAh/njQjrkcNPNjIiff7/Uy8ENTAMZGVGH957uxg5H
eMEjg/jwEa8T8PPhomapYJU2aVibH68mrxp3Y+5U/g+W6WTYOT0vIFjUzKXkgAK0p3tztXMr7ser
gj8WPJEK9anXD/tPZ4BjhGvUypDkJb+HZwlSLQY/AU5+wM/iX5RP4JWvdjt5SDajn1TeIfRkcyf4
755Ow8oXsEATtCQNt72ObG1l5rJ+B7rmGcorPJqz+sDC7mSLW1uI+4ORNxWAFcn9Mf0n1l2paLB8
HgUFY88XgUbOemLbYB4LKZ7l1jQaZHAVUvlEk2NXKC8DOs37gB5WIEBITvX5K9F92XgRlvWEQgVF
tCJh/3/dKf+/5gYBRrglVww99mGLxxlNW4GbHs6lncQ67/LG8Gh1TLPEyrM9gvYBS9jVhMEICOq0
uYMVj2aEA5aiFX9XshXy1mO4r7dvnA2p3MngIRRlrwBdzgIhSFaM8idmaHSZuGaX+t4xfJCbwy5Q
IwpELzA2tBDCzMAmIVfhAH1WWYp0ig4+PUWAD8ZA6OSwl+F9UFx4A5F/hL96HJ8uToGgUL0uj0ZS
7Vi+MBPtPYgXBJpC2w4ybxjIHCqCfa0N28keVcb8RxEcdDNtmsKgzGSS6uhZa6c/ufHtEtxBg52Z
xzXEXtFnVfX3tnEdx2WYqvfzZeBvxyf6FUUXouQBssQ5ag34x59T35MSnBplSROKkGuNCJRRkk3h
ReJbo49Mv124wg0Xxhr+Bdl/FY07Jt6PQumazhdSGmMVxdK9xYnAZZ5NV6Rtl5nYEG7ojXy0PmwU
8kbOIkQKKbe0s3schuNnCy43SYnLn2R95hYoOI1iVpZCCqOKKZeOKi363h75MpwQ54nKLRcyQhXX
xf8Vge0XdLBdwXZVgUNRQSpfFeECyqt5gGBJo4un6KH5I+70utQBoMQdE6oa6ljA+lgssdzV+/Y2
Ll/e6+h2VrK+4VQ7DbAIFrFFXINgG0DvLSrJMWQgofI7zK7cSunP0U+h7DfVbzt6wcbEFLE7Iv8f
xr7OFtJU7Vlcy2kIRIf8t/L3lGYcTE3ICUP8zuPhCC3TIkS20mJEszo1EMz6qtM8v9RbCoq/eQ85
HjLQ8vSmkcsTQI5G6vghzyFotryVb9MKHhtdqC2xf4T+AToUKIDU8a1Iky7echsKgCBEzNa0qK8F
oFDoyY1fZW4Tq4JBlE/VxMhMjRHzhSqBGnT8lYlh11VPRzylJmvgXvQ2btGNIlzGqSrd5JS3Bqs7
oCRNRn/wH/SSb/bUbRus1n8OUZOC+RexJYjU6QS00tZW3ik8hSYzNbsCegkI0LqYXOkndM8QPpM9
WrApSNKINSFokVNqjbb4KpyIT2g1kjaxAP8s90UJPn1SDQdvb8QqvLWtnFOpPMB9ormS83GkAapr
Jdq3ZE8/dAaG7vu7mC36orF8ijEM2gemROZGu+HSd009FX9J3B8Cv7W+oLMa5Qnnk3Fd7sTCI9YE
QQaRpUvnbV76ozOaOSvgy+5FgNwFBddgzDw8WKwvMuvJoBJDZWGZqwF1Tm4KHyYkMuFkA+hOF3T/
BqapYWHO70+7nqGrgu0Zag89UqOB3I0qwXjv8VX/5MN/sr4I6b3FdDmRF6iNhf4WfPV+J1/32i4Z
ZWnjuIXobxmLUb/v5P89Hyr8A7ibuRIQmx0zjy/tYPvgUFR47MKJS8ubIkSARVWVR20BqgXUzVws
xjH8CHuy1r8KfUNDEuIQeaz6agRB4FNz9hW/wyr6aHBqyabFJW7mi/uajWe16VVYXvWnMxYOmhku
ofKilH9gcXFya03L0sMq09WBAV84yG8+9KUhG2OcVkGARKmrUKrQK1Fl7g+r/h9rIq6PopxZ/I3e
5nZ3f6ngPl5Gjsnpw5GPjJP5Wzrq090HsP+eyZyfD9bd02X373r8ho+fSf0woZtw/h+XVc3pQ3iW
FYejXZfv/UbQCafu0+B5p2KO4rTVLHXrw53Zmjt7XbudNIzGceQDx2qrvvdhjt3wCMV3eLOZW4RH
RKGAd49/4u1C4R8oA+mO/rDF9C5jONSXmvBDR0f01r8ndgoX85ekXnRMCwNEAXnEM9FwZyaEUoxt
vRX9fulfvouE/V6BUckJ/yyPEz75/Sd4EyD2/zlARukXnWD3idC2FPExw6Grqm37Uy2mbscLdrLU
cG/zRlz27n1Pm/QG1opgYJRYGEJQ7ekLd3VAp8/ryfLaOLoKK+/27ggZPdKwE4g5LYS0v0/tLK76
FqcPBy7WJlVnG5P0p8uwOAYCog4qUL2FBsQh3CtZe0oYirmlkJ28Nm2/MPityiVY4PEmLGbQg/FK
Xuy4P3pOknMXMiBSwcMbjTjBVM/RoNCmQV5baesaOkDnWcIAASCpQ3F4L3lzbL8Ajmgjf7Q/EqtR
vpsHXYEIytl4/3EzQ3OvvqBxynRpT8mOE2EGLgLAwasBVEUDih0N+fD4OjyAwQn6IOiES5lsSVRc
0ZSeqU0+lCEuUFS9voj12ZEEdGsynlW6ECJlKfgQmiE0fIvmVWlrAFyYhwTWrtd+E70cs1ou85Ky
0/N1kxQk5I32XShDPO4PApxAjLrbct53HaAJfvRzwK60AF+UfIE7QLn9MCxs+Of0g4bgP20+YoLt
9PygBSiyQajTarwnYGfkiEzg4xVShhHBpcfZLP5HL/T/5u8M9xDA3IOY3AUBr70JaTjGwAtfHXfq
uqnOf+8w8AdO2qCisKbcq05gdShFEmgqO+6D/MwHE3rs052t7bDf8bGeDlosPAQSf8muf6E8iJeb
yRWNQcUh0hojT/QU5vwI8EtWMWDF+zxMDP50bZFvx7JrTPpALZvweSrZz7dsYR6sbjDdPYjMfv4y
l3gRcTP7J8BAavxnNrLnXaeyOQ5xB38/NMa/wEOS5XuYPQVseu1nGqyuAdLVRx/S49scx23RVJSk
1dYBw5+OsOZXhA2n/hxdzH3Sn4nTNugzemjylsR/Yshqbkl17DjvtChIaetsGSEM1Le9Um5hSl3F
iZTMUsrXRVCAXv8Oy+AihFqtKgttSS4ppPQm3+GyUVyHhJJA7rLCy2NgkQRibBprTpMHovsK02Co
MU9CeAU0i0Gfifvq/+jj2OAOuRrYRlEqEPGSBRnCe5ie1AIKiTr3mCdbak7NRIr0Rl5iJTXOGbaR
9CR2IsZDHm7jFIL+AzGBuTHq+zpA7MTY6cNo5EjVGJFmlyBnJi/KChnaww7uBa8vhJ76mFMf3Hiq
HYIc97ZrgzQdUJLNMEq5+YuvZOv2GZL1aOE2bGfdCex/9PIkEf4t1jH1+55ywp1QabCSGDzMM+PK
xQ4+TZGs8q6+JD2s/HudJdvdmjlkmowZZCK+83c4vzWlEveiZaInnW+eWVT+f1asMAURMg8ccD/4
1qmm4hf7vcYwKQhQNXmBnCH5FWMPyvXX1C1a/EsWy/Xos/M2xuVCAC+KUnaKOt6CfD2jmklLz/af
CFwuCQO0ImdSmWHI2beWAXnZuTDK9PSlw8vkcJhG9uACwnEdsdP1tTcj26m8UQ1Z/7Ja38dgibay
6NwhwMqhko7aI0FD5n+wsT7IqVfqTQ1j4eapRXFiQwsx1meQoBVz9VRZNhHs3ZErivLo5nej5bo/
GvhXA0AnuAoVNUjd7jlhBV9VtVwl+giIFWFqscuF6JIFn7ZwDJtI4dTpq0PjoCwF4qSiRArM0KNV
9QvuX+/fWbACnZOtk3d+Ztsvca8p84hVdlxO2dq5XHJ+H6UHY2qOnZEeRSuS4caUC3QLRAJwDAJ7
HksoWwa1rOsUXji1+k1TOztqWeGoZzg9MM0QyYFOoe3VYCntAWf7yYKKjp1MWnBLMjtJwrET2hjm
rMwseyuzGgXoQDXkg2Kr6EXxW4t9ePRcoT25blm7L+/hghLGlhWQmSkc9suk3m5lKibZReGoXaaw
rUlkpupzXviqeqZNXiWhGCD23plYfIGGhzy79hn+3n9pgiQPZRJP3Z1TB1KmQT7GDsS9o7iZ5Dx6
hzznoTpfff19a06+xYdlx/ciQbJsdm8ganvthoV65zZCaTJBn805VoGqbsICa+ll4PSTiKAEALa0
XIu7RaPo9xDk8eJWCW9lZvjl4Vfppw7PG+WdKxWTJEa1zkMUH4IhH9rXRqqXkGzLxfVQsfK9ZieX
rEytZyLPcWikPL8f8sbaH8TtiwEaoZJv4oIhx1ytXSwCpVspNjYkCi5eQHdvb0T/0WIQgJyFAJiC
Oj/GcPkbz7bUmE9ry7zKcVLzO8ZN8BVsPUVU8seJtLebMaWSDpeCAgwNt0H3TvFgMGGdlSOsrQqD
VfCiGjNUet3KTdLCjeBAl8EMu0GY6LWuzNy6JLH0UK91SMTP/h52dbpO8HUQJeuk/Ukm6e8ftY2M
Gqt9eHHvOgKv7QBDEXW6WSpaoib8ZmpLfmVbVEDku3TxTrMbprFGyWjcLMafRGlOpKpCBOkAfrnq
+5XkmfrmnKIRI3oAtuaDT792AjxTcIBXUdsCEWNdGB3CKf+HcTnqcgKJb4UaO7HBNvk5whRtx5zx
kmhJ0eVEGz3U9uYCE0uoN8CWFYvx5psi09gCTO/xJ4muT7YyRfHahB2RdJ40uyTH+CEvBPJoJDT+
oBJ46pVWL3Aun3Y4mA891qXL2YwsfLybO+zFdXhZmMB5CT3WVWKaplzYDe6cZec2mgP10CO9aQBm
rWCUMqLc4HDn4QuAgI2/h0+4lndwLBWYHVqgjaKBRYPCNKDZ3c4DakTmuHZKdjKXZTPUcIOv/EXa
WWh9nlZcCAqUk0XR0J8MsZ+pNPjmM9vIiB6WYmU9xMWc4ElpYHy2FHylz1JPaz5eIpUplur0YhxX
YwuLrwdJldFtKbrnN3orgL7wlOMZ/5pp2MWR/7NyjTO4T7VRRt+1Xine88/B1xuDQpxBfr7jylDc
DZqGkgVm41qul0B2HBH9CAvzzU+zoFcgAFYDZU0PUcWvPJwzsafZu8XybMVpOrGd/tUqBPi9C2a6
qfwTC//2xOV2JPluui63L5T5wy/FR+J3QROBEdCAcL0/ULiq76Uatvip74rYYPmdYZ9xkPHpQ2YC
ZFuYLhuYKGFyDbnqX60xxHBq+aUMYn/Swig7ZgEa90+W7zafNd4SY4dV6P/LVau7oT3N8kUtt5DW
yniAZBv/JnwxpZFLaKUXxtKMZPqKcc6VzchXM7LfaK7kggN9dgThkKcXXiMCTuMo3uPvd+8xsy5d
tLTtdZX6S2mpVgNw3zGOn1U/5CpI0V3tyKProIM/iwFTkqyV/ZFHfY6F5+dsXBJ0NMw9ebAIWwSk
rps62Bkq3bh4c1KpVB94fPvhsL+WIGtzzfh1uCjuosfciETQL8XqCXhlevxbDGuKssp47DccySV0
lypxQ1x6XjQx/eUvbGd3ECSEBYZPwFv2C0cOkp8SB3cnmicmlQo7QmIfJOKTfwH9sdc2AFeb0VMv
UfwO291Abdw7dyvc2Gd1UKAaBMLhIuK1W+lVZZccNzZc72no5xUz/I63NE8ZxOjrXwdhfAT01Swv
YBwLUxZZKlG7QwAylbjUWCYIsDMole0raiBU18aXVTOlqjF2bpZe8cb/1IL6TauMHxz/pWNoRMYW
hIXWXn88gFEkhUG9G9vvV/p5gxSl3ruOKFIjqI7fjgGPWICVyRvH0GOR8PJtu3CJkBgNNg7TiZlq
Z7+D8YzdAAXiBU2/JT60/KQbZ/bxcC4ePxaFMGn153lEJXCyqPfd4rEN6nSVNt+0KbIPHreKJAem
+J61w8zDYMAPfO2OEHqdcfoht2TXndWQw7iLqIwNMzWYugYE21j+VyTOJEPiselcRqVhw5RqzFo1
RSNCVTUVFuh6GguzfdLaT/Gdg5IYhZrtO/o4RKWSod/26fSIr666L+KKnK7iIH6aGNx7dqG8bSTN
rBhnDIEayMn3pr0OKd2xEn9p1slF5jBQo9UvJtHT2lEiJ+rmR3OcDPQ3q1Y0K0cRd8Hf0Ns4kdCX
nn7KDCthy3NhLffAT37+o9pc1Wz2zaG0Oz01zQKNmdVaYn/fm+tJzC5Ngxv25P84Jex2BzRAB+XI
2o3QSF6Mg8UtZhK9Nrj3JeIvGHTQZum5JlVUZzFHf+OjFEL5LAR3CFpM9SN1sVtISUx54oRwvhUw
lbPX/cdP2YvUv2IgZiVwfBczMpFXJUSau9X7WszAI0o2XbdgAtuHMo4W14tf8AgJuuDCUetc5MkE
fMNb8LiNKdi7qk205KqPX1BWQ3komjmsdJS6K5BD2yGvoyZ5814GbIAPTjoGGEaDSR5pzXF8Uac4
45lKK8TljvYq4kC1/qJFtpSsqLBnBifjys+ugRlPRgT3wHbOnozJzI9VQf0xTHdonvedXEk4mt1A
gsdJworbK9ugvIXLZhhYlVSz7az0vgddU8daCGcWUA5xFfm/lKUPCeMjtbgnoXSSCnEj4i/BK101
toPwEZa/jLrcTZChVcbqHo63oL4g2Oyp3sCojIH6WDX+wJx2DAuAqI8JHuNl4Sr+iJMTXz2ENZgw
zHTglgylfiCObwJmeYENrIoly3LLFIs9oFHGa+RpepikF5RyBkYzAeonZNH2eR/NEgx1YajefZcp
JBhyT81JnaUVx9zuiAui7UuNEauULFFhu5tG8zJU7wajcimZ7aDsMgIjF8PCxbRap6q0Yak4qcW4
zx8WxOHWFGg7ccr+WPyBnhjZxGeePLX2CrCB8dcEd06pIhfzRpWES7CP/6Ir2JXQggl6uQ1X2HhN
uoliGOzQeVOOINSb/PIzvsGeIsXDNsZhgtlE4Pxz4cBCQ+/6X00xf1njju++B+Rg+GoiDPLOKdP/
xBYzUIuH4E42eD9jsFllwxrPVQwatCgFrJzIk7eXbnWasBBqBrXzGvXqjvGddfrtw1qEgXHEz/2O
FQCYE2UvlXugDXfwje00Z5nSRmscq8+w0r7NoZ0zKwXP+HVaQZARYqeRfnuHyUjMi6rXQlXG5+aD
STFPb49vt+GPkjyshNPX6QJ/Qar3fNtf6kyKOEM98Kr1SlkTc61h+76prweGXUmIi3kVhjprNlCK
i79riq86xKjpa4gOKJzebx+AVfFFI4SZCbp4hxdfTE1mhKzueFRnlLxGD9Fg7JvC+LQLWEuwqlVz
uV25OwrrrIoqipS4rmGXLm8OE5NVTNeuuD3kYF7jgYtLAk4jwA3BZI0T8F6nAAfXtew1NmpUisqL
RVmWXP9hBw3RN5uR8Muk+9C5ADRROCuJmp6hg/oKhgLe/28P5pwF/p2BSo3TnkDKDWI0iQO2z9Ou
Dc09/Gv2UvxQw6nrOL6u2LbUPPv6PD77fV7IYNk2gACbvQBxYmP3ZXLa+P/Zlk8l5FWe7E/6fff5
6W/kwffMNK2xZWrlT61/pEhk76cjx3e3qPWlK7A/g0S2eO538THIHY8scPlv0rkYNlUA9DikIAK9
4f3lkX0FlsGGTXBkemzZyXJJoo9qaNiTyejjF/ujGk6CuYK3iSHSV0Z5PcdFm0jphXlIcl0S1sqb
Q5Z8WyfUk9Xm1d6O0INagVqQLCzKhkEYlwwCY4Fr9pq1sljd3Dbp/lDnodKnKSXryJ/DT3vVbclw
CE54/5gOT5T1BHvib+M42UmErLPSUUvEDMHpkctJMgHCUact1wXB+zxjh6OOIIapVjArnOM7SMp/
Fq2QsgOfROnKAVgKgaLNtoYSwU7KxDXrrAiSewI9zuuAWOCPr2UPK4ZDzjuorqkP/cs3xujAWnf8
gGLzGdHaeFjo9LLzSWAy/Qujh67yRx67exizetfqfQifzHTyM4sdUjELV9gS1oFyKX+o7NWm2Bap
+ipkFwQDpOIwTAPgSsxuZltz3jb0sLbNZ6lA+7XROU2EW8TXn4leD9D3DlB8h39esz0LeHfGdK9u
KqCRPtI8Olqxtb8TUcBAFIvVQnNwgO7Hr5BzcX3IORWVMIdvS/m4H3o8jtOgenJIueus1DuRyuoH
0e1MysS2bFQy+Jl7j2/qbZfHDepsaZxS7wPVAt6njDme6PYoQLr5bs3YxYodCuQvmfVbkLv7T7qE
kuhtma9SaT2uXIjbE5FP54SH8SnNGlRPUa3SapCATbtkoemkSjke1EmGZpmna4Ar7p8ZXsKUzVDn
oy2O+FD4TOLKr8lPHMS4NqxjjhPs9a/k18/WEq7qqEGwZtjvbnVtnVzDg25NARQx4TrFnAlwN0sf
iroa2yfmRwwBY3zd/UqX6edwErGlecF1mVIoy2aB9JFC1NKnawyiY317BoN8KVT2LGCKFckdnk3C
aBIgdzyfVbmqhBbtalQsbuNtPf3bmfYj9ZxnCs0fR55RcAG0gNHtqh7WlK/nNSexqFRTY1tw6o6B
wyCn5Zp25b4kiXpRFtxFWUpK/mVL7ZznOonUc82g52G/FXONM/BT2xq9/qC93oUVraM0O032k+uH
kf621hKH/MtgQaPHXYKLToFmcHUj/fiFGUKumYoe4VK+nGRenReWnT8ZGzxflB2pVJzNEGitfP81
/3IVGGALqVnWSNLR+5dgGzGD3hFFv7RQdqU4XSzUnM1h295VIIk1AmJIMcacNEHdimHEaeDidvgC
Ubzv/ULYqmAzHXEtHQNMIk5opsn4r21kxdAib+iXyOqvJW1Gjmki7KwD7nod4VFGDmzvr2kZgHy1
9PYVlfQcKpT02+aOxYWBiHT356O11nAmbtpatLw6vPMeAtUbyIEHZsBIc/1BQZ0ZP+vuXPYniD1X
xiKCnM4cIDqrb8yqzZkC7cR15qKur6OzdtMVXFRiOURif70nSOAR+MXNZ+C4mFO6dmst7DJNmHS5
SZ9r3rYc/T6Hmelo6ND/TZCVPocMeNfZAA3MpgMVDoZH/LhOIW6pPNpaiwELNu9BtD+nrqgCNEZC
hgf+SHAE2aKZQLxR+6W2WotpSuuiDptGgaQFIfkhmLaMceSQE418BtqRLSdynJmtizHZ3TeOOtEH
YLX0jzpI+OTSERUIyC79dQYBCNVXCw6vhhBT6UKknNHgHOHRip1AHs6UIamI3WatmcDY9ylpfkIe
nsQdTHZpsExrjXzQM9UoG+nWhMRgH7DvANHZE4iEeis4UwjXZndxl6aNrvKt5KJzVhEz4UOP3uww
76ixrjos7GK/XH4lc8HjCFLk1SzHDgL+17q8ZFqKAznHQ1B0nsLb1+autaGMbnG6rtebwztLMOch
22PwvDne+f3cjDxP30jgNxv8eANjEq65C7BSIXc6CqJdm5M047UbdkPbxV+szpo9747yapxt0FNe
9X4j712YXvD6YoyhZ66RSpF1+yFgA/AGSXsDR+EwOUwIFeppy4zh5X5Ltu2a/3gOBluXO1MplDyG
c3lENGKILQNaYuiyeZzgLgt7xwGibcmPuf6SQIbOtTI1WUhR/eTLrMrukVl+eA3bUT0sXvH9YHGc
h/c4QIpgwyVcR/s8OxpmUahMU22vuv1U4XgoAdCicAZ7lDNec7KN6Y1G/pzCMlzdpmEfarryEXqp
xXemrCO0q7Xt5GKKvZGvdQdBNW74HzdSMYTNx9nAm9YwLzyrikLJyErz1098HxRIQF/92H9l0VD8
/r6IT02IjB4YgpkMkY+QWCNs2+v4E836LK9vCZ6YtbJEH0S3yIabpwo6bt89djq7P5f9Z3guffo4
fFhnl/6EJk2VX+Tb67DTfgpeBAmyWaHL2nhMYSCQGv+z3wblbfrqEXObBcnJhbVgOzoHoGPOcSVy
uuth/9xQ3pM20KYcchevZ3ReaneOIY8hnJ1SPq4GBvp3uBDUggXg9J3Tzzqum4v6wW1vNsmgcCum
5xy7HBJNXxtV4hD3rT+KKklUuHCSfp9dVLauC29Mbw01FWYbChnuRlw8pdOoF2pcxRIRhaiSedxJ
9qIPaWKklDDQGHADgS05UZbIsJfcrLAy4BADIyblhQDXpULPYMo6aZuUQDhTquVrvzMnD1G2Ypl2
J9utkz0eMnWiT8a6TFmnrkgoT35W6qkTRepC5XePg2PrVCjws8fYn1vc7HgaPvo7oPcllpPjL1en
+4f0DrcQ7iez1VXJeu5wCYG999P9aPhN3WF/1hxxHSeSX2CknOU+ATBbj2AWJFBVdy0vO2oQv0XQ
dlaNMVM3I5QUWt0bsfeSGehs/0sH4k8A4iRbpNnIhzBjD1NK77V353SUWLpDs9FGQpA29olsIH8d
EBk/5t6d2Cd+TMSJOfrLVbMF7IGXK0fceMNYJVsYxb5L5oMp3ckNaQDJEHmpUb3T4zsOCyESLEKs
FO+1MKiuhZyQk5Yr1IavS0AwrL884+hjqXH1vZqnLQMHB3Ktcc9EFY5TXDz5ZLVw2m+j8LoNrzab
hTM6gq3M3vouWxwulhqfumLZaM7UNW91dsRCRHzvqrurCWrKOt1WkfpIAQ69ldxaTcNOwCZYVSw8
TwJ8V8TtsXTeBcSJkuWr8FCHcSpFd8uxBC7OV86qfb1MOBk8O1RAhCYAtDC4jKY8mNp9LBJiIaha
W9nmq7XQqfghJERUcSF2s2SGAjr+bSaV+R1/87/ia5/ModlV7/7EpMpI4pYkl4dHsb+Qyj78q0US
/rYlxEiAlrjpwTQt69pynqG0WeZrF5MPrRhgKKO4nbuX9eaxmB3+4wfoV0WiSzW27lC2oEhZa4n6
HqDqz6YFLFlskU9FARC+P1Gb1d9oEf2f5i7pd2Pexc2BjD0giqsD9B/lrX014XMDd0mLxd5NEvJF
V7PF1QDvVbOCMLqw/RqM8WzsZAaMwTQGS0v7QbF4dAGHaXjNxsQ74ShvDuYDiGFhR/s4Gc9Evi45
v3c8rlwl7q/hO/dzyhluX6MCW1lttdXEuGIlcHuAPI9Uv06H2aTfdvdG/aZWgAMvaf8dCDKsFYba
hAcjGSb+J2vFwqRM8gNMygty0kiZCIa0x1qrAxFYzN4Fond6t5PoK+75IB4Ot26Ht9V8eO43UKbr
djKvOsmT1kAZqybHvdmfZkyKPaBTUt1zIBxJJpA6S8CTVE2r/1Ws08PJTjXtBQZZImzst2iTS4ON
Gjq4TWLJpS8Z8QVSo0p81BbIb5YSo68f/t+tC0Q1ueCIhxT9fptR255CWL5w/xcDamXtH2X3jTWb
UW3FOLpg0NgF5Weq9sW0cT/GkQxTU/y59yy+E1MzO3nRNrLZJZfYdiD+nn0pJKEItq8wRSdl/Dau
lsX0a2/SPkXZ7XktOCLxA4ae3GFigcrJA0kSIMEuk4QFkcLMGQqgr52pk79bGMc+n4ELfQoTzk1t
NLfSr8P9rvjuLaiTvwIJqzfiXchBHEja57Fmb5+xj16zIfGuR0pIAZIOfrKP67gRG9jlSGhYUX7h
wy+JudAWrmzJotg5pTPi8NcmHzEwusRXYNRbq3VAMlmdmzYVGXUFuiosoI6S+KcS51FSK4OGK/Cs
kYvWSXLuFILdjWvPo9Q1KRUv8yDSKA2XgHriXrtImfNh5fRspHvcOvzdridq09kqbY/4lZdSnO3V
EnWSGlkSNKggddu+vIuq94AKzYaaD5f7QKoAe1lE2zdHkw7mWWGGhRz9dyAYUzYkb3yzsIrRcEJO
j1egZMwSf1OFfk+Hwq3GPgBOryeDRPQX+oo3N+9X4hCvPKQk4zR8b5yEZllTm0QijttNy0N/VLpp
qCxdDGljHdfNRoUN7MFvkuoZNcCZS7uyWj7kb+mf2Gh0TjWdMkSDbHZ2n+8WhhWboQoKpsIiJ4gW
oLmXIi0PYwZo0rCuYtBr8J3sdgL03j9JUJVVOrOEq1hwmtddcazVENwssKIBMIZtapnxbKX+oZJv
SGFN8QMEuiIV1L0GUEVagoWrB3E6jhoM7n2ykkNTHJVemXp59oWKEnG1zOKhYtfVmOv2VAmLIuYt
UfZPailZHZUp9Rb9fz4ecXwy8gM1aSpHon0/P/IAagIu3ETZEzLn03/Ark4RlZ1AXQvWjlp+ZXpr
/vnI5hGleurWNGVUuOL5jjejhlzU5PBC1nYIovszJAbssIDfazOhGQ9YRpPrNbNlDmLpBSSqHqDJ
7yb3SQf3Kcfotsrb8Kwsupfyj0XkZBvGhJxuMcEgOfuIK8yDDTCrnlIA4qnVBR7Yyt46V+lJClB7
hcmYCJfbKtCeGLzut0fy3fz1kuoGUNJORnmL0isp7RAtPEeL/ozt4voYdjAKN6mTsQ0n8/wmG06k
jt7EX2TP7TILXhZlOV8rZMNLAbqgRjpUWqf6MHXXyCtBccqmMfDPHcFI7oTbGzjXoPySNEMWjmft
Wxi8u9glxSE4rhoc3lEQaHCxE2rMBLIoXRIc8PSITTB7HmpVGLfG2EZgjC5uxLA2LxngD1o0QiCa
b4aEriFlBHg6A/7G6nLP8z0aBEsg/wLZVm4kpycZF+fsAMPy/w90DAhtaYgHG2Rfl5D4ugiHnYOJ
nsI7JITgU9v1X5ZZ8oZTSEJcjRO4DVfGZuZYALeYtVI0DtF0mni8GP9WPjAhOuPi0yXtUB0KZI34
wvm3vZ1gtxMl8uryj8VbdDAZjCqweNxuPWs3CqmixTqLOQy4rGwkwLbnDvnoYpAefDvpVPQ991Ij
/qwl+7BUOkqEz4L1r8EJ/1yrF+XjT6hKe0CSWqdYDgPXHW6NSgpHmcqRQESu8wisBtPc23/ve4Rg
+iUV2NJ63yrTy53qD4iCluHTalbPhH7Xr8QaKlEmNaIJdcCUOcZGkIJ3+2p26p9i8927B0nGDXGp
TAOsrrVYWhRRNn27v7b7qah+Y5C8jR+SnqLYSNJt9Ew7CiBJNR9RLYj4jBUDDmYezpXDQeQkw9Hp
4edyw5qAfxOp/qpMmLD8y+ugXMU1nAa/2CsiZ4jlwQgfzvkVWVDEeIa6JiHoPfq3geXHiNCfTC6p
H16psR2mjcQSfSFEpi+c6o4RFP6Cz0clt+jp0/KPI5BIAWpZdLucntzY4R6+8blYdUp7GRLD3HTh
bTnZOcEWJgNBCXnTLsgEDL8iYHctetC4DceT++yzG3/qZ7Sw6wXOXEM4RbtsMqHf7ug21khpqF5P
gywqdAs7MhT6ifTq69FTcNhvpsx0tTg8+2zcyerqGmvpp/KZXtAKb60aQgZ/RA3Qq/h7sNronxXp
P2Gm+7ISeAp2nZKbxtTeNSGCwIeC4e4UcpEgW6PVm3kQm5ytCFIqFdscO3kuZmlL/1cA/yOpid+m
KV4u18QTyyZZak7i/mfb4byglOD6KhCumvU4xwE2gTSAKFMgp7tz83W9lqrMYqcawDTdzqsfyvRi
ZSZl2Y33DnlCgrDdsvxzqp9tZ1lCcYK45YUYgPwQ9emdXJ4pGc3/l4M/fxgDRyJaB20vfYqa/tBV
RClB0ptHAV5DrPIA6CLceVdYpiclxfR0VIzATrVVaibdOJhKWj8KxaAWLaclnfmxFq46LaMciH9X
spZWn0/eAWjttFw3+WI70El0N6BUU7EtUuoZER7SjazpJ7aSd8+YDtipukWRWRLiAWpJWhG08ROi
QHUN4qvNOX1VtviFDfFJ87RuVdomb/n33GX1SxjquUyuSX326hMY3ejxX8pfsKZ0yRt6d2buyWiy
vqyqGo5KqwGMiRMnK/YDIZkhTDzP1oxBgxrv+vzhbDPs7azvHJiizZ2Lq7QDVVPia2/SrVAUUFVX
i6tMkScwNJI2nNFUG1parW5bJBS5J8MEprH8vQuSdENYZkRLnB7Z9kO0PTLL8f6IkE5jugAGDsyG
P01/VTDLMBdXp9FfZZW0k/m2YSCoRLnlP9Km+Ya1zU68TqvVFurxL62At3Gmf8rkfbsGT9LcdKWV
ZDzAjA7GIuNdT2Cns10zSDY87NfSxueOk+o6II+pne59xlMSe7QQDAcL/0vcvRrwGnQZyKJB0BS1
QfaQm2R9aOCUDu7KDldQRWalOWz2MO6sODMxGj9NRn+AIk3LulqtFsxvWZSYDpSigi+dFrvMK7/4
bXSDDReqli/G4/DqGCiw5bHJysopjjBIY1fPQ7rkeAAEkHz2Ilu58v6kRUWaq6uN+26uTLXzopwP
CLc44CV9HWgmZSObr6gMmGskyux0J4rRijPuenEpOnplQ/Lgcu6KstJcxQRi75NXAHGoP7RasxN9
tmwkRfY8OKjpcPhErj6oiFZIYEF7l4xSj3aQZTPfyplPkYNMn00EZW3o0l8sLRb/AMrKF5iGLhzs
aPVGyV6hfeKHlmoE3cCU2klAgdflcfldut70cHjpAcfa486I9Ddd9rYK6sDmvqAqh9Za6lfEEm11
LhsI9n2b/R7WvFzxwxsnl08A48kyK8Ebu1LBU6aZJVcuMhndgjDHYnLoCAFKXhOIGbQf3lkRKpGP
PKQ++zlD1+bG2FE9zRCwwlazqVtrKmy9nvcwJsG+AFRuRKWCfjMCJ6tq+46OI6KWq9tVxpdcTvwB
w4UPrjWHOoGMw/EUuPd1AoJtj8S9nvEWkaglVIYOmyV/97EIiVbZ9ZVY0vg/Kd63PI0xYVryl4WW
ep52/YRmOvz4U37Bpq61yzWsWZ9oda4s3Xk3NDE1xYjLh2rlxzMvZfGQ03xdjSccyeDUgtmTFi8a
u4mPvNk9npSnGQVHI0YlZqOAwfk61uY+rB99IMGNqG9jwoS4z5becfwNzMQ0eggnz/LG+l1xDS6Z
kWhxSx4xns5nV3o+7issJfgq5q2kl8KlgEXwHLbAxOUc3brS89oOjRmIq3OAeM7M0ey9EaghS+z8
3Or82LuK6AbuEUGUgqbLlQQAUtB/ei3ZU9ZtOGJG27lkp3K9DqJUV26V5xH0ichqJV3xpnPk0uUp
c/dOjB+EVdtjKxjxmJO4dW4iCHVcspKgEJPsI+ZIyGRJPpJENdO230GPShZzZYVKQwEyhP48bNfo
QJkvFIXgSLaNitHyVfpnSqP+lklm1jHxdbFj7Pdpz8JiyKQ0YdSjaUoV6O5p4czdbG+4JNaMREBx
jrk2nmuG+4r9ybwLxP+IoMv8tOPm9hkdZI/lRCBlsthlEMYxZAKkLGvDTtzd4TqlLqf8kWIbDSni
cci0jtnNNhIJIhGeJD1pJN7o64qR4ygtfLx0njAYuWDTtOS36RR5yQIc49YdBmmXwTeUUHNM1DEy
ZWoKHsKzdGINy7/D4kWsSd/Ff4XZxxaFWgGIFyslleKk9KukVrkgbuYpEVyjtTIuezvn/nRhO9xr
cPdUwCZ5GGA+ylEoGiDggnamxvtubbDaFy4uRSG+f34AQL/kkReejfnVcJCtBHeUJwXigqT4OO3S
5UdVFm2NIyp3ArJdqY9KNfEka/qzivFqXEhMvpbmrvahfaG9sleLvfub1y70tF4kkjKtfOQB51bi
7dlxt4xQaoNo1+XLoNHfQ+y/ynwgSbTctarkoqCvqXow6bBG4z6tiorxFfLSBoXsvMjHMQuXNsBz
C7kaoUSdr8k0zhoERF6flam+eVYnJTKYs4lLsqccdUvgLhEugS5fmOFg+djFyP1OhEBCiyqhOr7n
bhxotH1gvtyihKg625r+U+TSSGBRzIvG7kqvdPFOawFIRVd6MGyg0ATO8/yhyezwz8lvD4ZIe+Vn
RlLWLehoYS9SYvW+cOFJCcAZULX99Lowr0lUpLr1vXkXQ/t4e/+h2zWYVbc1iq8ArIN6C8YX6hxR
vmUtUVHC5AHRv6CrhyGVdPFFJkVsO0LIKaSj2M23V5XD62kBk5umqLZ46davr4/bQyvq3Z/4XB85
iyYM5JRV9JGFwJhU9yrkwBgZkIfCKdjHFoiZ7CeT8mZc/HpJaoAn89AI4A/HPjCCbVlhztnw1pDD
kG2PW6e0exzBn/oGr6wN7xJM8yqJS7tIgKmOXRGUGT5o5qFSHe2QSsaSMdHhFk/nES6laUYfpEPN
K5eCuBZoLXx4QAU7aEp3G457Ll+xOQyvc6Iu/T7ZjBsBDSkOmw4wuf7DjY0W/OoOb1tNqJklMIE1
za6J2eex6FZlCkAmQEnW7U4KbtRPF1AGvsRRMs6EJCdAvHAlzQU7kDKY6HjeQOmP3C00ffwU1Dxo
UnORc1xK6wm+Tlmg3a4iZma3EWT/i9JKmHAQvel0x+6ac41nuV+R9yPXCrbIUxhwexlJvT2aQpZs
R/LlaHedTUkIdllaDjkKyTYH/INOZ9L5+4f/FgWTPvp5JHwqVcVoTB+R7V7I76XFeZSvHcHDH7cO
ldjfrRFSsfUCK8W9yId4kjML3X7vaT+e+vBTe0PLHrLbA25FqDZfP0Vakm/v0aH3G+2T9UDrlc58
f8F1dvYRako5Qqc1XRnUyXyEaQnxXMI77g3CwXIp5rdhMkwSH2IMwNQZzaRWT37+nMt2DW5etT1b
b6eU36h1tyjMfLc4nm06iv3ydnZTNJTRyg17qXyDTn5X7mu8XILlwQdrsO4+/O0HytxFRI06CNGa
fBqgvlyLABs1VRASDMTvqD6bzXK6Ti6Gdpmu+oI6qxKpK1rHT9sTClhUhIs8jmJTXpUPv2uny5yi
Tx3/RpGB96dK92MF/5/mnVDSGHdXgyF9THV7Orz6NekLDW7TB/KOc3m0Sb1IwefOQhhuufBSiZ2z
HZU5mYKAqtNzdjFJAXkVnely4DA42Ur53NY+13EkTlls3Spgbc+nYtZ0WpMnq2ys8DdBqrooDm1e
ry2wWj+R5C5ZnSX2L7R1Nw1b8B7yhhqOTdXnnnvry1fMsS5MByhss4HilC/zfRZvlbuOwtMIGrQ1
jZLQoJH5444A5h3BDQt4sUbuCoqPQbkaNhIiC7a71W5hIUxa733G9b4pvfd29hGahHyiSnhurLV0
rHNNc2XdGLU+OTXRzXv786SDDrj4I65eg0ccKgqNKbXWdoEIQemCwsvQycxfpZXmMM087x2Iv+Zt
ShAgWHQEz55dVdFDMETR3k15FgTlfNQj7ZjQUs7fDkYOb26fkQE51GBQgFCZqzPWMIT2sN3VuWbq
wunbG4ImFxohMgo3FVBJ1EuQlqwLr5yXfNymS99xVBXM+frOCloTQZoxqBHXEd7QVv1KZVLNgfV8
PWU07O98jdQuxSrS2lOPTkKPn18XwA3bbZo+YlbzzdMFaP1+ZnVvAC24/Op+i6lRFd2zPLLwfwIU
3HIbxqP7kS4NQ/jsEeVjh7f/oDtGxfpeEkyCL+FNemzcIYnpTH1F1/zzZ9SwX38P9DG7e67wZI31
NVS1UIz7wC06swNVcEsw4mag+TNfquYdUsWLFx9ioBn14r0vN2CSsB1bB1cLKXSx/gnXwf84Iktc
lHr6oayDB4ziKEDql1tYc6L241l2zEx9khvtlO76kPtZtyoivWF3MUYiFw3G8Hp7/d2UAumzRXuK
5Cmk4YV4RBo6/mBAyYZgyhJ56yXPYoRFY20rGdqLQ8L6iy5/phoiiRbViQmx1GJRHXJnikcXYv3L
ddoicQ92ccniYNNqlLqmyU29n4o0A6NUNZORrC01fEeafYBrRkNPyb8PK4fGIfCmKZM/Op2P9IrQ
nBqaULBe3X3b120Yqkfd72khbTuILpMo2F+IC0AZDhR/UhffK4MeC4YfZVoR4bYGKR0NkdFEHJmk
46Xgs+HO8ZEUxtigzURA5U8UoEIjpUg6qH/6/5vmllSpBkpRRSTIuNRZGH9wfOX6I7O/+eX3wKE8
xv9nqcTFm0t35poEKye2eP+wwx9xosEyFZaoBbfMtsOAOnzPMNGpT/2cHGprN7Xy07lCTliRVT2Y
wxBnRHzmkzg/KbavGScTdSYnBCa9X28Xfy7P53PXeKP7Y7MsyAlnNMNtdNf6O50yAAjCdqNHVQpw
vbcVaWbXSwoCfvk5arfeAleulEuZrO0CghVpx/E4eVSyB2r7ko0avspetr3Xi+AXQp6Q1xeQzcWP
iOhALF7X6dH7dCLe5Oo0o+CKusHNYt/G0GLpuH7+7QCSBoLZxm3URldmr5klyr5LF7gUwspgT+kU
pnafA1z/WGWZrlK/4EmXTaKXWXg+pv6+sIEcVLpKDWKL+mCgpbTlr/ew3VqzcbY1Dhdu/ljXUipw
hqGMzPYnasjKp5tC1MDrJW2HdaM6PM/mLKQVXtwEhDtnpFfJUBJlSFAJ7uZXbo2kxmkkjt+BZ3wu
l1qXI1nb5D34tR4QS6cOS7EuPpIc71jy78KPT1XhqNKiADEITEcTQKXyxC/uQdfqLYeeiHrHflMs
erLQ3m9zh/vMHqfRdnWMngAeAEIbDwvBfv9YDKn9qfjScbTCvtZ1YFyZL+OlIYpSZJ+kN4raOwkW
cvI+v+H8rjHblp2DG5/O2HVF1eSbzA194iEXT5teFbeIY8etn9kG0wJJv/QxjnF0U8a+fegM35wM
jZDAfOVN0mc0GyPqG3kLl6ULtP1ddjV1hoAeDqPIbfWXhWzzRsdaMLR5BTk8ymmTElL/e8aW9gtL
5yWnIsFiQZG5LVAVH6vb1ee4gGnCjuBKH0Cs2jijwm86WEfr3LpxVed/vypOT3egmGR4r8j/9t0O
rKIzQxdreexc4Q/xJ7vhJ/XsEYRp8fbgJLos+xiG/6FrGD63gVaxfucq9zAOQy+cLrGPTf7GQSvk
cVx0l0aGM2hlnzfBG93WiB7oMZZJyeLndtrGjLh8v87CjfTVC/BE4KJesBPZHzuN7066J4jdhC6Z
9OXVoiWDnMCtSaaNPC0xJiWfov1u27kCURnrL2LPW58+P0Vzp8vNSapD1VZ5CUvZ4niFnjvcsxYm
AVTDM/Z/wcPoLnIgycw9bTM5qsb8ior+4IeJ8BFZaMuTuvRn7RJ0iH3z2pHaMTyrOKbyKBj/AVsG
RSiAS5GPWDv0PHFLjIxsmz2wvbNQEMJJ1IXKfckU1chqktUAatca4ZIi6fsmnDdZsBMKWxrQYM3G
3VL9A/hp4ek8log8+5tAqxShLB8WkAAeKUHjbFNZPGIisuBuOnw54rOmXGIPq3uEoRopwWKodni0
KX5Sb/Lcj//JiROEt0Du8ByCcU9YLMMW2JivvexiRMDpUOTONKrKNJ5Q07UXY8b/rKc8GR89vjOY
DThyoLHtnpgnDBP2zegKrvPtBKQh3X6UMhIi3Cwx96N2vtieCKPV+k13mULFaVN2EbGbVv3Btswx
Qk8sVCCgSpGr7SrT0CXCANzPDB5Pef0zYPh8WivHr00/FIarGxLA6iid6O63DKWQ5aArfvpqJ3Of
osydp/srABSw/OKURdIREDC11CacGW7qjth9PK319NZAgkttMJbMh4CHlh0MbaP1U7H2Q6KcDaC2
8qumfBjfIOJy6kcNy11JshDXEcJMtI4JQtR45Aj8WDK4zOro/6t/Ex9gvIbAyp2a/uImw+gQv9aj
2A8HP+UiaB/FO1fo7tSGkrqclQTV4rSNLhr7gjJnTQ0/3+WK4HhB8EVI+K7iNO3I9fbOj0PxmBnb
KKeNolTmg2ro0sX4jWAXtgLcHHWsxoqDm98TVcC++tGq7JD3SWR0VnomuyTpM7sp6YiDrzcuhAb4
Wu8OmGybdDKHCZfYo3a6aUJe8fRXyp9ygIvFgzmSm5IzIaBHR10jimF5Yb32I4GKWKAF7NzKfPbU
DEKxND5hv2M12jLZMgTD9K5uOb/+8/bWYU/oKsokjVIAq7Qx+FVF3L93NsDDqLtrEqwQ40o+E6iS
miwuJvQYLJpeloPUbgIqEBqWj9DW4DZ66gGs9Tm1kbOcjnJ4OFcUFsmFwXD0hnDvi+/JpnsTu7Co
BJPr+zWlh0OvpSs5Ew0LrhgW9IlEyfZidX8WKX5YpriNCz50RssEasKvfA/U/utXcjjA+t8joqaF
DWu3eN+YhIHlZM4apHanjCUkjFPxwq5J4Cp+FH8BgRx3wxq494Fg/3csiGwjSwLx+BOejlq5k2bT
2dLwMme6VTkMoBtZqZHW5q3yCuFRhgPEGWtCE2ZTZLYVmPk4Q7sTKjuLO6t//I8PY8vmG/M0Nsho
WlHpxCuOe6bZlE/7fxBXMGqBPTEOtQ9JLiycmn9i3E18f/2oSj+INdMbcg+/a6N1J9LPhbxwCKn/
uyEM108sZ/+gLOzPdD6rwJAVB3P3jE1UjwvnZPFWexXUJ/y+DcVckzXPMF6j/H0aQmUfXo1d57XL
9znYFah29Km+/eJAvkSvIMj5AqAC4qokqCCUyrk24Y4uKsUGk6Gqt95OKkcnUE6LDMFUYGyezbhK
DDl6Kj/INs18Ef5dlKHOBp60FPmUA1Ns2qjY0ba9NTAV8ukej/69/uDbcu7BXr9arLXdArBQh3i6
7USQjzNVFjV+K7tZ+0M93pV3FLTIAnjlQYNFtsoCxJ5HNgy7d/oh0lDOPZDax+uHFJg05NWp5KPn
5VphzrBIU63k8pxM9XMsHQzQDt+Ni57QoRKTxj8yXPD+ufc74NHcF9y2yi63qiOrIa1lcGJaghrk
tdMZyDlEWIDiq49wbzosUSmZpgwR+7kBHJu6yGU8rStbJV0jN+aTGhYAIIUnImYLu7kw1AdsuCot
YTJ6xwEyNFwuCeFo6PYbKQBMq7oJ42Ge1k3yv/OxI+LrmO5x0B7dtoK2wn3Y9pgRRqilWnKgRcXC
U2+t16tXwjEr6LjM3r9EfP9TliFVzHwwHY/9ZqceihCBb0I+kmdO+fT9fDQJ970vCBO7A+hSekyB
IsO1H6GkS7ybT0de4kniNyJByxBrG0Da/J8ShVde3TcUituKmHaZ/Vh8AAgxwHCDiqbLoKH4Dqmt
z8uQm2jYUDDueHawVjvX4eQgxEy0kf0TiAWP7Um87CXhDOcG7S01gTTKE5juYZR18b5cbeJiXPTH
J8cNaYgfYSBJaCKG685IyTAScA3fW4rj03RzCo/tlzD50hZcJ+Ni1MsUjkl/iXVPuxdKMhTfJ/Y5
lbbh4ILqZ79bFt9zchn6C2GI1ozT4WU133/DUo/v91yyZq1rKR0SMeKK+5O6G8ZPn9i7Rzlf4c9E
A/YVfcCUGHVM/lizvVHP5+dcFjEd4X/orIQphhoN/qZ7QGpohc8HXytCy/KBs8tX2bHjic7e9TaM
aUO0fWHVFkZ1kXg2AjxNzrWyT8h7JbPg3tCisNgFdP+bfJuOAvn/zxSpUcOybU9F3ydQMzLYs4kw
+Z4lSIbHpGDjSq4d1j2ZF4WXblgtWNUE56Y2ETJzh1oHeadDxKGjssRgvtkdkOoys1aBYnlCZe96
4f/7CiIPZDL+WOCU546nU0F/fHXexzPzSZ+t9u4FXR8utYE0OT9P82+mZxiCUBALnoF22ME90d/V
bnQP7izEw89CHRB19+GPEN0MWOuWWdYHND/AF2BCVkjhtrN/pC57gVEIcM0S7yi0FUEQo8bMwxYt
C0ieGl8f12rPDgej7W8jnploHSd2zAw7ogup1lXjT4lB69TipGcf3bochaJKL2iFFG0YeO80P+sW
D15DzG3OAF/szgKzIwlVE2RYU37yRkfEjWc7btXWquYY+IdqjZZowIuKnTmGtE1yQnFas4DdsckO
eqo4pRCXNFY5P0K1mMYxZ0XTLQpZ3csmqrQmoIU/f1NJSbx6ietWSFR8ty3uVz2VvjxGMz36Zn2R
OQtT+ElI4LNPwC31wVw4bkkfQqxooL4UN/wjlcSq+mM8daGq0K9SM8r0OoYHPHcRHX7azJ4f1Oxq
XFr9/Jdk3hzlKEFDe4JkCn5jnLSYhLTooLyD+zbdU35a+6IL+pEkF1WH1iD3/ABhUPxKTt+v4ZTf
mhb0srVhh0NaSBZacgyAoLCLaGTV5vIPgZqBEtCdYem4toxscT0jDten9Scug/lzX1u1dpY13xVf
Vc1ESZRAlSfBryysXx9d9co2Cx++KwSUVcFpmWDkV++8mOkiEOz3iVo9VkK8sTKMZZ3YrHqk/XZY
uh8ZVQOhOMLxOVDnr8MuVFWUJDkiaQ+r/KspGcW4J3DlL2qjTLmx58zfu+ikKfML6UxgksiSa96t
NLfHuh/LiNW7Lg+0amdSfiDdnfWpCmGIubZ8dSgASekzO/K003NQdUT/JfONMResINI3fsZOtNVG
B+X/QSfx4+oiywDd6Eyuv0tQCS233BiWxq8fYGh8eW/yb2Zgu3lf0T3+01+SngbJxiP7sjmIFVLj
YBM/jy/p9mEXzbbatackJAKziDcVjWWu3V2NZSK99VRIc8jLyUNa569qiqL6l+D6z9yEc4TGKaYP
oIb0Sgnw2Cc2tk553WkJZupqOlNw32Yqw6PT/5lwZ9YkmnsIzNN/ZifF5wcefIM49ZJUX+Wkw//2
0tTBoX79Vi4aa3caKMG8U8yyarDnOfhkAGQTZIPzZYtgVuWDCGRJlIdYZqBhMoGDyDazw7x5xyvd
+JAfgfIhEpT3x8qFMW6A1c+JwSANwdaYiqPw0dfgc3M3uHvbcGhacdqioMsaqOjDmfnFlfIF3YzA
wgS+Q6G8iOfFV2xTWqSu5fuqwI9KU7BQzBDNIudXL+ihVSjV1NXy2ammJD6zfsOlCtKBHL1PGCFj
+LSrKpc/cLeJ1su5OFBC0A5/zcX+OTbZqUObDI/7iiJFclGHJeLI/UtHaPcbwkfweEo4seOkdem0
VSN4C7pP/yCTFoe3BMYQWltu/xefolncjNKowBtcS8Z3lr4BceSes185QLJzhYocrq5tpg/B5ZHS
WJHoHR/xBDGE/2mQ+Sk55Pj/jOwMWNINKER26rLbHf7BrmGLqrCQppNDBuo+A6AUkJQod4yvyy3k
/KmDq4OaaPbdYUp2EkjxRHOmLC8H4xPEeFa7h0Hi0QyPXtS/ee6KoM+0aTsdh74SKBv/rWyDQAfu
802eBxbymVmXN44gPOODMiJUrRhFPkWKEGNlkp+1yCuehJXy4iBW5Ce48jrUSPj53HU8e8mvvXDk
WULPDWYOIVkhWrdcLCvr7TEoQtf9C7k3njd5UYWhBvyjINFVTYL06sYBY9RAi1IlJ7xHdheeOf7C
aDoP0O2Vpe3ZkJwl2AyJYKScu5B7tF5iVsMCzIJyc84qmWGOjN7ELW4f9V92JxBUXRWNAI0+yK2z
K+uBwwA1naVw3pbhYU+xvrDVj/s9zLCkDLmqxiyEykUeYV2TV0Z4EnSh9mk6uVvRCKSmBEUccv4W
9b9ZILpwNdtxDgzzY+0FjrkEXEQNJCWtruMTbCJ8ciUB00zekO4uZSZqzAsMHrPUyga2guZ1XOP5
PBaNmjBtdOZlVDI+nGZSYbvKDDXO0UCslXuir1AtisDYh5Nz+Rx16+PtRrmBQLInw3EQfMx/iBou
z9ZclGhOUZG3uYhrI+/76XEbVSv6j/IHZSKAJVxOASJlrlGhh7L2QOSVYNNjrze/Ax6jM51+r9vG
heaF9pD3JzUosd7ciYPu17NqJZckNOVYAhmIAV/PS7e+pj+Sc8H0rn0sz4NXfDPljQbwiK52CH3I
eyy5U2bTrKYpWbzpCtvf5SduwFDqiZPoIHL0MnMeaNr9S4U44NAjFJJnDiOwQlZy6CHDTrH7OPlG
H1i07YJLLkgtKW8bRi3e8c5Hno3RK3NwCXqapsByOzB5cXAtUeyvdWWr32hKyYt+bIL3LMccLVjn
9RZYYPXQMHO6PIUMTb/RKqmLtEP4sFVTYLGj6ib2JG9K/rIPpYgRQ17zwOgDiMHGMpw3QSO54Szw
s2wvMAWk3/frq85pSubt7XOIj0Jo+DQLE66Qs+Y2mvCOCcnKhF30JqzIPiMkQvqRwr7RfvRS4Ny2
Dl6vPBVmtiuIllNYlheQoYYz1KKwg2i/vrjRtS0OdvHNtM3zku136lDDoP2VAlOGt9yS5wZA062s
oznjMObfm7Kcdk8h60ufrQnpFgWaSjpNY9V1YkyFrnwmb2tz3/QRCxC7dvGYuVxfKQLzM/t4IO9j
64rOVlkAI7HcIWiCyGn87R5dlnJIuumlv0WdsCQyBho0k0T65hH+ZIS3ALOdkAzG/B05gu7OUy/z
m6V2rFEs6kCDKyeOxqS8CTxZ4piQI02KX+x0u75pOPRPWoMLJH/XLrPUpgETVXeiWzB026x1mO7k
1Y3VAFHEvoNcwjiCsbSJexjIjBa3BzBcf3Lw4eqHlTqszMdXyvDgVMVTc5sahBOEoHKyT9a6tGl4
XveL9NNWIZu5Oqp/kBv2TquQqDFTTmzO+zn3JPFCQr4/76qMVcP+cjPPPYWO5RT0fGKDU2/JylwG
peUej0cEqi52tgAWizUUPt4ScCblsx73i6LaqY2w5SLCaf4/dvR606E0IVqJqS7Qi83tXfelAjKz
J3eURakXFAcl4ztuH07ugtrHTYj/MXBEHzrnDH2yNNYYgh9zqafg7GM7EoM5MmqmrYLBeNFnwTfx
tbaa775TKpJMahYGSfjVkED1HtPaGFHeQ2eksI5yyNC7N/MK9i59mHVvKM2l3Z77IZI2nK5cczFJ
FPK84r52dNbXJtnw2l4IT4QcOTDTy2EV+cq4N+O1JK7AULana4N/Lh3WsqHyVyGs1L+u+7b+Yyyx
Ay5T8lD9CT8T0MQZqR6JLTRQFjG8TJCkKCz4S1luWzGxakkacbErYA1xCEkf7j+axmbGhNbLpk8W
889xHrLV3PPNb3v4CeglkgzSlYdxfDesfeozBtMJNmxlbv/zKF+Yrl2pownb3WesC/sGKvViagEE
5ZrrAnj8iG5hFe+yUJpp4Gn824HYg1TaVcYvcwYpey8EFevl1QbvCnZLaVVTm1ma7Zmo2bnZqP74
axOfP7T8dld4eCdD9fHEapSP3SfE7k/sFwGlyuNNRGrgSaCanfAesFP3DfVlcDKSO1kskeiD0EvF
MMyqLUz7MEiMSYQuvpDtMUvRrC9LPQinV80gY4foaBYpdA+12z/ASFSgvTRqgDLuAY6ODJLVHpF4
oV2zfDmOdAFCMF1taEpH1izTvYfvEtRTNacoxbFQ0a5R6s2/r3Sr7l+6K4N6XAZmBrtVZIbfjH23
faXJ67blKCu4lNMl/azvvAUwT0XQoSuTPnqixjXVmQkNnKTKov/4rwILQYjfXKl+jtW86EgFW2Ix
NpjCf/m8RcLUD9SI0kZUEt2NlGHOpo7i+dNje36kr2KeMOS3ZlueFS6b2yzzTEio8t8BKoOfPPgC
+PxYlZKPbfk5/byPA1Po1dCbkmXb45bcrFPxctEnaRyKLhR5SMuB5chSaA8gDWFHoZuP0f+rch+T
QznCQ3nNbKxPKf9dhiIAjzqJ8DWCXTtO/qCsoUx4pLpRV1cRVigejqaV7tACRABogUNMusmcN7vQ
WDP2XixI+U+vYyPJDjwRt2ERCnHFbFQ83D6G6dRKykze5wYx+/oDaw1hOwd1/ddi71vRdN8YoLFD
PKhGWPpQ0POBYyaQVKDxBE6nxHf5kZI1I95Ed3KzO1D7GTvsgeZV8i/XSK93iy7/ZkWlkqSvwhuu
LpJJxXEfxwYczRzd0b/85kwH//C7uiCEA7RBaHiD/KxZ/ZM1AHdYXegQhjOBJNwRz7J+bidqRXR/
oo0DRoUacD0fnVIcwh79s+4ij1XzYlPgJTqbnba/CZzmA25F2pO6dx1SKnG6WWjolrEtvJzCRchN
9RVAtTiQ0i7WvoQwFelJVyKyXkJS3QEOUDAGO19HjTAaYDo5pRtVj2IsDQ7VJ6x+wNlxS5AfxXAP
JXPKYc5s0gAMvr0OnPfcdMTLckMfXt9RmzkALwQYsoBMRvfJNfpoPFsifOctXSTwc9ftqrSTW+vd
IslZcpPh0B3iNIAMa0r8IpDWv6rd0BlkwPYcOuR2wt5fUIFr2WKaxJTLTlQqlds+bSDL55xZVNst
/iErzV4PbY3VhnOTfHtHujktHPbB8QDRND49JaeA/YUkT6CdkCVYnGvl8rHWONypsgZKxVeXae6F
gKnu58OVRqyf80R3HwZQGSHB91utyENpgUf/l+/elCFJ+6ApmycywvTKXY/nY/yxrvkcnvwZx9rs
z+H3KgkVtwXpFWgW+QQXvFzCBZnwFvE2qUlT4Yra8HssedKx0hychtNJ229i6JVxIeCxpf/my67G
5+Q78czlWIBvq+og9zhQwtok5mniRmi3tkrH7oduGrPWq28gBTljnq6rQg5cgWw0lgLwi/FFCk/q
uiSieJAST7gy1bYY6Q7uCQWb+MArU2xGFGlRCJqanfKe12DUD396ty68xDxtNCpJkTq2hZlxAVJQ
mX6yxQnRyF06ksSXmiURvwUhg/w+XMpInxE/leM+stqnDrGVwvY7mQtDXmhXp15P0G6jBMeJtlN/
8smSAndhnoW+HKBV6Eba3jmsXbik5gpDHeSRXLq/Xb0BrJ+at463ciItvlOmPWuQTy4LnsPWudRU
iDUyPnRbw5jHwinWvJ5o1XWP3/auyLRQjOP8YbfKjpc0rGC/A4fZwTJzZO/aLWzlwBRYvhiqnH3x
+FkLlFepdjD/zCGKDNjmt/JarxPwQ3QL1GkCoJFWelTB57WZgXwY8TzB1mS2R6FqVNCkaJ/fFDtK
VFWPgfOX1/z/+7aea9Ta8+me72hZcbNy1XZyO9SeiT3lL8kpEMRez/yJ2yzgvVe6DDeFh1idCg8M
lr79XIQkaEganIjsgim9E8HKdsoUPtLkIZY1KLnhKR97vtX0xiqgM4oDJXDngbGEwexmNGLo1dBQ
EOJd9RcKZEDn4pgoK8+iYDeXVkmOc5/t8YCuMieT9ccAewZc5EKCbZAwnduwJbr2xB63JaSRJ+0S
zILvX5yn5gfNlB8Fnxtz5IbcS03HOfOeEMqqPdGfz8lsX2FC60JBW+Jgk5e0a4DYNDeZQsfFiFiK
chlWz5lp5AGp9TC+60vi4lKd3eX+yoZSmMozKvviqB6AKxGxlXs2VFZllWAzjok+bC9iP4E5mU4D
dOpqgeho+MD3D673bxFjf9sh6LZWJRPh1EqVZBagzO+TsF/FcXWmuu/K88SpXh0IGSCGXdh/Qny2
LWpebveUxPQKpAFtEusbK8HjUjR9o5/RscImZv2Xs/QTijnLCiI0L7RVBSbiPB7UuvWc+7584pSe
r6zpsYFrUCMlXplhDv79T/2XnQ1MuhZWrX9Tt8MeCG7QDr6NSUfT33i4NZinbX0dnPh7VzohNJtj
dpW5LHssh3f5H3+zRMMNxfbRNWdUNCfNA6x0QokRQlFoFg7hRRfdnZ3skvRWFpXPa46AASid31Qs
OWCNExFIW0PiPr9S3eKZm+l8VajwBBm64moKEXN+KfZx3dSJKoFtWbWqd/6DNTL1LjEVPCrb+42k
pR2YfZmWtI62yLQzXTXe0SeBODjXlo9cN71xkaGi6PMp4+wnbGlwVWH/+aRsAXLKtd5M2ujNHZg7
5wa8yEIAXryeWKtEMguWhPQMNDkkfEqAP8wuWazIXp3AIO/uPGXXzfGIHl+VhhAiMMpXnOqDFuWP
7zxZbU0VCDDQDlzoS8RygkZIugsaUbmGJd2fVm8C1lMQCPpM6F4vzwy3/pfy1dzHvClIK+EGQeOg
1SbMMp8GFBVL75dLg1oTcU63xJMIob4DNZH9paHaolsrkjGNOLLY/r8+ow9QC+/xoXie1r4UUCxE
8qUgPUX8PBE4WnKJcFn9yC/Bshdm50MHd6YHM4iRVcwJ8f4nECyNgYb/4tIY6FbFczeZ/nV6JkZJ
P2Zu3BedMCJ3GFjG9b7FBYDjgEAMAXXTQuK4U8iingekgH1zWKIl3s3bwKInO6LYOOvepJMkcyzq
GB+1Ebe2AnAMLRSwHr96/A2G3QBzq77i8m66AcJWiJ/c3ISxUSpoikFQnP6SFmHxTpNUMTP9GGIe
zTZVW/G8KLHXtJiTKHX6A9+9+tJEWAwrCprTfhIcWcXl0VKDlqZPMOYR27fdyf1ORqnPxCq01jG0
CwojfgUUTryZA/EI2sJZCDvUFC/BqlXA8ilP7yqlyUm4km+zQoMZGi9YmSPIo2uQ+GJw0+xdgLRi
k6i92gGH4Z98wzI/mMv0Bm+mXifdIAMzZIJ8uJV6sekTKBkPmW0cI94IhA11qNmxajKr44ChmrvI
nVXMFMuP6D65khqsaGTVmH9M8PsJBsVh7FkbbEgn+8rdcdbinydZHlJG/T5Q1gwQZvQA9XIl26tX
XJZ10oswFI1ReRrlrDlQKPM6y+eWW0sYzIApmxzQ4MLy1CXg4SW7kEdkqsiF2PCWGls+0tqGfIyW
MGuiFYTYwJo0BHNB2ng73MR33fcepPbpdJN5T4mcQEuSYbzvo8WQylnc4U5BRMyYSJB8zY42KjVF
7XkMxZ2kGuzSe2FV5pdd4Z5T5HkF9nv4Rbx4K7M41upJXkfVNRDWPHZ+cDv9fBo+Q6FBdut6DP0J
AmJURcdBA7EJWg235KCgCNXLz4BSQ1qTZCjn97RZC/Y7CemrdsnRbFwo2ZjtB1dVl2wKgDc7Y2CU
vtphd8XhFQthfaczExjxSzIJQx7l4eTFt9PewJ6r3tqPp+63tHgKxgtM5ax8HTo/9URNQ+XNjWFR
q5V3Prn0eqVuFhlaMHdR+ZkOJxowOMHVG7iYEW4v2w6maeojtLr5Q2tEagXv+R/WeY6hNfbLYGFg
XSrapZHCykXQ8sWKWs0rmUHEA9+uwI56cz6w0QX3/4plOdSDTfQPAEMeHJJnc+1uEKlSgtdc1o6C
byN7TEOcCwxWSyg2WFXhNbG0VsVrZbTkr2+ogCC8BN3EFCvlw2rahm1xHBrQg4qW4cm0xSmD65PV
q64UQZFuvU6lBdCIoijGMAUjZtvnx1eXx0D7wxfYD4OsAgA394G+NW80KVZGNM8vAjhyFq6NoY0Z
sVRnS08QwFoXJciR3bsb4clIqIcku86QbZAfUM+XlKvYxwY40HnMxBUi/1Ok1Ee27JzBhVMkiJzK
baCHkgnS2u6LavaAKawk0ExfuUt1rM7TS27CPxmhCfF1VVV/aEoy1RNr/aHgozveCCYl7IanKFew
rYfWKlVwRbbFWgD3nSJvr1ziDz8tZNYk+by3qAYUIBy1hMxmP+9gmmEJUbaRfBR1jTYN+iH9QgVH
v5od2vGX8RTuPQUMqntTGJSprn0j7YUkwPD9oHutRbhUmmU1VBJjkPp6XvmW2IbItPKNlYZ9Gf1m
jfJGdOi+8KaZziFSbRbXPnKAA21Xxng2HFfec6t+Q7g78g/dM4yrq2QfPnmMxsXKdDzX6ciXmASZ
X/T1qaJ7d2zodaw4rSOl8SGOgVEB6oFBcoB1yzZ3kBO5kDexa6fNmjG74IFoRF00E5AKF7Z5fpEz
K83TysxG9jk1H7o7EEa/PG+nIMznWLd7aaob5sC2A2ZoOzTFWs4uvkzNq96uomVqeHRAApUhflUd
77KgEuZV/GT9i5euO/ny3sVrQmYd3UU/t9Z8j1lRZWsxvtc8ej8ctYhlGSbUcC5dAlPMdEcti+Mf
AuhGDebmk7GagCtWfiUxv/pMna2IW2LALP5M/qDVK2ddmWbcQ11J4APoqly/C44+VHhXX0OOTAcl
RR9V6UJMx3OEoSo46/5yYHSiHV4SqlAWzwckpI8mBtjeEEZArAw2+r1bjpf/caHx9cIo/ivyAKJU
RNtJJ1jPgaIac26j9vcosEdpbzczT9E0Kwskd7Ah22Pq8K5XGw+XRtj3C4BF4F6Zwll/AweZ/Kv7
crtAad38YU6ue5n2IXBgfBN3vvXG7Bud0QeQNvbRP8O48rj+JI7Ssg5QPglm2N8Dg5GuS9Ntxs56
L3p1axhiL0Mf/6mx8YSAbnf2CsrU7D1XTkpYDMZQDKbNBj/bi8d6I7wwTSg8zAQDvWxyoNu/xzsY
g8ZzLPTy0SzSYfXrDr7fiTCLmmU7OhG+jxZQclaQr8HfSrOXuznPpdEhbK6RlnQ+xWdsykS/WY7W
+5foeEIIzxMsOIWnjcyiJ0IazXtSxM296QNq9KF+dPn8KP/qKFCkA2JwA1RKjaQRh8OKCJaqyDlp
IiNn+7QzUStaPmwiasFm5Xf+YWYkSj1iP3KZgSSVH6xJY0VmuAb7kEOpZnSzYFRECnCLaxSOuyXT
RT4S4yepIxQO8sVLEEIsPqH1wPSOnIVdAL4/pmxois0gVbClCviKeW8J6HKdhwLgSIK7WSy5PIFL
dZAk43dfTrWaOMuQNSUja2Pg6uTzKQn0UBnfQErcQGxsGrjqs7lB3y6PhB2Nh9TU8hfO03x/Ki9k
GtNtFqC5czcBJ8BoQItnO8EPyJX8wGLK9JnwZ5Oipxn3oJzXsR0VdC6ugg1U6x2hmW3Dj3TP5tg9
5wbyMFbba1AoOy5y8m8/RaxRDv8CjX3Uvvww8aRXBz53zKHYwBxmNB3wJ5hmZ4F6CxmaR0ty6vyJ
EO0I93k+9Z78b6a96Pqz7I7taeuS/RLa1wgGd4ZvPf9Jpes6UkUoKUj0WPYvNrxJ6FQ9S6btFlQI
pNVOie25OZgTTNZevlt/zCsfjK4sWUtpSzS8MhNFna9okaj3m/is1AdF7wylNQ/Lze8PLypE3P/W
mTZ5qbKPEWKnM1rv52am6SS88/ufeI8B0OuwFEf0kE0h1e58KM8xSLRRUk50a1xEHaX8S7Ygei9n
Y6683JeTzbrE2BdGV8r9mJYt3sNzIzW/YJjJcnrPw9OEn+aR27t4j+p5TWC3+hwYlX4H5GMaG46L
wQoHp8ymEWtC66tbEsaha1xlPNRwLwX1WJIlaMHhyygP2RHYzYOOPhGCN28FJ+k6nP16PeO+xPwH
ChOa636w9IUEcPfnNsVMojX3CGu7CFRyUVTDFuMJ1PDSbQOg6LjSBN6rG1ARwtEBXAISa+JSFkte
2e2nf8tkKl2m0HA2rYmBSJK0v8xmdygitImoilxgX4cmRriNik9tn8UI/af85V3h1UDS8VReIsOT
doNWFVhIKjsjCYnQxojsNlkODJ8T37FOG9ls4DrXFoUu277NsgqsGxl+xdhApzt6aF8K7S8Wk0Ls
3ysbGeudRs1iDvLEjmWlNpMwKbxH8F0/p/9V66ivjHnyhpyXHZpaveIfo8XneWfiNV13LFFd2llP
APBgLJEiehd2T2xHkqLiqc1uSW60YLTC9n+iFjAzAbkkZjAPT67g05Xox/yV8iHKzAQKUZrVHQ+u
usOOzt/Mmnyqqd/fgSTQKNruYG64T1myomsfbrXzlF/RftyH6vNjhdXYSSIK75golvRp05ybBc4T
gsJaAVZ7ehQKcv5igcbZRiFvo2U8DWwWhJ9HeiW0qbWnK94P6V6yVG0LHnxuhaZfbALcE1i1RJjI
289uW9Cwy2+GGlFSNPxtfG+RX+TU6+t9W1bBmkDQPjeJH18+b2LPWxsLie8bdyscG4IMzL3IJPRJ
oj02eAKzRLnwf8YQ13nlj5czSMkTbmSjTAnsX8ffR0i79A1BJ3SDNJ4asTszL8WKBbES3Pk9DU52
ojN6cflvDXquukQy4OvwOXDBYsV8doBsx2FHPWKQzWFBTry/S69idLLVgPpMPPotCexV/ixNR5Zk
bQtuCOaLVNXfFyeX8Blh+js2eJMKlvyz4tpHgkco/hfGlzxZYOzJ9YSJSTZb7rPcFlGLvWqvKqvL
kZF9nzS129jRhsrm0opkbDY9GDB/CWN+SBSrR9rC7+JPly66eCPl4gX3pS8GnEeNXe/yHxqRazzn
r9Gs0R3YmdDAhUl0uf+mCMSn8Wof4SE8qP7WwYr/AAL9eG9MaSaAaDCkrMFR1bwrthUuuAF7jtvZ
M+Sw7vFZMdin2YaWBlyyCdGBx/s7RFxp3MPhSKrSxcNRWQ8e+Pou5xQbGEGWjKapWYTU+Kwc+jnp
dC31LFpLRIP09UhohG9+tAO4f1n+dBfwawuquPGSlAOwgM/3iMv10ZQO3fVXUKCm56s4t333wsxH
JwPR3V/AVbEkRjAQXMnoJncMSJhb9ITKA+lyS1cuXqTvw8ujAGtmjnlaXcG4yE5YkgnGLTUtUpFz
gmDN9S9J9ESfHPac40G8RTlPa2uCpOQn9LRH0h0BbtG1BLHU+ti2D8zdXSDw4O3CuhbOxO0NcBTn
ybaSOBJRz7c/fF7MML+4J50Ts0azR03iNp/VuKs75+UEbEcJcsmXveWL8/zXJtr+rJUF1BkQz0ut
nJWevWRTsw/xBs2UW/3Bx3TKef3Rt1Z6gl9enBF+xDAhvZEGEyqGog5Ow8uUn9fNbaWdYwfqHhw/
5mUKhNTSLOFjwz+ezyeVVosDMvz7GuJjeWBcwBc0Czbn7GRKikYfS6qLGKU33DJtU99VO3/l4kat
iQPpsrfapsW95PUqEqqW74hRwwBqZd8AUCJHrhvPJIPzaidUThUjO9XFmvKg/D7bagcLTj209riR
54m+cyeYovcmW2bk94Ys4+4zJaod24AN44ISjfXJhif0FeveC14nqAnUQ0YYNOkLpnNLj1Hd78sg
bQuEkafigtKOBSCSBUBe/tDG64Xusn7dw5miNa2/Nf+KukEVORqcuJNYRPywAOnIlu7LIIw9F7XX
GHnf/4mCkcRh5yAmEp/u6/920vyfTJJv1q9QrVQB9MFgG/58oGADooMii2obWkMi2d+jh7pMUTt1
55DZReUCNyL2b2obzW4dWRSyAsamh6B6TTaZfic6GJF3CnyOxDehF3q3yND/nnr/FKErCI5o8XyD
ppyk1Tm9eg8w8tmzCKXkJP7igWjRxnVDAM/N0I0OZGMY/GY3eUzqB8N2eEuEunuPh+J44ztbqnBY
a/pXPAC8+rlnvkCd8desRFM9Vl5Ezna4Wwbx9TaZUlNW790Dy5pvDqXN5w4KGT/YbuctMQW93HWf
i3so1TohPxDyzFvvql9izWGbSsaoYj56X54TEmFT+HmveuY6SB4xL3OC1/nVIk+divA97q1ofqr0
+OsyyWbVU9jbFQ54D5mKabIpuwAHcocRLG1cZAwXpne9LoVQODkdQXKbIDDcG/iiz8Qy4St7BDcz
HcoEyq41T49kVqudvdCPRb7piKa4D/kqcyV1XLghf5FUf3NRvVwVcCk3tjYsVOPV31OeVmR2ydld
+68SV5COWzcaJCfZAALNLe3cVP3IqqlXCkQexACOpj82udWm17GGBG6xemWtq1WyCPP0tWcWwW9Y
GIWd5s9dyVkJMSv8tFJ1WrvpAaJah6H7Ym6o8c2lO0/B8n//rgHo338JmNvBirD9DutQJqJvK0Hd
zvwExskEPFAB/0b9WiMuBCggmnKIpXNfAL3G72r0RLwSW1rnQ8vXZ04ciGNdjF1hDo5V+cmwADEU
tV5t2HQyG6pP4uHKK+/VLwivHYPKgPk9aXXZjOITJHY9NbYyeg2HJ/4HbezbcvZMTQsA26590Beo
OKC2eA0sbOD7AKNnz2wVeLm0kajCDqUFYMtQ8sskwm3li6HsMZLZQm4AyhdRCxCMNHLp7ankkXfl
br6SxRGdIylN7OSnmZfyiIbp1jI/XdfUqpKVzGkB9dzqRabY2EJl7NgvdHp8NLOZMHtDbzDMpHx3
BQAMaIQkq0STTK0mo/8f7UCp2YaW3LIiicJdq0xspQSeUa66jUBmrmUzSlPLzlKvcHVsdnu/kwCA
ZoGum3hJuS0+R6uHePvHf4eXsJRRf6EZdQt78Xzjge2VPr7xcJRayrfYZbPMhxhMuT715fbCiP5Q
QmjBLgTqFh6DZqEec8RqwZgZXyhBG4WTcYoyYk8vV+/wJ0o6aaHuYdbiZaXCqQIIYzZuTNaghOF7
fHNITMo8bOAzHHbw6kA/rJpRP+Cg9kYjqpxMEwQE5rXzE1J/ZBa30AKY8A2vdRtTLkAHcLUcn/er
w2rRPla2BZ/rozJusUWyezajKjfTr0d7Z175jZgZ9m3mJlAMI1ZMevmbj93CDijZFDt7yrEDYCBL
s78eBBnk804aTShyrN2mCj/LTutckOdTM3pGJDMRHsOMNSE/YUNI0ZrCeI+kyntACnMua3iH7JJ/
L/itSEul3jjTmJYGnzG4ddzCfpwf4q223EtsYAT98NS+k6oTFjJIdsNxmFpNtgaekBam/n6F7Atb
nC8ofx013rUd/U+cjPe2Fc9klN0Vit0EZZujwKBKbqlRrJY+VRezz+N3fnyZNaof6XPz4XVxQj/O
euI0Je8zaURL+21BSG71NXB9fETHtGzDbNz2d/QXhuJ4b3FbSFKtK4Kz3e7nFOsWKdoHGze3Zu1U
Qvzk7rSIf/wpHWof2QIwecE3LgtBjrs5bomdD0S/9ZKPzt4W0dJGHSEyljP6Xkn1iVlpSqMDrj29
cwS/E8XatyUXjDCKp0JBPTBkcw8gzErT/mXBEuYp9KykBqo974DPGnN11W279NROgDEGzcm2AxIZ
unz4SWBBUvssFZKLorQ4RI0RYn4+x0u2dPmW1mJ0a+UD7V9uktaRTblHdLZiYq8cCvnwgkbMfjaW
1Z698NofUPE9SLfbjQ1cYEQd7N2G7+JhCtZI0gw8VrPg/jyh7DmJx4HWQIqceTEWjyg+hB4UX6Dq
3KtPv+bkXEElrD6X9r3qMfdMAQNBEMJpgQlvAf3TMtaU1r89KiGoNfohLBN97u8PjZpS8BTHMkkO
e/yxFoHYUnzexkMgiAYfArWpn4m/lIoRoE331mVw70DzzqNOz0VhJ9RhbLZdRZvehR9MG38TMPvG
z2R3Ym2VfWxtQ6Deg5iQ2TF1mi9csffCxuTqfXMGVUWPcpothVsPZ8kdyKns3PtGONIZNq+r4v8A
h37RTi5r+hCwG6SVcQaJ+Vok/NNvsVt2hshIKD23p7aUOn0WEjs+CK0TPoa6DOhJuJIT6a6KX9yy
AmGjDytXaNlmBFR8kUFJMWy9nEjWFDHc/q1rNUjT7RqLKIors97Psj/QbNqcJHzDit2/o4nMXIAb
YFwICm+mun1Z3qEbVQ9PlG7Y8RgrFcPD+hGOeJaFtaGXAgNn89AdyEsV5NyM/AWj4+9ijAmtHEFB
r8iLSrjE4vaqR2BXvbxltmvYyK4CRAKHgjvUAVrN2j/3EQIcHTmYxMnLjDqF3TyLOmnnlSjFieS3
k+0z2dLJ+969JUautgrbrUV3Sf/ZziTMxuoWRChnm6bpNlD7t5moCmONywdS1HUjgDpGrYOdrbVh
NjR1H/zA2y4NKquNaP3uO+6mVX6j8tLe2KEVBG1c6prgSmXFuXNCjAJWtE26UelqB2M53BSbEM8p
Hez2XI3vpu0Ppg3zkoJZAUkd3HIkEhMUmikkTSjEFywx/MDGy4310frIQH6QVn7BYF1z2Gumgh9F
wdfiRL/CZLGzmsywe9P9MuA5XqFbla7SrW0DSggk89NuGbuGA6AExcRpHCdnlaihffhjohv02fOl
SmF+upMT6aVkBaKwpXh1QV7DazMN4u9V8adhuthOm4BBh4TBgPyeawFdkeqX8+sMv03Z8pqfmK7M
F+AMTbD4N7jmI6YEDOSIhrusF5+y5X3akxXP2aBc5AypVLTqf8wuwoBTxGqWcEZEJOCegkfj/TFJ
BjufBgdzTH40/6vjpA2kvfQb+UKxR0IDjpILpRf6OrBtbaVA52l6JBn0R4tdlIkOsroP8zqvy72U
x5DjkS/bsnDz4DRu1Qu6tvlqrQVYJYBIWDg6aDH22ez23HR3zQqwTAlbg0MSv4kiidNqv0o4e8Nw
stZw8TBwmaLiNYEyZAPFkm6ucr5A3PjNBMuOto/7NNQAUSVHZETfyI4rfj9/A1pPrRd6zQAw4YYL
OJ7f5hUzAXDBQ19MHUS7HnAoV85WNAaoDxyHVa2ptlwrGFlWfZ0hVMU8vJHUC+RsazOPGJDOTdC/
BTgn6HTFWx5+pUPgvzYrudSSa1tm71a03pOaYrwlDI/yGI2Z9nxemeLaK2JUtp4auSmPhoDk6HGh
WFx9VSKL6Nj6bHcjybSE3ucjZJZIujxeec3idDJUiTPvBRCk3YDwhf9EDn8eKw/XgVVCxhVWrDV4
tqJC0wb78l2BximDlHlLm+cLepqXGozgpY+cZdQgcoKDF9SltBNL7pr5o15ejWiiaW2Vgra3CMzY
63p+OmcnPXoZhPtTBtE8X/euPmPXVaRWlTaiOpYtl7DvTIUIm+Fmn3vL8p6ga6itQx0VQdpUIP7P
BDmrVdnSA1UAUu/Q3bzeU7wkkbfw8jXRM2dhIosu+fhpW4P7ZofO4hg9jq47Hz0pS6ttzUEvhJJH
XHsuKuSh77xskuTYAHqjol+u2IGr2IC4GJFiEZ6N9NYbLm0jQoi0ncLh4We2fN00YqbWYLFN09D7
TAXHSbIt8M+2L6xMHhRoQpLw4viQ7RIw4x1tHoBIcKwbixxu0m4zm5YNO6hBR8k2eo3BYOb2bzrt
MoXVgpJI4I5MHt5vjiU3J3fD1jOw4xvCxnG4YEhXSWRFm3oOyloCsJFGGtJ40HHe5hcjvcyhBw6Q
xo3wgQMoEADXGnzdpHrKQLkPDoJE4YZBA9qDdZxw38BwDvLP0zcy9/hwl52/jW6z7jnBze25DJTy
8e6KhaurgsxvfYrnB86UjyfsbiTEdxdDJZV8rnxp9LHiOO1d8IZ3+bu7BqVfwPlqUKoMZm566XUI
0JivMACgyxbukkzb8Il6z3dTjOnXiV1PF38OFlfx26bXocBsTX2rxYXWWYeSXm5RP7PemJmyk43c
g116jGwbBmmGsW0eg4qHRCvZq9BCu2FDPvO/gWRReobeuT9dSG4TxAc8U/I8o0FyzcWPzIgkrwjm
vDtwigqWP0oLytzu5LmmByfso7C1Cru59ecKJK5CXtE3ZhQp+EqJckvQboz/1sz5Bwue60hShmEP
iDecFoFXk+gZ8HWwOCVrsb+GH7EGEZU19Jh44d+etbWiB44af2G9gTR7E2w1SuEeNvqv7oz1l7B0
6zFR11R7yKvPUHCB7EJXKLGYyNfhva61/jEMaABOt473ZMWA/MundwvLwpS8v1TdIFkgU4wd2DDW
DMMQM+mq9hOx5Rcp2vuQiUAgD2fMZ6Eo/Zc9H1wSXlKwTH/UR/hCUbY2r4qUm1USWquXxPcyt8K1
i7hqoLYX77to2UPBhuLHhF2yNxX0jXN7dFM48b4I8hObQ4NUSiFSNvid0FGtKVOf/Y4rc0HpbijN
JWOg7/8cxQonNsMwa/JwSedkQcQzdtklfeK5D84CXxRT9nzZsDe0Il94sgfnDE/w2bUBchkUksuw
bIKG//LRbaWjPLaPucXYAmnqvxNnjUu2XZpAYybMBFI1ts+sEe/uvX+Obf5cc53KXF+8/s/fQRYQ
zd/woGwPUT4af1oZdtlLJ5Y+n7yEa950LSkZU28PiRTPZPNIjNo0i7xXu64H7ubPfNEltPtpKBPY
+r0rjVrIq0ohFwRrv8n26Zz1k3zPUrrDE17NVBErajpyWPpFXMf4zJRiLRAbqE4RqhiNHiEfXPdi
Y+lKSdvCI0QFXXpgQw/zR0QqMWP6whd8TKzCMqA7P8+EwPXar1zVGhB9xQ+kiLr8olwHdO6te6MJ
4zO8fj0OQde1BnH6D7HtldA0lcYy8sksMbaO768sbxInKUAq5DH3LIsqaDRXvGYdp22WXC091ANI
CfwDqnLm4y3dilBniw7I9QlGRuSLkXxpr/WpMjUzAwS0O5QLBBPDoPXqJiJh+DRYzY+PQvQt/Ago
3WwlqLJqIfz5zW6gzchvpK4U1b7D6r/PnSmhnlLQTbwLav4bI7Po/dpsSaFF/Zw4grb/CGVvrlXt
qtNuvO8pB1FbGO1uyZ1Xn7A/VVtaly8UkBP+S07GugRgGcSwPgwFSxo+vvdUIbmGTyVamSlEycEG
3At4m0TqEHD68MBTZY/R5LpWigaT6RV0pec80rW0Iyx9vFJnfQ9vXzJQfwJ0lyvK9EsMGULissN1
iDNB+ByyOHL3QFbCtaWV4EZewfrlK9DrF9xgYt5qt+LpnCmrRgyHF4cxFswx5H4i9YCEMV+gycGT
EUx8WzF/IvdyRLPc3ohcYPEoe4el23ZU/3+46Hf7KcBjI1YRPd9thjSIRCFOjeeC8CFf76ZD80Q9
8z48u9KwcRYjo3/M46AAjCxOOHL/PgRl1SWJcROI99IhzN+cU9NZrd8RRi9cHKrBGJ0CWVkdBy87
DdOr5yCLLmCjZ5c0njJSVCN+3+fMzqpusDG393mwIoLXNx3fefqmBI2mBNbFXnZUsxb5rba4VoSk
CCL4k7NxERzkgIiGwe0Z6nNeo2fXo4amaURt+2wRltLHPlmHSkhwyboNzC6ubQwRSg6LYJBziB+R
rqMCrDMMRFDvq7GFcqmopFeyn4a6Pv/NuQ4tH85YeItiB0zTRGibLJZiiNbKFwyzh17CckyRRNX4
pS66lHfMGLwCc5USVZU/6XYirwRrIrK34KVUse3FrX6e6ZoWwNueQirKGIr5aVTOLXP5+yf/45zM
49x6pEA2p+OzqsnlAJCRmmt3Sjx9D93i+dmtt6IUtzKOpMIRdkdot1m7PyGtrGgElr1Lhk2lD3lI
yWw/9vpGXrYvSg6qIupv+YHRrmqIgX1aTRzG5nfr6tlH/GXCVEGRsCKULTDMQewhWbUndt4ME3jU
5oVmxrOBIM7kd+UG+1he5eSUqDy0tZv97r0/hTnFqgW7XcfwkYSMcgTJNjeGsoxYepi3LHGY52M3
w/F+DWYqEoGHra3GDb+fwfAH7SDUxZ+M7J0NRt4LBQHhmk4d/wTN+G6rnlEnLO06V5rU6vfQhsqX
cynLXsl0K2v9Nd91IOrXB2QeNcKR/MxhBRcf4DHNTdixQBOem0PGct52mYE2+zyv409Px3FCzKZ2
2IisAqQUiJ6K61tc3X+aIpFEluBUfzpSWY5pqPeZy93nqz8uGjPfaLdOm05na0C65sfbCjHfc/rr
GbFBzbRaNu0YTfTAvyu7I/+e23gAi/hIeosOqtH3IqMTGSnHndbCcR5j5Fma2SeThBkhU5gWyAKI
QFfx6fOkZ1WVqRaDlvFP9b7Gnfq6A2kpUsYpRAghJPL+1XxDADvU9QLvUeGE8919Xh0khXbbScPD
dFC5mgVSeBSMFhk5qzcHwiEdM6AcC9hWmpRZIzOithropArjEeW695G058g3v9AsTKqzY1R+MYpd
33iLq0wXNWSL/Zs3ThLoc/TYICgyuB3vUcLe9KfvluFMcYNukdTVtfzMiPgpSURZA0TUYRS8neGR
D9jRN8vPKMoci0cRGZHyVk5qk5K25Fi2ADzs5q8pBd3wHyU5bfyR0LKM1mdljuEJKuc9ve+odcxN
lBNkjNfBaUBh7HmW+cqhQHbN9pZQKIovPWw+35sw5sXLBPXe8dQZBpuErGV0wk3ATAf+dsPbsytd
k6lK7G56dlhDZv/o4YuUz3yFGpIzIRp60SbKDgvNzQLdVMZF3Kfe3DhLqOdG3Aw8vdHenQ8jlLqL
9b8WHFmPKekSmWskJ5Qs/UYqwSbIvAEyyo/ISDHrxtYErW+XWJdYNDQSO3d2XmLkH62XoZ2huQoK
w5Lge8op4AYptpckq04oyewyiV8zba++8q8Aoyx31XqTiWpmfjtktQ2Xfq65ESHuHtprx2Q1r7B9
sAQX85UzTvwPvZE4VYx71l7ZFEqiMAcEt6ShHr0N2NNNaQgJKCAfifPk+BAeHhsHU6r1EA1yK46r
dmGsnRImiyhCCuwvL9bAYo7XVRD4K2OS3gt/PpH3qCRMvSJMXBki8G9ZuM8CZe7IIa8fYDu2XfjQ
OUbXr+ndCkTznQL2VJYNwnqy030Ms4vJmjNgzE6w9L5+/ECYosvkT9esNyIiRZwkLcd7AxmXc6tP
T9wj0Ysw9af6Ag1CInwXdqsfvk+/JXOkYJfacvA+RH7X1Ue6PQuTbro7w5pwBFq9Z/gjBC96nMWW
E9XlRXj1jkMhSSNFHTTnbW7n1hyx1YOSxoBYTQHOYBNo5kuqPVx/W35lbOyybFBqC2cQnYsACHuQ
7FguMx9jJ+hnhOAqpu39+wc9iHq/s72lQvTLvJqeFsKYrHJ65IJddFB5MSRlDlhLs+9c0Q+pF029
8iznKq9AxuIh+BwNmioEEkzUYId9/jgNZE9QrNGo64Pl69Mfxmjdu/Ez1/kNGjYNHycsl0IYgDw8
TGG5SDRahJW00h5r4LLiRHRxC3yo/jAPI7nXzzSUUlNlguAlmkMb3X1I2W0I+BAT2lDGZEqcyew6
9yosfArhRQhU8c6SH08d1s0TmdbonYvLg+GiiBueKrYSogutfEKZk/bd0047m7v8IkW7M4jgqT61
SOS2hKTIn6RPLXCQ1Ul4vADEpE6GkG9rtb5xWObvyG591+QW6njvpyKMslFCpBE+3I5d5VxHPu7i
TRsMg6dfApMQvsOaQitSMDOnEX/Tl+sVqC6wezcHlSwS253l3yJw+2vHOdr9Y9lYMBSvGJ5U7O3M
yyVNjWZN1/AXjQAfSARi9J/j9jEXaeCqahtOlAuwyqyIJtJZMkaKA6H5q4JxSrrCuRX6um2elDzk
pdjKvARNxucBfiWAjF+zbD35LSyOz41JUoPnsAQWzfXeW4d8OdLNuy9VAZevm+urMhhleg8byx1H
RKzTTri7K+Q6O2cLXjJ45v7sdUZ64KMzXkVSejqEuaWJ5P4Xa8SZzlpJkcLZ6272PxEGERX0AyrN
NYq1it+cAQNlpojlqm3PrprbxIlI3d2wV63tj5eSyLHN1NtP5FXY1fH+oPgqI5LpmPcMnZpatWMg
rnsE8mJ49J8Qqak2PAnWYoHFIHKClJFAsUThGVOy2t7UloJsOhdq/GQI5PG9BPsufAEw097vKFry
1fwtCjCZpd4RRbX394HNOXuByW29Vx7dFneuGU9LZSku/0yU0Z89ryJzNTyb42UB/fhcUzvqUXMo
0r7woR+M88aRWX5Poqh5v2AVcDMbbGvQiwFzV/XJvHB0vBYprdl07noIzmtFTGwhcLCg1UL1ww+8
OorxpKkcLlB2wf847hgZSUyMjx8IYT+6FQn6LBXAzmJma+22Xm0ey7n0Xr22eHeYJ3aEC2ln5Hui
cLjIEtb9GFGDJTUGk5fSQoA6bmdJ1ADnTs/pe3r8WVJvothrwr+Q3zx3F/ekHD/2SMrfrLDcgEqJ
Vd6JGKFpXWZ/EXdaJbbhTS7krHA1h5eS+UIU6eKG3xP/iNvIhqu8+nBGPJza/h7lcr2QbT/nqTCK
9j8uMAfwJ8ZuaJXmVsZ/Gfwl0UL6Fv6r+qAdoMbBYLIN3EfDVjZYtrP0KJ93N9Zq9JeGpCAWpL0L
cljj5v0dnSbvpLDOzXWpE2evPIjLm+bVVzF190eaFy/ofJ11tXTk+ea0+I39Jr8sQSXpjqhJ6t3x
kmhw/DVSL/YD0j4AGSpm5Oshx2dv32tBiMDKhq8S/F9PQeRNicm2JQBhKILpmXcYr7Fo0AV4SfuO
o1jJ6poeCvI6shXUW6Bb8FbC/byxw7ltvDYwIe3XcrlsR8AXn5v6hXH3PYNPMlQsoo3KYZ+rbPZU
cwLoJNURzJrCCvgDFUx+Aq39e068EXLUlXK0utKN+r1aBeNHoUzjmUYssM2R+CMDz2b9+Zw6TIum
s46C+Rh0wkIcN45n6J/mN/ToJWHohoBiLe7+W7g0YcICIqqOsRpoFqD6M3iEIiSxUqjpksvrqbpV
m+2bFHGK02eROevDcns9hjlaBmL1XBvJSaKAm9ULaT7sl7iIxfp0pfHMEtfk5K9gMIc/MlkdtlE1
YYDKP12jHPkAX8kWDsa03mZUNp+mBUFa/1FX1HBSQvLoJ+R1rr/Q7x5djp+bM9D/1gqOFHp2T+ru
eUxCDVV+xs75DmTJyPMt4mfoYlx6EqvhkgKZzc8pbCZSCwPw3C6DUZr/XYdQsi3IDTjy6PBXEVcK
wpqF9XZr+uJTmDGPP+JfkYNN66XXDd5CL66dn0b94+P3s5OCle/bFDn40Z1fu2n/F167Zy/VeLx9
pBZ14kTkieRs3EeqmCITu7Xe0fGXY9q1bGc3uefe+1JH9kCkOMO2JRTMnXtJWpaotPF9P3QbDjOf
HVD/Rp54hdwDNjvZvC07JeJes2bbhAVt/k1Ew0IFwOdahnVGSS8ttuAkXBSPsoLpqOlJPxzllLF9
SaHZhJZx+auNw3LlQX6mU9jAYpo/yDVuNFMV/B5y+rDRo7F3cYYjKoR3EtKvW+tMbQrBGF0fDV2Q
eY+IuVLGd2hzCdnATC85xNyorn6Isuex65YbrRX2jmKDR0VcNI0zReUFsn5GwwvHrzHMkCOvyVtT
prqbaY5eadj9f4Fgm9usqbCrjJsZ8pKGrwtxSgS99cBqDltK8V7n/PZeRhvS9ppoDQhOFoZSrjM4
Jw8vLuMfP94Zx1iVSkcyWB8sx+XNXKHitg7ouufFD5KgH39s/6S78mnfcZeIcmpDbtcKW8fkeH4u
rVQJ2DJxX7TcRsw4aafyXtXjtglzaGvpQV4cEDMaMCb1BAqrXk3OPHY8OfqnAxTqE2s5Pk1vMLMe
/IhvR056g57T5XO4gxFa7errbz7itBWiOcDjEmrFU1BH4HsPMZC+bdypyzE7bQN9cnbdE6fVgLQm
m96cPZoKX+OyFa4VqB/RiAFwYX3oNfTduIlLmeto/XnkHDZVfmiAi/mTWOHHvLIQXwGshT4yu+UC
48RKOJzM/yhsxPizgkgY/IrjM0bsAkPKu96Dlwr80StBkk6ObqPs6zjUDy7ugBiKtC2MGuivGMJr
3is/zidA8VVMhRLPUtLQbg4HEvdq8XjZ1rQbP0M3zC0g0NnXxeZEUoxudWDHxE1RKfzVR/4BwjNh
1/V5GLOzDdgT1j16RYWNrxp7iPwz21gS3puKJib+uQqG7IaCLR3ZM2o5WLkFvRAEbO7k+JQ5UprJ
9sLh1FYl0lSz6SZpNL1XK7UvqzGBqP1coyb2uryXSIXUVk3XiooAlt7Z0QHuPeGbRLMyQGdtp/Vi
KhwhsZ/GgZpqwj7Z8jCjUCvw7TljNMxuUUv/wK641n1pIMiD7MAq52LKU4kkJHryAbQAOBY03YgO
T7pBgXjuaNs6eG5cs3xdgtrp34L9xUV5qkpGh71Q0FhSeWLAb+MBxAHzNKE5bCbKJ/W4f/aA3/Q/
mHHQgg30DGEaTEf6sv5QSNWruuSBV/CRICkhJ1IZ9RQHPl9R5R5qpWG8lY4cBMYgHKisNn8O40Nk
ULBA9yYfHUwk6kRmjL7iqGua5nTOmmVFLy2OmIJ5kjJSlWA/zUcl/s2YonKqe1sArBWv37Bl7iB3
6joPw6fZVAfE6CSdy4oB6HtRp4AkTe6SxVWZXQbkYoKcURMcNFgtEqjvS0X25LElltka6qoe1GyJ
mCaL/JjjGn0D9P5aYxPeaN9dGfqQ2EFYRhxqFfYuazqSjDgQsjg7Wh5Nqomo4ubSJCZerNIh5I15
IW4C9xIO60bqOWPfpexs0f54jMJqhdTPPHDzK2NIIJvgUT0TFjOE8HTIw5sYi7cS7shHkR1ZaN0N
cScps26xFebcRkn4Yu0XEAqclBcST2bG6WauUpDOBP8BmX47N95VJpHOmkB9iHXCpXoUlig1Wowi
q7fLX7HC9i3wrvp6R2HG4AOSe3h9ZvML2BXebcuSRZreie9Aaue/8HVyHK81PqxzvLqrZMKNjIIc
6raXzbghfZeaoLpiHdXe8qiAAQlfkn7fRAQ8n8bHi180mP0jo4+PZ9aPlIORWNqugBwfgPm4unpF
UoHC27WITq6GezSImcN2e50bJhUxjh0iuPapY9cSRYMERylTNBiLLVP7Qwi27qDOKEtrAvLpcFv/
GG/8Xf7XK7kLe0PICCnsqLKSFAILS+3sGx+w2C2Se9Efe5bIwcgDpp7X5LiNqgPsHWM6e9Pr5QNa
79fK6dPmGpCQg/jPLunhB6i2DLap56VV8ubf2cKqxFW7c4n6rR7DyS1Bc4uriHQnz7kpWX/dZHCr
mO6/ye2wQUcO7vgSFvG58ZJBScJBO793dmS8WyUAYbGt5T2E/RBpL4ypdfsOP3rlZ+XLFPbIjQvk
E+1sCgUzA0rrlj5tuG2a1gS2J8WE35KVP3YuXa7EWmIKMxGd1WOH7HM0NuiWmyzEfgta90mjIqsj
piFGHOU2k8KOdXF78Oyhw0+2cPn95iHyUQXuOv6w6HgyswNYjyZF1WRsBejRUmV3iZrMfsX8Nb0D
R0ffNvrM7gX4eKors2AwmPtvCpPnmIrPp48OFqOvtr/iSd8TqBEiFKYGXI2lgOgVEP0RNImUkR8K
Fm5DVekcMdJZkhSiuf7tUbBPeODpu+WGJ1OYuS4Ga4nqFsl9G6stV3lPfultRWU0Ob38Ko26Dcx2
eRG2gi5wANfNaLOF1mUMgtrxdYm2yUMkPVbwvSQasQdgTiWTZ6HDhuU8LxEoHz7CZAcu9kFdym3f
3BIM/2WOX05dnrMHbIoSufbq5NANzIZSQvqgiabkX7V6/UQHSHoTpYDlXbIxK7aZoF7UxceLQFs+
hCcaezL2PKyrcHeyZreAXrpII3whBAMOSbbPtLZsRb2R36zr9EkTNGwIeM21Vo6wqS7QnZvEBzNZ
K2dEDtjAcIsxlciZrZNJxfmvJI5ztoW0gdkq3XlpAKw0JluWia2cPgogv2mW7IZJxDN9zII5MQPA
Kmd+8QECSsA9Y7xpOahVDF35+5NvK0A6vtMYSz5AC1TjmKoe6S8hQq696EM/NQOg74l4vttqatzA
3YHwR1YD23YXvI2mY6AUbFLf52aaWeqSs9jpGAw2XUb/Vr9N5b3hYGcWSyHMPL1bL0wmS3v/jPkA
yHjxuNdr/kSjVWnkY96oRqnZLVxQuDx/Co9p+k8ITgMPdyXId59cmN5BLmsnFYIcwnKZLMSNkfS3
ZbAxRxtIeqvLdNf7ccvBvO/Gb8MyCCGprDAi1hChtKNFQRDYG7NoFijRZF9EEfph0mtDW5KgrTuf
Ss7+JkS9qJ72t7wqi0aFnjZ/MbvqdlMqMAIIl77ntlt4OceCu4aGn0j9xVOX+hQhmbgkvxGTyChb
ccp4s8rHBzhcB5gwhh4WO23v1/72+QjFhumjo76xAzCO4cLEKzF65tI9LMnXmYm8oxuFLsE4DxeJ
hpi1QCz27b2lXKHdW3TxbU2SvVyhsn2/+rqPMRfTNcYQfozeC1DdjteQvyLflYYyGI8R+LzB9qyG
SfrkWGpZdQaHg82d6HSwiiceR6+Qjq6H9hou2fQMisq5PZ6WHXtwwACd1s5D2Bx8Ie5QyLExtVWh
IQxdYK2eKpZYl/n94jRm2JXJCcUStl64zEfNF6J5P7VG3zlDOpM//OB+1TT5nquNY4HDbAnT/CFP
MBF00sZNc5CoPCpDQN348neKdyKWSK1BF2q+DCQ52zqrbUcYMd48ZZ7G8tDrbA2PRcLSRVKbiuOt
GpGpOtXvq1Q+fMkLkSiDdmzjGt/3vIfBM/JFjPjqag0Alwbsu58I+gb+Mb0BMjNLPlAn9eXKUqOD
ACrC9fj5Tl0Gdt7LFd/qtlExxlUhYbrN7H9Q3nKaG+9yeB//FEpjOk++rmeZmhWbUiEwlNmT/2r8
/G1gCkD7DT7rbfEUvKJPOlhCabuG8Ylp0a91S/gRXPNQcLKVhWA0U4L30fc4+D2aM3FZ0IzEDTx9
csaTmWvXuAH3rWh9dgxPipP9WZSmF6rU+3TGFEA9NjM44VPJnV6+C0GfYkf8yU9wo9LtyzCaLFUP
Hi+dBKCulT9xbgUt6a7SGGDC5ISpj0tW/XVGsOHQNyeQ+draC+cVNcvgAZ04JPTHcibnq0+jlafI
M6Abb7PaC6KfZJlQOXO7+AWSJW/RrqfbTTre4BIg+Kmant9gvs77CSkhYxt7xeviOAIZIQIHlcYx
2b7vPfsQa9MVHx8QVTnyf+E8AKmhQImBhNlqBYKxpd1auO/Mc70TO0raO0YJLZR496qOcUzC5OpW
3mG9iTcRrH1iOmVdMGxYG3/TT7mq+JCN5PdqOesTuLt/leyjqVoUBiEsVCx4V6PDYCluhrpvqq7Z
rmnWdUsW6NxpXmQw6q3/2jO6bPUiflGO9tnA7jkMROxrb9V6Oor+gs+z0mgLnV7dEDK/HHnPLuYw
XK3pmX7G+Pupq3gCUOhyRt1pysEdlG/IPIKEMb1BTiYv8apEz42BVd+BiYc6DqhkIZDGgm5V0+XX
bWeklfR8CycRQFtZ1ajxCIhDYiCi5l4eLFflSx8mcbKlECA8859g5BpgOXxIJtASsvpENsOaCUeF
zEFGZSCNx2mmYqTDSOd5INe3O21SahE8bbXoMHxDONxyqSrvAnGLufanhn86gJRdizTSIIlmKi1S
obeMDCe/sOqNQ/y3pHMmXN6Zp7I78e5BJogN0t482vJdsMcHP+giTpkGGbl3Fb4KGztFo2dMw8CE
5dkgIXntzMR6qozMaAzUpR+/QUPC0GlsLt3gsYzmiJQruG7jQFANa+VPSMFfr7rMKKZf7h8cJS6X
zAB+IJpa5QXbB4YVALmKNjHf54kb2xQeRFTZj166lERVvqZoyhTEU7QzjTyigU55JbSxglPiCIxE
8YSbExsfZryeW+6Zynh5AjOyK/ct/3fVfgCyblHTWkyecYveC0MUPKs7ZK4V+GqDBmRDMftYIA/5
912vOBZFETeOCPsp7CjsIznqEc8W9rG3bjRhQsLlxPj9e1kNqc9Wz2S7GaQXS4F3AxQxCNcv2ov0
JRKNG1YXBR6jHOjQemArlGbnVLVFZ3WRSNSJfLLxiYbeeOa42fuNwD583GjuU/gi7swCY8U4N2Ht
b2dOwKYGrw8ZicNDA69fw+NHrF2piI/n4YxYso2XLCjdvXzktkj7ME8gG9GEAd7SncNV8AQAesKm
hXfSmMcaZoyh5kMGloI/QqVPEs81gpwoSQ1r053BZGgGNIt/Fx0h4jOJZA+xY7LjqtkcTA3WcbvD
ztaD7H1cGxprqsRJ57iBVm8/mpnuIbfAyEFdXkIT+T7xddKGc1X9iR7W10CLtA4nozWR6r7N8YS5
TDxQeILgGmyEjiLHsS5pPO7oGKNAst6T9l7x51rU4ijtBjQKaYahAgpGNHIxW06bhsSgLBYAVTgw
CEuiCyPIAwjr5G0J1MYiC8YDxS9Yu+n6drdEv1BknHzYUQUHJPhUxnLkdbA+lyegfp+47VVzvIum
Od7vRBPz7A6UztU+pUgqW4fNiDaOhSd9CnGK8YbNsAS5hw29HuQpgavNd3KcBGGC5jW9jj82E4q5
MSjyBJtGvoV7hEvApX7E5Ys9EjyfOS2tCJGaxUXYP1qUkijf9CfQQMbORLaCumPVSt5oBBkM2CEC
B006dJWHMPiOiTlpLHsAodU95Nm5SmRiTXTq2LsPKlK97AndaPYc2DpXxRzB3Psm2AafjwAozhVj
r2t10E5+zChooOlyjoL78aUpDzGzoWqLMvC4opSFGo2UlEZV6kSoTfHWiY4V9hgTzsIFd/jd9Dco
bWiMYgNeRFfCbfFvMjUFx8euGpEJC9j+pkJojPTUn2BHagdFIPjyaC+V5l5rdoWgws7Wot4LlhsS
+NAAWDMNj7YYfyIx28FBmcsCJ2rUdvU9TN2tNWgGUdxKMHGMuSyEGdeJgs6Vmi6QrhkT+G7ma+Ka
sdEyru1MhXTL8fPPmZ0pYlZ+MiYRofjGhJq3LjUPBiCSg53WJfjFGWTxgWF9CGOcqx1hZH9KOcfv
1be+HSh2U0wymvslmN/xjAu2HPvjuWIzoC97KwX6tH+Wxw69PdUynrf3h9XI9YGEU8xHgg6onIh5
0+wM4ff1T+NaZnvb7zs9iEDfqQ/ki3aUdbEC4RSe8wcqq3927F/fvcOagHsDCkK52s99YIG9coY2
YAW487gXbKMyS4BpflKvUGWQYYdK/N7bhli/iN+55F9vxiCVlVvBWRJE5QzinINF9En5Z7Gx1vFn
RcUGU2kB65RU2A098g1KvT3EiyBq4BDYgukbEpiy/wt5F6i7K50sHSVHQ112g/P57xQ7MC4zgnFD
1h4lP8ftIfDfehwu6SfGFnHTCmS0Ty8TRn7iEjhQGP72i6eQvYsamuf5t0+e5c7eTNUkIivXhFc1
uY+0r3YYoSzX46UFaeboYZFZqHf39tcTuSl4D98DqNwKGtn5w1oa9v9MqVSGfImGNLpmHruzfigs
SFWR61TnHw0u9dPk69sdfPh3lo04PKcUK0CZUQtVjffrFzFXuXrrdzRyIbQPeHahlNuv7i7p/Ahy
HaQzJrHfrKipXjcXPpsjL/cGD84A0BOG3y1CS6es4FIrcduJbbK+/pNKaPb6r/rJHdvYfa22hm8M
Y9pC5a4M2TOYfTPb7LsVamvMo4/nR/lcfjKPH2PXu3wvqX7nSK+GK1iAFVCF00qAbjG4E0NN4LER
/AG+0sczXd2IkyQj1cJrjfV3Z/X31aZqVKKfD+Ni2S527qK3D1d9wmg8WBAaTTUI1/4HTi1ptPG3
Wl9a4utXRrBGfrqxSqWXU8q+7wF+jQVDAwiYqyo9c6TUZ2f29e7ddQpX06nsDQF2N7hiOrLp+PfS
JcB8oZbvZVZTiGbzN+DW2XGgEmEFuVODZDfQVTPCnIo3nR26WUURKkr8sW4VAbIzEbkQzTaKhoB1
BvY12npQ6d9y+DHkeKAcgUymb6JnXF8NzimqBJ2buM4dWljmCwgt0RHZgHnvozdx9NEV2coY60++
E477NBBwgV63pJix/zvJ925IojRKKHo0aTy8qDwqiaPt6mSbC2ZmleCrpffpQqI3+owopr0Libfi
27bUCfFBwDw+rEfGi7X79tK57pCgjCr/o9wv2vwSVNO3IW4KNVeW6XX2MtzKESQIr62gawnHmU1I
YeO1i9nQSgxBXD+qgDO3dnkzyJrNrWvTbXASkUf9RkV98CL3jwlIw6BojQ3o7EvKGx3ZIk5vAcpk
5lvw0eyLyOp/w8hk+3ZHu2q1gqwo6cvSCeS8lWKv0HR0MQki79lWIsuIK8Twoy9km9CiKOjB+Jvw
HAZU9GVrr+rBjNDZF+qVWhlB2MJTD9wypbIl3IqVRta4OdmNScUWyJv3eY8i+5qh/B1wjpkFcQy+
ciwCNsI/cALhHENAg1H5roAaFMvLc/B2DtTXVOqZVRgH2AlNgi11pQU0O6OLsLBO8nMP8RaCVHcA
VgqEX6EW0Ei+g2os0NdSeFps17vC6QwngDARPAgFkAq+vUaj8yCmanA/ssZXH1MwCzCDq41zOaYU
BJlDhjoG1SqBfRM0jBAsV/Op8Yvj+n3JqSeBNCPrVkpYY58EGxlxTVvAfOg+hvzLtffuyip/ls41
1TD/noRk0iHrCQV/GfJs2BzkPogsB/h9TXOESZ9yQ3BGRx5hXTlgjWVXhnz9rYYAyhnyD/+1PoRt
vuxoId4OXQzCc2NiF49HpbaO5qLGzl3ESSuoDORAGa5MKOVZ1zqeS+FfFdMK+A93SriERGNXlS8k
AWNGR7tR9cvOQ7LDUlhaiatMu/tRm7Mi4Y5C2oHrpdVZgxSU8DVDC2aRjUvRIbQPcz0UQbrfiZ2V
vLrUwzhQokrYdl2N95nDAiJITRqgNdy16ozVwVX4nLXfEcB9QTz/cMNrk1WKR1Cb1yh8vkRhsLeZ
TEFsc0Kim46EviWv2cfG73aJ8+OPPDcrlSKVbnKFq2BA+hKTtXbjjlVls1wnX8NdjrICnkgZJ9Gi
gBj4EcPOfIXNUZtjekV0zH8E0h4cVVXAkwe0DWTTkbiL9E1Y+ItoIoLUXVFckLGpB8fLhtG9P8sp
EkIoSJSfV4ZerYHo0tcCU/8xbJt9O2TV5XDPXl5FkbQrQI4bKjlScYakJzzlK5tuuLDue7EFWX22
DwAiorGigE31k3YQuCVtJGw9Q/ZFSGH7qdpK2rPFyR/cZTxs78GutDPSWum4xLf2CUrIL4IYJeDc
h4CveDleyOACD+U6rB8kOsYJ4nxpUOgmdRGaISOrPklS0I6Dh4+kUjpiuE1hVBJXGKvQbbSDvxUI
VfPM9llAdLZMltr9k37Tzy1HnPY2z3LetYK1bUbO4WDl0knfhArysL7OdBI5/MEsbH3bkamaKxWz
OIqXOVGGSAfDNK0q+K8jSkUeUNzgvljNb7/9sEoSkWk6DltAmCv9GlakB/PgoaHdjAvDsAXjb0NV
T3YoLDQKT/O/fpx3V8TQHBh7uhj56gcc5UpDjfzzPQBXU3e83Phj1e6krW/QUJfDk9593588AONL
s3E1KRMQr4UffYQeNSubWfV+VOejW1y26UizpHMdos81U5u/EXz9djcEtsBYVwQl3xZWH4DVZ/WY
n5WhYJxWhn6UlQOjFgs9/X3qmMKCRELusb4pIZnFnicTyS/oK8d5yqi3Q2je5CfG5p7ThwksUOX9
ENtS458xooUsN/kTUVuPxt1MXnie2E/HPN1tgQB+a0TBFUpOJ5dCyF9xpppr8H/IvelSo6aleyVV
uZFgZ2ZW3Vw3kPJHlA6Xl76Fut2woB60V+0uPyLCCadM3Z8h3/PPAxclXmcQIi9+NoG2xDyCQQId
T/5kSQxvHzeLvh5Ow/eWByRSKZsnRDo6XbtBqcy5LdNLDscQo83i4ybXIkuUZ7mfKslAFje1sGnx
8alhFaI7PI79zkpf8dOCh0AEDCgli3YNMOGNvHWGaMnGu50PNyd/p/JBS5vKJeKhVF8q0qqzBR1C
iknMfLjd69QWPFbxcRhNt+Tv2J2WjsVbA7zirqpXI7iNEpTRQGLqZrwgavdMkB/d7vbXjK7qgJOC
bKkQLQN8ZwvKi1RQWWa/eGloMbZKV+QWzyg9zmdZnCATpnWKLuG65em9LE0Nn2bZ+cV1IeUXg1d+
KA9Z8A1+yba4LF9gk1yptQbEN8q8ukeXnKHHe1exI5KFsbIT27HG6ePJp8P6TaT/h9EOoYHtaceI
kH2lGJujkfHx9yzGWOE02yyK7gNTQiGJlENGaR5W+XSZ6/4vlyC9fcBWQudOL2jOTCsiRZDw3hLh
8C3sUa/yHnjgAKxu8M67VFyddLTuUQDQqtK3Y3RPlbcE149BTZZHpaQCZdkuCcuhPkEeCJgs6eE0
e2h5963MsVF+765VvPAI5b8IpseXT7D3dRKADfpNMXuQQz4pOeZcILgWEuN9NFVj3tI1tKLVVFgp
oOzx6rvXo+dqiQJSOn9ijARrMwkm8Ux5aArP/8xnRDp09SVt7bfoJHRW7S1Zn8+scQqj6LDDujp0
Xqq0g/7ih52ffGPS4o/gK3ovXidW2pxerYZ7a5Be/92RQ7dvBbJ3p7+ZHwZp4l8d91HcyOaqz13J
gxOF6eTswGEnRPy98gRt5juFDT9VMsFh1pwvfMiyuTybSlhv40gTWb1xvEl4DFEtSNjKLdTb/sv6
svAsFx62N43iGSeLIsuvjyzu2zLlBvTEEecuWCkTwPoDMAs4GvYiuXItdbsqKZPBBRhicO/MDkG4
mQWCr/tu3u15QAh9hWY6RHs9sK+03E/ylODwoC8KL3Kajh8jDkXBH/kVkAE6tYIQr+eASjQmHcfI
4GfGV34sMs9+fRlMnXFbCKETMzdTna5DQIFkt5nSue4RCIoyzyXeLRDpIIrmL0gI1I+vxe8G8S9b
ziwv7ToCo+Awed3xLBTovbbzx04//5ZBbyPscJlNVnkCcajSpunO0srmDIVwNnY7cETux2MmkPna
x0ACkdqgB3nRcHbams3IggykzyuDbddXcxsTHB+PCxKM6yZuLRfIzRLPcVOYQCzecPBN7yg94gF+
tIbELiYQkRrafXqF7AFP1zhK6lWFwTQ9Eetwt2K+FYtiVLuKi7YBE1BoYbsU+o6Arrbu1cWRAc0F
csBCt1qIlYMivhXa2xDx3ZVD5AbI87Nv7Nxc69AzP4l7C7LCnkVVVB+uregV/f2w/fzRc21UwC/C
RCL62gNJIVE9pIrojfUnYnczVTLe6WxF5LqXRjVgwXLW3IrXMcm6Ngf+QorE3CyFIRWdcXYlFGcd
HD0fSc0OUQhlajD4Ac8+1M/XNFGsdXIzzxTQvONUXDZonrqd1wZdTypgwsfHH7lBdqXBo8ha0yhy
unqrkh5BAkAA1TEnFaPtYKLo4nKmIc4xtgN7UZoFlMNuZAA3O5PxGMDo7TSL0Uo5bxWtc0KpYt5K
FMrH5a/AsFzLRyrtxtxp74qEWgqgMY96TvKaDpBNiT4Bq0YL+1EuIwK5yUEihK/jAD2wXxhDNlvr
0Hr6oqcYWARTsg77QYajpb7Ck4ZUKlZXOXEkLkM58aQXvKTeX6NcseLr3KRkvrDUgP7tlkpYr4Uw
3TofWgdoCRYgZjCRMLrW1SaGMsLWOYw6ANqEh93ELKj0C6jOdGj2liBwhrHHjmwcBO0Xec2ZMfsF
qgbrkISvHBU5EkMo/aKqAfps+4JmN1c2OXKlA2pX372kZ5xk8rO/AAkAKQ6G2ePM5Sroe3HtnLv4
rWagTQ2P+bI7DG2fBLtDJ9thek/zpBW7/QzYpOUf86/ZhFjXOXjBZwj4SLPcnvzOu9EgloMF9ML2
YUffC3lNy7V3gfz1lAu4EpPHIGgxT0hgGp+2gS1ClohiePPF6UnOaeWxwzvUumDPSoPXnvjEo3WC
kjtChhbiokM21Ggt9ES0Kt6QbDXXj/AV5jk2i4KP6D79zDZFjp+czaCDAKIicsDfcJRecg4bNzxH
7IxW0L7yHXvcISd7Bv6WQb/eWmkb3w4SkM4tobkqejmofPn2HxHeRxqWn5jR7SK3shXG7woQM+OB
QFT2iy9Xs4276ePpMZkNefBr0dQCb2dg9mlxFVzWrg+eTAAY2SN4BMtgz8IELQt/2r3L24HjFh2v
kHOknYo2TT8ywC1tizMBJVvl1tXMzN6uUsA9PrV9qW8/JHGoGggxGMKMPDCs6l8vCOUR7O29iM25
v6vVlYsG2a6UINB6KwyKikZ5fh7t2cpnjjL6924TXuxqXA+IF+CwtVGsOE2jWUvRBHOBBn7vUo3C
Vgryav7qeDrX9Mj2N6M8SanoqS18CU37/Bb3mmj7hnW4B/A4XTjKLRPzb8wlwR+O7lYKMQejLUJb
IQzl27Msr2cTbZnbBHKX0/+wkJLQm3i+61VGOYCiWToA6YPS6lOrQDMQQrArDZMGRXUxhvQGdZxD
qUU/Y3taXWOz4xw9vmMF7uHKk6f546m/7tM8EKyH4agU8GAyE/1usI1DK7rKB704uIsvhfsVmRH1
TYeVbmeAkIQMX1aSUENnQ4TBmo0o7c2T3fJltHCa5xsIwbVjwzzRQwu+tkzZchOZv6oT8V1IktjT
vqH2UNEzZIMLvhvf2RP1+IqBeV7+rpvqJRYQdJZwvUo15cIZMM0DnRlCdivZ3+2m+4t3SI8x/oYm
NVUE9SPLuWPKpAYqg21CRpVtIP26JHbDTImFYr7hi5XZus4O6DlfQDuzw0tsiZGXMuM6T21w6z1U
CVuC67g3RJE9CPVaxiFlJsQAF11usSSXiMx0lLlQN1pvgkxuX8zX4wgGf4c5e6bkGTgWYSzWG8/E
lrK4APuzmtLnTZtKNZVgYsj1IsMB8ldoBl8esbOBzXSl6xAl6sr7GDpJQokyZHSGMOnL1rBYqj38
iq0PTaTt+gW2o8dNItQrxoGVn+WW8BH+VMYpYmZYv1f6aLEk4qR/h+z5iE5Pek5tEiK5cz7G2IYM
tLyRCkyLs9b58OzZcpXAXtYIwxt1SM4q8eXGeqkXmC9UU6o9FMGgYEEcUYf//gbJ3IjFHig5MGZe
9EW+pS/5XYgFHngiQ649pkbOoRjm58b9IUj+YoiKiwaXrMwUGLoCeZHiN55Sd0UYdfK8KLBtRP8C
B3j5+j1ppADr0ArjOL3WjNHrTaQfpZrfhaj0b/Kx/MJ9Ra29Gy56Hbg4ljb8kdjakUJ97cg9kaWX
o0WyQz6WfmDgIH8VMZwWxkiWsxqUqqfLf4wPla1kxtFH8k719K61cFdIdRXItAN4uJwli5iDLWse
YeShVgkb3H6QxC/TZcw7TB0pvoHiYeDyOUUuMdQW1/yAosr2YR8+KS5Vq/KrfKxF0MFdC9AaWGFT
AMWYr4w83cUFBg4uX0dbkgfusFN9o+7RIJobGQoRYijoXRnclgUgg181FWuqYd8E4nV4AL4LDESY
OdSBtiE5UdkGfPw0LLQUlbr3R7Xel3WPutuU2KqXVZAl4CSQ/P3BCQpqsDcuXr2Usj6ACjXt96Ld
EO/rHRa8B/MfFB2mqEYulPavL4VSEXxrXX10iPb7VOaRehqkTasysjnKv3v4CtY3MFTMMuIlau3V
tVkdDzifDAqqV7KpNnkZK8t/LrFq0h/nBXQfRoBK30kJ3MURVNBW0x/ybezHCTLVVzpZzJuETJO7
lzq3nlDkzp7KyeWJuusZjxiNNFcMk7MEkV5W/MH0cJqvXVFIfBUudD6ZNQ0h7PqMX6Y/mOH08VBC
eGzBdrFK2HgtlY/AACAjZtxzmYyiWSH3vUXptiK1BZPzBbmBijajShIdBOt24DyCMnzaIibp09lA
zkza/E1GIXCuJRKZbZy8P2f01wO2QzyG2BlPwhc0xSMrGtITI+mpA+ZiNXR/LipWvHRAHlMN1aEz
U4PDd03mfJXT33g8u/NaApfkaJ7PNSLs7rZY0zsV3jwp7pA2R+vUHml8eCS1SpCp5VQd7eIB0rWf
x03IzQ3cS24qOfeQ4lIVqhwOsmTP3f3tvfHT0ZFZ8hgdjsUXofCG+EsU85yX0Pig8AHWsMZWZEA0
sOtTxou+m1gU2W2cZs+ujMqxodImDdCyvQFp5u7NSLBD0sjoeG56wuD5z0Y8e5dPXwI0IkQ39x8D
ecutvauZOpomExOxSL3or9uVtjuTAU8Kis6tEsDHEj1npx6ro97ip8I5NvF+/f339VgJJ32GZY6t
QQQb1UbiGtsG71iP1337e3HVoQWnSMWlIbtxCj9oSNyK8JXmELJOIrJIBLrSgRaWcfbZ5lU/BIG5
yjagAJqvIs3qcIa9tub9sENYEvNuGhkE1E8Bbrxh8mEKExy9DBWTSVnCtIZJ1FihqiytF3WEZMDE
9c05+W4AzzaIGPv42s37qGqgX9jzrKMMGU8TOF5Z252s0no12zRFi40LHUO5S/hX6C0PaX3TvHf+
gTuKdxS1zjj7eJz3GYiq2BQYpZVDyp9afvABXMQL8fm8kKcCNyCeGesZto8Ln1WX8GG1piT8a+vO
YXROIWvR3u9rIlh5kydCHs0cXHLPKVIvI1/MSm149m/VUHJUgMo4ipL9uKo9fSDQ0LRc1oJN5uDu
4J2y6kc9Zi2ocUNfAZxSm02GJ5CrXuQQTJEWXqTpwvI+Gyy8+R3495LJJ5gZmL856qSvYVchdHgx
4uuBOMhJLSInkulhuwWw5o/neBRK/KAb8IctRBxbcLF7g/J+9GWjFoDG6BWUiE+M4TAIKUQS+5b7
48souVlwGfxKp+a/iDVzsETbusO1FBlnV/gW+j8C588hr+zFhrWHJdWoRY+CGgCI1jGtYM3tG4aU
PueR6TMz1itMmtvqKBKcsy/CmTbnjg/tLzhuhIBhSc6PFlygdMJ0PkvJgdyGb9+lPXWb/XTBzi8R
xUmrJNoIYQQKBHDbK+1X4TMZNBi8NDuISJ1Vq3j65tkNgSMDRTDsJrkDUQGD0xJq+S0NXJ24jVvF
f5YWFj1FqLJwcf8UPV0FF1ypxd/Yk67zu3v/5vJu6nWUiNjqymcff0wPhLAaBYo+7lCvt13bpmFo
VbpWugQMqPcnAhwD5m6CatKAeXg/sinz46UgkubXi0ImaSSl3mEVCErNm5CBqWSfsZy3yV6i81Qw
V9yFn/0s+dwG/LD4EX6FLO/XTVKJDml3HgugnpSluwn1Tmi11tCMhgzPP4POX8oqEXsqpqYzJbau
jkSv5q35kbtLVK27NyyWS3hl6evULrp8nQlaOosCIlmOM7I5hZg9uPPBii3oywPR2vadl3t0UFz+
m6nChQ4nIy22c2KJhP/kOsFSJd7qiooA1kM4nOudWRc0BVV5+8kE567opdgdHzfGf+b12gVQOgC3
zO+WQd6KeiBIgaqRlkh3iDGXmpYnvqZg4XsW0Kq25G92y2/YKEz1arBG6uTqO+PQVVjDsnHFS2j7
ogQeaT37TBrBAPL67gyNCNF+q9rjUU1cM54lEGZ/cyc/KRHU1ZeYIoshLq/HAxUgnG0CBvjFcBDy
TBH57vsRwhIpRsBCk662+xrdD2GHx4KH7dGKXXiedFtovcUvmkHve3CaeJSKBF/fU9GHYDy3d+In
6pfp5ic55q+rU7tKbhMIfdZAIsOpcr5X8EzS+ReDwfLeIzsDZ1Mnsj/DOYtDNYont6RvX4ktcm1y
mfHxAOLBDKF88b2qVkrJVaxFipk+IYP4a+srBQjVxTVoUEzCXOWjdauo4FIJTCUgzmhL9So+coVm
2YOO4SbUMouZ/bDKHbZaOH1/ooVhNjZKtYExW+zeUmgzfuQl3KtnGL6R2VUqCmocTbexMZOuvBi8
0qrDaXyEiog73JAn0fLe6x7S53WTuuFcuiha4XaViw43g4tUREo2nzwmGz6sUGor3JnC0K5+RMWM
8Damsg/ZPJ/tjT6qNT9sELA4gCU1AZs7Lgp36EUrfHhM01VGckrD7+Cg47q9OEk1dJZw9ZPAoYkr
Z5MZPUrZCHWyDiN4if1zhEbwTnsIkYlW8clFrpAJQ9hgfCPQttEkJCJ2PjZyY8HHgxe/0Xw61ft+
H5QJIxKAfKwEHnUWsicpJqawJWFbTtcqJinZ7VOnlqskmkGSjzdU203H351ku7V5isEILlxaD9oV
CGT3BYkCZgpu4xBnqCSQ051QetuqisbF6tmEu7BhbZMDWVXtfwrKnYLL1GXrdtmXCsgEFJXfNjef
U9G/t1OQi6wLNVNgfQiSE8LXTvql2+JfSVm+LD21GaeqJpoqHCUPZBvpbANaQIMkFyNTvYkp71WM
cfkqWDgz/B6ZrhNslze8oA1a+D+lxK8JQQqURgujSGInCbSRdE3lPc04zrdQ3Oks7l0rmDBSfg2p
HwGRs1XM8/CkvtvT+Z1fsX5yXfDR72rHrBiECtuafmZtZ7OCfn1dOW8L1fllu5UyL8ARY7Y7BJyT
RJ6X8ZWFXsw1SXprPE/JEu4Ni4CFYzaGIrDjHmnyjf18zgqg5liOcfvHqhJod5LN2Uz/kjLkynnA
tl2iXzxEvI+hPj1ezNkjB+zV7Twm6MtnL51T8z7ZDMPouVMvbT/hGQqVMZYLZyTvGBMKPa7wh2Gg
Jyr0YfC1ZVuZAXo+7LiGyXdhER0u42i1ITATtJAUxnPWPC3VoUfExSoy3zXTF0UlOxlg46bz65gb
3zI/D0baF8hbNIauo4b9nr4sOwovoTzxGyGauva8j5/zETu0I6YQbxBEyTRi2EtEO2fiIqUffDtb
16P/UjhdQAvOUUdtDEx8fM04LPXD6PcUEhQaxYjKBZv/hVUKDj2bA6aGTBLUBB1ztJUs3vUi1Y9/
dR486odBbpH5C+btNWw8WF2JJ5d83W2KBu/qYuybwNytkh/ZmWehmFnqzP4gpFytdQ5cJ/6vupkr
ryh4qixFEMxcSq4OrXIdel6QTpfmA2d5jluu63qOY5s+apvb6bkovefEAh3bSe15WIiNZZGG6NoF
Qp8ru2fqiE8poVKvBtNKGEvLNSbFLQeLWXL0fZFCeX5Y5ZFO37NAD3h0zdXpTuJl2fVE1qbuHABm
KwHnuFCryhyGZiOP5+I2xt67TSwp6N1PQWzjoHX61eqZ+tm+6SBSGkw5FMwSIIuFiGbLxQPeHCLL
/fXz4D8AAdxc2RZO+3uAC5IeE1JhEEYlZ1VMLvVJJPdKbRiQNRxh3C0Di/1wk37c33i9W9C3+3bg
4/vknpD1QOYJH3SQJ/VGSGiHv4kwpxnMgA8U7Oqcfg+JUCEDIN0P6RUnVoTNOfMdsbod3Moy+WZs
qFOfDv48WqWRLn7s/PR1+m8qBpUZGF/egPkmNh3zo+Qr1+a0Kq3kNQsn3y7C8nlWBAd5gq0coBkz
C02cAkn8Vnt+JUgvczPAQZvNIKFjyetW7QafFL+eWOi7Qw03ueimTmBYQPRdLtezFzjlcCrcPRdW
oH9yAG3rQVbLOYPYH3tEF5wCr63jHEJSR7eU2k7M+HT3zJM5Z5UGd6ScFeef4CkvhjSxDfCapj2m
V9nObu6sRMuRXffJ9tXyBdSpv+5mIOtEVF3H7MLyb4hq7D/Ihr+ZvQGIjPOFNtldxCDW5v32qitS
SnMtcf/Z67spdinrjg05J1buUGkWNchbzoOU598Bjd1hBHDfhNzcp4Lhx3kKlb85zqSfJMybpzAG
IdHz2LSPb3CpSaqNM78NY4NmNc6pFbyl1KJbAeA1vKBR6gohOJfzx3boANjt6LJ6NROMklPLJ3l8
gpTFF1DCKZ9AfByi2QzG4Z8SbfqszST49oEecfNdoYSTty9m5RD/j2MdzXhchxlpGoD/AnevzQG+
5trMsAL/Teiy3B9mTpe01MWiIQ7ugGHIpIE8LNbDgTr9pVGkZDojIiyPHRRzy+/7zykwWcbQjDq+
6BHqSRNNlTsHksUjeEBrQPUAJzxn2wizuHp9Y9NRmNE6a/Z+Nlb8GHz9vrHAeq/IgqMjsjNfuirU
PhObQlkrIY/B6iXkCJProRsswysGVYoM9/qIahO4z6BbWyiy76Ouc//inxjSh5mXlk+11z9PLaZh
2+m+cpJrWRwFJ7WX1xXyW3Tu5shiGME6lonx9iRkBMXzg2EjBM8FnlmooatS7GFsvmGsFv30DUn6
TVxAWDqEqRciKX7zahX14FP5B7H7NM60WBzL6s26kG4IKVCpuKiwSsPVljcOErE0fjN7AeMqvuDg
2i61/zRqAVp1xkg7Ng2nwAsKPt3xxBEHoOkuZfVDO8TGZU4bAefslD5FzUl3ZHvahb7Tx56gpwBa
m5kcqjgen2QPz6MsavqFm9QQ9jUM4NLlybFCuOXrfXj97ZClZOCC1QvtOHlc8irQeDGrrp+8T+0a
ujJ2oW2LXDpfEcyZcMrQIpK/XBhCPZLOdvGzMpkh4Q1KTUsQdTc3IgVFSgUbCk4S7a84qR5HH4l+
x/LFdR9dy19mLnKft4RCCCZZMbGITYh1sqZP6or6PbmqW2VP3FK+96ZrRUTc3FeGLOSM2sIs07l2
qu7inP7R050vlD+5Nkw2crjxZWkpdnxVh1jyTdOm9gLW3INDYglGAp0o6prQhM7OgTY0V7zEnqu8
dTuRiuYCX36M8V14ZhDPrF/1e8Z29El3eXH9dU+jVLquu+QH+2vkaRWQzi5hCN3iiBtDH4CsGYf9
u5gWpVJKUzG8cRZf2Gj7rwxo2fZSYqBihQXexSrJywmgZIcIndWF2OIqVuwYwsw382e+BtYH8ATD
zOLIXezFKEImszlsu0y4wVcol9SKz4P45xo74TGgpi8UlqKAO2ONeMjyJjxKxbcvucDgb2Xuihey
tenYgNPBkW1RzjNt5Cr7dDOMwaqZUisc0Km49mruyV+IfpIqYAb3ToE6xHLJnakg3AJg6EmxFWTc
d9wmO80iCDvuI1Jb9hgbhIdELmjpU+iuFZcCk2G1rZf6fB2oWfYO71iqc6t+2WOWt5HAlbOWtn/z
Kj4wHlMhWOU+0l3d66fqYP3gnv3m54VcOZEX3ztcvX5U43g7f8wzoNos6hRx2sww0tNDatIYXwDg
sGXA3WgnLE7ydQMrYTSBMJT3T5JtVTsYaElptePU4jo9rugiEfpTtGxLPSpbSWipp0uOTBPardca
xG3voSb7Q2xnlNPzQ/zZnDBE04JcQToy41qkGHTlRr3hkj4MGzC0KA57WMS/YycmHlSXuBKLLcW6
3U58kAKy8BYijzHCrehrN08GyloE85/5EBkyR3S9iBJQVQJTl+CoTH+21eMbZaEgto2KTjJPa9Gk
Bnx+0hviU1Tyc0Fz/wg/B5ssJSg6fe+C88OlQI+MAZi+kLs85OsdeDwlxd2m8FLc3Hy/6orrWOtt
AKvxNHepa9l0quAfj+0lbMukxuHis8xhOkANOQA6TnufLPecIXISbFg0MkCJkReZdjTRSBw3Alp2
cjkBroqzykD9pxsYjU9Lb/D4JEUokucH3J02u1h1D9CZqtcyC2JJLzv1XIy75p8DiEgvfK800Gzj
M5vv+F2dVOBm/qLpn16JQusipGEbnOd4sMx/Cvyv+hRbOUA470CvznM3DpmVc90WeHwd17FXeX0Z
crtybArLTrtvsK2xakM19SqSc4OhCOyFgrTuc2YVOS3MYhyNQCoDjPPgFwLYIZYsWJ26/7S6XSCG
2xTdP/vUE31Yk9HAaQCFwcNDOETpsDnD1Yl0ZbBOdgB/CS1smV1I11stDxFRhFQ+AcWLrpFM4+UW
QeJ9X51pjuIAj+rWNtWcNmejsJDclryIB8uCHjUK3Jh+W667wTOssm2avnwg4vzarCmtHrvbZS31
+2Y+OXSV4E7897jLEgXMR83gW/MrcR2txlLJeefsusmuQ7DBY6yVTGgNerIoLVB4ENzulEXLwFrJ
J8MbeCNHMu4SXdo10vEinks/GRiXIdCg3yeDr8wL8j3/KSjkkjYlIU4AoYtGI7xVarcQnHsQe7NN
82GAK7dusIumwuEu4bSF5e0wXEP1EvudEGDgvdN2HGmsGNc9W0Fz0eW3eU8YXUsvW+nItzCNuTbL
+WXQnqi0KxhtiXujpyf8Aa4WDfqq8pYX5QGEe3cKuHHhtqPQHDVkFYX9DdclUzkTDY0THwOy/1um
TBIjMnV4lrbyP3f0Q7pOBWcBiYBGlmKsDncKfnKbfPntuNEzwjwhOjDFZ4ihfE8l5gQ4nhlPV8ZY
4aNAqBpYm5Fraa3g8XGeVJEF2J6ISZ9zMNbWHvCXnrFmsgkQ2/4msP2Q3scE/KxV4nldV/pQcr0Q
yIU04KAwjr5JqwAqamdDwXEftiYxQZQ7F5cD7Y7/J0l9whpIQslCGLRtgWpDhY6CGXXov3oIBY1U
Y/napBQM1khBw6Uodg4yEwT1h699SC5ENPsZLDJ6mJEak21M7coa4faWK/Sbfbv5PkIBVdUKgHJC
zWK95W3ax1wlJe+Lewy1mAxtOWc3J9fvlSj4qgruJ2d0wvvNd77d93QlXuzKpcmACT5BKUKrujeC
M9aKEGv8oYvIWibjw5Ks4VG/i4XEOnrTnYpBGRC9N0qRimJdACHXTwkRZ4X6+Pj63k2vjMbSrsVe
rtCXDrOnoKrotJjky/qYl8yVNgnCynnuBPIcYZYMXahO/3Q0gmaDxTytscCKwt9CqpCce4BHYLGP
pvan9UbrBQKU9XsbrFEds+LSlReJ5xE5g+LNi6yh+HBRRj20wdbc89MuXYkeeC/0uoJ3TkRhxG+2
JEoYFMQBSsvC5tnJeM7T+Eri5AdILXLRa0XU8EuCBNAQvPjbgGirsStwilGknZEKmb5Lo2T50R6F
abNIvFPw+GMkLuvUZD5EP+5wxTs43tGQh2V4D9QBkTJM46cxvsKXpiOJqiJXOY2f3xtOX9YBda03
jwvO/5C2dsWbf4dFBT5zDNoeUH087XwLBmwYk70WV7njcl0bAY6gy9R3yl+OAe6RPcvuHyDBaPu8
QnSwDn+rGJ+OMiiRUBsPRylY7jY6W2FACt9/YSXGSrkeiRHkbs6futpYqeDs3XqpqaX2MAxfeX3E
Onda2UMzQt9UpoJCBKb8tfamUHOk/g4XCqwq8zCkTXb5VW17NzAoWCOryBqDS4i0TgvoLWw9zLU4
LFz1zFUZCycbKJJTCeJk+KdSTARORcCBb/Xmi35nfOwNfuxq/Fe2Dd2jJYrWWbs5JYwrc2K1e1aR
s8mcHk7oFFrwNkWKmGoJYmwD4AdOkoN3ALoAQm6+6M88sAjT3qh30CEMXw3LVWvToD7dG6AV7zlX
G/1XHTGAxVUlYJ5dF3xxQVh2TY/l/sWmAdhAaCoi8BQDKEyNUF0tMSivoxeuPwvr3IfknqHYYEPb
IDsDMLFgz36hqdoPsYh7nOKIgR6vwfFyahxGVIGlwGgiF7Y0t0X+3SvJbU7Hy9MMY9TgGo3ivjtg
KUjjfcEbKDnJ1XfEi7DuwhbjVIJUMWtw8pBSTW25sHtbKySDuTjgb1JqGLKEOgukEUw7QS0xyowq
X8AOSx3nZDAtlK8ao9Ko5+3rSe2q0IGzzCtT/n5hPKX4VfMI21dHxCDfvugPQUA9fBXqWDayH4F3
atnK8dg16fenOrGpXcAsElrGaXMn7GgTIr3477ROHKQtW2LZYxAzbtVj8q6qPAFafAl6l4DzRHlL
G+yBJ43cMvy6Sy2CA5UWBgIp5YpLFT1Zff0QmtOMIyC6wINLbd51Dlthoj/mulvWOwcoCRca89Py
zWC22Uzrq+RX6ywYGXLOy3vH/O3Ns72H35jnZ81neNea+wIh6/0BWG/XTf3wjlJgHzZhoMfF0JyS
015czGfgBsBnAtn4tmz7yVbMadu55C28jbTQ4ZEzBqDNDG62tquU00HXcNFj1ITaVWUh1MScnyKS
S1puno1aAFZiKZ5OPKEXESdmM0nkWkDP1y/OpsfQ4lhmUVrkXvbOkv2xUUCH0gXrGYYYIIOw5r7m
9Mx4mHOsNhn50M8Z9UD30mGuC0Arlrd3XYwrRvn/d/QQPhvUxR1flzEr754mX41Ax7FDPjTH0oJz
6TAaa77AChkzVMsPTFHDhekeOgg+qYsMA1ro3u5DPREkhzvFq1MTyrXGVGwyQDQnAcZO/tGPF+bA
E/vHIQSoLrE8Ctb5fO7Vx6S1zrplFnDwnZ7TB6e+nple6GVVfj/IURLFs5MbtW7bPJ6tTDRXI1lM
6MD2KCSjOkk8psvjqLSs7cRvNhzH3EqYgxJ0YQBuK0mM47jgYz8l1ekvsqDNZ9LzS7Ih3GYEOC9p
KpWXAd3xIybXoW88C/SqqmBcsHfqR/SrTl/H6/paK+ZPPxE4Y0Lfn5gohFAqnnTHOvdTm1/oQGys
6T59Sg8IgBl7c+YY0VvyvMWVDnzYWwOTKblYHQgwUGdtGqtKXgNZxkgwd0DzesEQu7OMbipiypbq
a8dW9FxKAv5jQhsvNrde+0Zm5L3uTuF+3jbcKG/nn0c2JF0tHmXu8Y4R49meXcVHy78z5bqUXlF3
F2ImFAbu32XtTcUn5HfNCzjeqkXEX9MG2zqS/Xjic0t30zhcBPPJL+74p4dysqCfvqah+SF25F5v
lzvB2fuDzofdtz3OLqSB4GVRyC+MJC4Ed1pXGqQt4BQiF8DE0/AjYioGeniR2JS2RIiLnSpkzSAP
rElGNLiR23HmnafGk3e+UAE4nDRSqE5fWmK/BrwfwwF7IJv3AHYNSooomgeRtns2ndjXcxdQ2r3Q
dgj/c1JqYUudK9yN0/rZ9eYOktFXtVg+so8z/v4C+cMa55F2Uui+3OMN71lCEA/FxFG5KZNAEMq4
vdEcoujR2NC/zAsjl3RbvqV531GwOM2S05I3Kfl7poC3sD3e0KYLC8lmbT5ogn9DNpKgSgFqpxT7
sG3o8XaRfyCxPvp9+/x8xt6ZksYbHe8jfb7ov3LQxoPNEb2uGELG+6ClCOXHBu7b2pXa8NjX7mLz
FHXf6jvAr3PVDrTSMSsLn54ts8ypWuYsFLMU0JHZtO7TKmScXYijBjZgCqeG43HWlSjMDC50H5gL
ukXUKPXc0u83WMnO7GMjyyCACjKtqCg0UYwyg7yNcwV1pF4rLJ6ehfafnDf5yI9LkXrqsrJtaSkT
/10Vn2IXw5srOYbX4iaop7mCIHMxiYBeKmUnXBLBzhg06mPzettT+ZKqVfxZ9SYr+zYfoM/mPtYI
YvWsUAymmWANE20xFZ5vdo1SwJbddRv/BYFBwEU36LBuXDo6L1RNsF+p5YGwUvcB64Pil+KYX5E8
E1D+v/4IBn5ybbSQZJvn3v2nL6X/2YWTBKjUtL325hcfAH+zXnbu+DMOXI0EfoUWE1dk4UhpT+rN
rzmGIJg+VMo3k+Ah4Q4VLwtuxvUfGH0kEuulFYTQcJW6rkiiFofOunyvgR3tihYs9jHWEBMWnQtE
ONl3Ao2xNRIy6424tUjQAQEdE2N0QCxADb1g3NxHsESpz/n9UtBx6qwa/whrKhB4wpVqC+3Ekc/0
ZzPsP+qvYZjPPnVHjlpWnSDx+tDRrfNaAxdGlv4+GG5xbY8yhzorhBiwQOVTYnJ/nesK0SQdY1y2
Z3o/lkz/Y1jJBPRjwawZtC03VuBEotzIe8HPK/r3B4QhvJNqZXkUp3itlvfiSURagdivByR+BHvn
DbIkoz8MbK3MVBltQ5mdU6F+gWXZOug5S1MyQ7iEE6XAahmCQt/xG/SMCq3VdN8VlarisOyrR70h
7NKAo7r1UxVDbOQ1UBlySxB3GK3mVxqcD3XDqkXr+55YN7UFmLBMe5MuWeIUQMvfugKLjDouFFEy
1HrLW1SWdfRFrw52sP46hbfAiCHY29L9TXX2WW0McTseO/j0/FwP8Fkp0lfF5KDa5DRpR75JEvJm
wClMbrRjGmDcd6E6lTkzNAbVE9rauObqcRxZLcVxSl6zFS1z7mtDkFyfpvpZ1zInz0lY0b1O/O42
fnJ3tY2baxnEX4IyOmVpIdXSx1fX8lqsvC9pFGNerzcrsp5meeXCY3ldIrTWwN68HltZxPNaO9IU
ducNIXSmA+sipt2OU+txU7v3P7s1/uottzDzBrYbunEKdh70muqkdXs+m/FGOgyfxXgk1N6gWO6O
KFzoZ1QxrRGVihIw0//hYZSSYKlkJwh2Ml3cwPJ7XEyQDrHiFuv1N+7FEBD0UexmO9vW0E/5PrgU
TNzHEfToNMeQ/rZGoV62/jTe93It+qMon1P5tbJpsj20SFKpji/64wjKZ237za0038dFlq6Bh1WB
3bQfxp96CLpiDQEErwX+2qS5jszlABggp63Jzj7ih9O2fkktuSel5AIvE/YHT76GewOCHzb8qbI2
W2T6RDEby9kBGiM8/Rssdlq4XxRlL1TdrflHc9A59UDWSCzIYlUcwNUbCqemlEyViwK4BohV//hi
3KK4xAgsgHzMLe0x6PwA5YzJQ0rTJrcRVK9ZSNkfFF3PiV1rJ0kpr8wM+uCcDNl5rp1R6m8eYD0d
IamOU8g2uSriHGw7w0eL/FaWee2llZHJeV5c049spdBXpUe3yYOouxlhX1CTmmfRoVnF1cH7wjAr
mboQzTyDX+UusuyOSMfIb4Fl1zO4i5o0vZqyI8o+4z4WUIlZraSbXS3yEV0e1eOiFET7leJU+6SW
6NvHoo7DXgxIhyNjnqD89kyJG5YCJrYUK9ED+4wjt/m+GGeUJTRpP0g8u+oZS3iD0BUTDhJyQrwK
legJu8ovDsQquPqanmc39+bgpSSfkyBSQQBKy2D90xRjYy0mgnmcfZHt1rQttxp0nZz/nfcRSui+
zyYdg9PjAYswAUf4QJiJHCC0nVY5g5+kfeLrk4hcj9NlShQUfrKitnNtDEODkqhsfmOqePw0rCIT
4Iux2W7M7G9KLfprhwlrb4zfA8kY4JOp/Wq6uLMP4q3Dq6xWiBmqh0akf0U5Jurly28zjByuQfPI
uA5aaT7EWb2glEU728YFPSt+6h88XOpI4u8d68XENK0v/WEPuE2qijCtJd8TGUhav7UyadcWhv5R
k5e2FrbGvKzDUoBJgQ7D9r0OGiyBsl3/Bjpy65LM2UVSAgpNud4360LuhJM4waowDAcGBFfUjRXt
/RXt1K/e/t17V+s3DT0c2xLKQqI7M3cyF2ytZA2j0E+xcpHEGpR+igXVT5FRgrdMqU0/Dp06KX4h
zr1xR/mD+tG33okbQ83jwkUGLRB2Zv89tRItwwG8SfO/QxanQjIQOkoLM+rVNg4AoW8c0F/m9M68
IZLIpzU3QyoGjr9xSAE3ymLSxKlsfbQ2Vk/Qe43BHEjWPRyNczN0MuAQoDtyYJi7+wJ3EAo7xZzv
A+5yeuPW53Pp/H8MfX6dyHvTBTiLD4+RxZ1szr1BrArEALkl5tEV7/GqZPgjn4zCZw+O7dApOSuP
DJw2YoKlexr9t4cOpv0kJX6jhLk3vkuUnnN36UFD7OFdXHc71/KH8VVJSiQCHjJ9xyq48ixKvNg3
MFRWEoPco/3Q2l8vfj5/8GwokVZr9+UiGw1f70pIzSPk1Fg0fnToM8M/BsOYa+Ta5g7g/C9y3ebb
V69RJjho58x2yedIEciCylST6ozqRAhvcu8/X8J2dm/6Xp4Q8x0AyfAgrKx0m8ibnypVk4KFMyCv
vd0N4JvpnWaup0fIVAMkiVwcRc7/h8Bm1oDXosaGpUnGeZn9zhDu2xhq9Ut1PMFMMHoiCoCyg6p6
qFOJo/skVKgoGL1Rt6vUf00dQURc8l97vUnO6u8pUKtiq7J82g9L5/TK4DCpXyMO32+/R3Pt1FkA
516I/bsW33x/hhJF2o6Qs3ubWI9bNwygdPZ/oos43Oh9FsafgC3kJEp87brVgHRn9r8eo7vLxWzr
XemV91HgQ4B3fWdTm5IAwotLVEMcmVDbai5I4E50BF6NAvDs1fcZoRx9ve1fz+t7LxeL7LzqGlWM
pnlxPsXyu1ON/VPnRWdnVCjPcucKYnYFWErCRTKkblVVFG2H15JBdthirFfaiRI+8jAd3kRR4SlD
NMB1Rx9qIhHRh/uz2kzhjck06kMREIvGxwl9TAoHQk1IvdPUCRZM5mtXpMqcYisucGA5Ck//r1WT
jMzq8BHPj9GzYj5Yy7V7kZIo/QgindLrz+TDq3qsHmOnM6FDubtQInjaOq4I4SMtkWeTlClItPGi
J0c8bhLo8DCQ7CmsUwFptumZYiKbBK/2uv6ISRfK5RaCoQdAw7b35M6fgS3jRAx09hCDFpK6FmTe
0A8KNXpiMV2P+JVKlFjdnUQEu/f6TaBrvmbatZuvk3xbeCGAFH3CmQuzwlnAobMX54Hp7/DpptXU
DPvuS9LdpN1/4m+B4ctTCPa/2OCCpKEOeLMAX29E7tKMU+dePT0ECTOhYhWG+Q6RzYD/FvFHpD8a
iNvbB1PAo9mm7aWjXGEEwwjBlJnOWejui3LBmtVrbjTNzbrw0QWK2uyO8gEV8AgnrOdcqJ0dP9oS
cURv5PgvKSVbV+7NWKzTDqPSgrwjb3jgvzMANVHMoS5Agxco7pwIomiWQbh0XGBYflcTy4Pg0g5V
BAlUWbUysOZ/GCuWJmUiJ1Ku75EmnBeaK1N4msS/RlFITH8OQSUW8dM9F98rVZy3qfJhHL3bNxb2
D4oTHsa8XkUaAXbsd7EoiTX6govvB11/Fv12l95h3cyzfb+moT6CfOZcpGNokE2rIrkv3l8s5xsU
uvRzraXKJspe42FqV6hNuBt/yDfJc/EU+q6MMsv9i4mi/o8y79axjTkxsJ9P/OKr55mf+LYof9Kz
Zao/eDlvDXrLBzCjtOzXWjNy1om1FfoGaAxA2iVTgHyuuGs/DS0HAzipeHEfe7VSEoOBudQ3MFZc
CnMSbnCLXCoHHscRA1yFCO+AnggLPWQaBJ6L7NupmCWkDJvWHlhsE9FSUh5jJyLTmpsc2n5PnUb3
WTuxwtWN4avOezKBCAhZG/AqJAtVgIAW8mbI0oFIo7uopWZXXn3+yAfG0bAD2/2i4Ziu8Dw4fauu
UCoSdRbLJPiNXXny6ovIb/IJfvEKf/UQ3VFKfWz5vBJtgO9ltyegYHjavaqkZpTRAM3XgiE33RV+
HfgeEYON5saG2Cw5RFGFd8LzPZ+yu46TzYPkzc3XBqICSQ2UNmWZOa8DnNMhZX+uH7nFmSYD3yZQ
tM8bUQ+3A6t3T7oIEXgwvDexitxcDtTaHg4Tw8FiFnLXL7Y/dsNdx7fzmWxSzA5lEfI5DvUmEhIk
iyl/NAzU8/yZsYBj2jQCjDCn5pU9g0H3OOS98HIqNndCi38PM84aAAI/XTPkhwpzQiEcV5ou7pZi
RMm3WbwUE7IhOcls2ef7Y8w2+KK4ErzQJiOw71I0wPYtOq7FVC3+AMst85U53J8POTxq7mFPnvGY
001eMahlHzNwP50fNDSAv9yIj5qDk+VvQVibTbD7V+9YGG/nwgS7yUTGKrlAcG/g6by2Id+jYyn6
9OjcT+Jc6OMT20S4ZPkw5PULVRTwUxXDXISgrb1Qk0NJoehbEkRtzEYXm9m9ck+rsBRgxUiPOJqS
BXxZUXk8AW8u616uRffnQYOf/GN6zvYr+wRj9K/2I321/PcTThwwovrNOJhBJfdDyf4m9nz/ODA/
yKlMaP9T/P3Oqh3TwRGXy0hTMfmd4nuvyemCspmwd/9Janih5dG7cAgIqmu+AiNfLyiLCJmVwv8X
lgvGfCoL5Dtop7TIjvE31K92nmBJKu3hM1oY90TR9Gt6o+vFjSBruSNHD7qrtXFfzzZXNA5J1oot
J+gdHOA2HZ9+cYioyWQx/I/7V50mMu99FP3YH3MsmUjPRFxh/KBmWJrh8cwqJMz5BLrGOlnSB2e5
dZ/NHPvSZqBrs2gFTHVK4k8SXUBIZ6liHF2E++Wks4HFpcrIdQojq9IsR3ViOQ+HqXmsKQL6xWzo
ai7hI/nBPqEPY81o/MXhx/vWUvPhLRRqMJaoyDIZf4vhmV8XXB/nWjqpJEiBTlafTpCkzPsiq4m9
Fq6jkk9mgt9bW96vFxY74lazE/ONv7CzaUNAveih+xXVOGEdZswn+rHGmzuCUlBHfEd5QDVQqC7o
nKg0KqcJkD/Wg3YNbIWb0UHFcWEkjjE2YVujKIiEH50YYMHrIQ69lbhx5BPoDxu3RaP3Zpga62So
2NlBqokBxyE42tbpC2iQ1vpv1vZAM1Ifaod0dj9w6m4EXgy3kCx7BWu+5NWouLtZBhXY25fJKzpv
pzfGWgN8BFhjuPjcZVcjxUbeLESNEsQCln0m8NEo8TnttX4JX2t1zP3gsYqgPhs2l/CrYAWqf7Ft
Qzyq/mXYN8DMON8yjRlevnFn47fP3Yn5ndCHMB8n7XphMCJdBKqnKxvLaYr/YahjeD5jIb2QfiXe
chxo72oDrMRXy/j6+lKP9INM5W5Orl+dipg4Qsa0PegmzY+G4BNCRSYRCVSsIRaAq+mpEHnRxeEs
WNcqZXEPh8fjpyIaB0rlQMRmdoOxYk6NShRFSqWCay4RrSNX4qh/oS6PUYY3y2zqClN93uPr/llO
/gUsJvSlImUvvRlMRJMQG5H5x+oxKaPyH2jBu3CyRe08LGHEblevh+D3taCFMAnaPC+7PpYDvbZ+
TuZA84z4gO3tJXrLFZt7kJiWCc9rGP8hUwYioQH8QfnXE70fwBfK0u2OPVaPw+pB+47bTSjeO71i
aJcyrD3VNOW88nlefjBzTGnPO1hw4P3YFUX0KvWTa8qhBiuTJ6s6Wtm/fUNDxS/I1aB6lDP0lX7x
aIJyI60XV8NTMtFGcuB6h/5h7dO+W3BlsUahx5Ex5q1doiuRSaWhcfUm66W2lfW3HaZn7L2rwv0l
HchJxFgguAN7SBhuA3SETRqEoiIycumi+YwOBCGo8/BlK7eLp+pD8NFCXpLUPWMPVVyDQh80CnR6
iZzyDnrg6W30y9QIGr2aglgQ53NfxZFBRBhrB+ADMZwVpqgkfouqja6xEiiduU3sZw6WtHcH70BU
hI4WtEufgqPt6x4OP+mQNAHOpGVnPwAuJVz1EFvH5DXclQg/jue230J4UEWsR7v8QV9Fgu+1cCxc
MchpgXZ1XSOGuPAdvfbMM8oYNF4xIr5R5KnFzS4AqgUkRzZ3grxSwHaIEagAywn2aYyJyZm3GvOe
OpJqJzM+df0V0TOwX7au1LBHTrXP8ce3GCQOFb3rXLJf3SwjQ08fqaqLg3Xw27L3V3cUs19RBAhv
d+KG2YxRGyzuj0KAdgLl2inztfzXgW0zuXvyXaUdtGMzYM4Jj9KcKAcQRYLSLvmdN23Km82GPAaD
szjfy5v3j5VMLUjqq1bbJV+Ph3FphB9hEsISfVFede5S0Xpm2t0NFmHACOAtSUTiV40Mt9q1I7+5
5AQ6kt9AHoLzLkkAA507MrZvfB/cRKWkDOf3sdzGNb7Yz+FJFBi/Y6ugpFudP1AGO7WKVc7KBaUY
2P2SvgZbTfDWgXbc9suCrXPfUtXu/lDydPzQuRCd6SMGJcqtk8kC34csUE6fOmCgXjqxif+PSr4c
sbmtaOoowRVgPm9+0SekTOlH9/I6Ioas66uiDwHYiTNjYw2mgbl7LlVBVJ9Jwih7r1Nb2xkH+5uV
athjZNImq7rWFN+GPIt7V+Qx2Klahn4JPPuukpYw8hZrJYWRHE/ZXKGC3HorfFfni2JzwrD0ranr
5U5gihqKnh8kfPMgV0YOHBbR8wIscvvKzgtJuV9mseUDcgx31VUJRFlJpQK1SRFBFKghNoeAAcSw
rQ78rbiTIU67Li1a+eojQCCDoEuBFFvoTjas1S/vG3yewC4MoBacS50qSXHhsxBxtac5o6aBgXEk
xV0cdAv7RdFLv+RThWNLhzslfqghB8R4Udp4WxvjhXJMo4mEoLXaauKM8HTAXQBBneHPI+YKcK1i
NuVHJ1g6mNlV8ytp28/T5bXYuoMWHB+OgsW7R6KYiYx+9D6abzsEUiJh2LevOStXBnXVceGOnnmt
5gCLVCmfbSLKTvTuS1xo9kCVVCr90bi9WbyvSY/gGgnLFee1oP+zrEXBb2PGkpzqfQjRY5mu/vVE
7PwTmlrnx5gJM+BT7oBM2mMtlkIcoY4077l80bJkSzdRK9aD5YvyVkQ7iGYxbOGyg5rFWjdoyZes
Ijs303wp30bnYfiyjUiAqNdpovUicIs59kOpYhYXu00VlD+7dPAlS8VxJ7GY7JZzrIDqgDX7QSte
yND3YqhP83q5an+zCNB9VVLBAVB0LXODDYywf12WlBEKmNjm4ub8ZGeK2gYuS4Igwkve0bmDPmIE
YwxSTZmlxlZd4jmJD6pEkcI3KTmUYHsbDTwnXysRrDVRmuRSEg2bKl9g28hPiMJ1Qux3VCEd+HP6
zh5drxC+XU/0OdJLTpVKtuM9Br4mbv+fBOYZG25sm8lhvEIl/6b0zDMfN8v9YTj4d3UxNqUYOpif
lyr1lK4L1sl3Xc2iL7RNmITr1V7bldH1JvKkaQeT7U9HnfGTChvrTZNSqHhm9YczulMqHGW0m9JD
v/cQ4z8Ftro2inr48notCseAJ3yCHJgXgNTugFW7GvPBXQkAutejqfttB1BwfAbNaRSF5T22JMUM
Xj+MrKa6SmvomsVjwuOcaMvrpSAuMQ9choJ/OGqpq0FP2498fabMntq9U0ac5PL0wNw5e9KRyfpB
Ei3kYpx3j3CaXT5K1/LqphmAyBA/siPQ4SBzFwGeW7cxPAE8TyamGs5nj3oCtaX/YdppGv3kpzwc
yVjbgEZeVnD3qIuvdJ6subBX2CZh6CXoqNBLo5YMK1r8ZbgfzyM2qdmWx6Ah7jOFpg6vwpMhQqk9
++trvkR1ffmEucqBY1ps95y/UNdSNZbn3LafvNmZ+tuQpnwBtYVa/bETXkeN0npNhWVO/FMC/1cq
2jQqZuk6oEteOD3Nbdhcvx/Nl7mqZcJt4TAUPYW10fgxSPBldoDHTszOqqD7I5J6hontE5UI8LL0
xEApQ8CVeRwlIKDOLKeKVnjlvsL7Ecnrqqbs6r65m4y5enzPs5+Yy8N6aV8erbcqtUAZE5lndT/h
a5GAUaZprloiDMVBmyUfybsjgBZ8cLehZ4QJ3p+ypcpR3lgs859HGjQtPyDlLVnWxTuigBEj0bn5
xlkRUTv2Bn5rQIDq6Nd9ORUXUOM/mpr57oKSFLr05daO0i15gG8UgfrK7yfSIJJrJx3VAe86/clv
NSsjABlwBbaL61m3pntgyrKSXnQTIwCsW2HJBQc7kWYFkI8s2fAuZARhKBn4MRMteHvuIesqCnsv
+/3WbjVdISRo+eZ+5XR82CWp6YXbfz6TpeoynV//97Dhgd0/LtXTFfSoG2L/yOVAA47KZhbMse9G
Tk/Wrm8PqLsUu4DsvvQna28572j1XUN4NSnLtOsapXebvUA6lB94o1wFFy6UhwbdyAjEmZhDJex7
CpPA2H8ZyfiLwo/v2U5DTQf5kbP3rUTmivOeZ6CIaaYfa2dz+9d3U6P/RR3hprui5BWSWfNz7O7/
H/0xL6AS7BpZ7nwnWWzoP1MGd1RZHeb1WgksqL3kJd+ZxpSYixNZg+oT4ZeMjb+25hls0h8v6n2B
qX3+XSNVw4Yg9K0dVVkVlDhkOo4mQku6Wpsfsy5De+oBJFXnn6znRLTe9gn9x+MnJg+sxjPNXO8c
1NUn8wXS3RMklXwacn3vAg1Z82WQfvTC8YZ/M3olDo3LHpP6A+FmdGTgx0+iwBlKyPOWB8EsKXYs
BSQJ1+E++0NiL8fRmyyQCRL9xXWfI1cyW6dFdbkcfTuoeeEMsOhkgSmwFfA8vcHx9yRbbvXkaT/s
bOkYzM5h05czjKuPjAiXYouVPmb8atDOvmua9tQwP4id0EoTg36Ex/p/VgE3PxZ3S4wfrpUTAeCd
Vlt8H5vZ8Zza9L4KaRDwKg+z0nNoEH9Vrfohe8Cko16Ed75EuyTJLx0pdDBbDgNVfa5EoUCaPybv
ziVSBc/0yxRelXd7qEyAdwraT2dqnc9SLvqAfSvOlyzhCPYpXk5IAXzWDcGBAycrMscVh+GA62ST
R2kN9ljing6Tf/mXwis+1tGTjr81xb1+KBE0+u+dOxl8DAjiGbUCBllBlI2t38Oxie4CDpw5vkIC
qBXQsPRfATUViaMza4vrLvY3wSiU/kyQlsMvbgVJUQ5RVqIoX7/Diwe0W2urC1sycEV3WKlSwURJ
LLgb4oYJWmc00r0WaOTrshwWtKIwrIDml1nTKfgiXaYjeBcRHcDq1pwXYl+A0p3r00wxT+G4vckH
6lyahOkyZl+pggeVO090szizi56RjUDj/xoereCKc38yXt0BG0T9CydcIeqNTlZmqI8b7NdKRq0+
lh+mno4GdOoSHXriMetBAluakhrHjfCYv0anyCoTq8O8crD7oFkj/YZ4Z8cPE0EFPnmEx5sea+ey
GKut56WDruAqIJHETECIZ8xYbG0xg9947YFXiu/DfXXKYLffzk39TH2bD/Q1VbsHahX9kj9w9lHQ
RX0S32fC/oKXTppV9eQ9CERiwOW1V2pvXOvZB+Uf1tJFbNyA5ysrayRFFF6e16aYkRWwb0HW8oYP
XLNADwyIpGNBbYbukEn8M2/iRhKCtK63imx4wZlAUHtrrTKatZhYjzbOYi9xNr/IdTE9sijy0ho6
WkYUrg0I0E4AZz/I9HRuu7a2Q5u/5XOs/RDLrmlseSVAG6l9CrmAdRhaa+/cp6jXcGKx+/mjHskV
zuSZW+r5pmxDOIGBg3WeHLMCmCEhOgrAKuF6fuwRi1MOBD7e1NshTCaNARjs5+bKqw7qQy+NCJZK
jJdQjrmks5Sc7tXmU4p3ICV+3uG+3Bw5a/XQWyRqpsW/5elZVv61ZKDn31WpTNLRI7muBXpeSFoH
qbyup4d1dmJT2nZCbZX/VBtBJ5t/4hmHUYU13xGRNErleXhboGtaJvqX44ZaPbHUk2Dn4N/jgORp
eTlgr/P6dg5StFgVZb/WGsDVLdHUGv+F1lfo4PcULVOjzVUCi61uM3rooGJukYNjo4oH2MtwQg9Z
SbbZehERUyhq+leStVz/miyJSSTK8MhxP0HhDp9jCzRam8Cb/lNvgp0MTyYJxkMpxJTyZxLtGcxL
nYPH3ScXPEHD5rZd4sYU+8mIIcAtYGNofyndwgAXAxSo+dyPSlpVY1M9UgDhuUqaqs6z1VfyxbYY
kc3fLUY0C14fNuvSO5l0aUjdYBF4lN3TlZPlx327kmyBwZ48TITisuVzSuXkLrXYEf0qo69bu7Xr
lwSxO6hompudeo6ikZglol0iHc/V6omAoahynB/6YcFh9LbIlJ7IF9ndzaknjkzznS0DlqQAp1k6
6KfS42x29g8JPNfV0xStpNkv36++KbvuE6qzmeBF1tBv9GCnweDk76klGfh0BHKK5TzqwKqxmgqo
zQMI7fLQhUMMAQfJwieBw24OkZZ9WoXHsisFvnI+6QWDgxDThJ8kmOMFcXdEMde3WnepyVPk4Xyj
fPV8Qh1fyVSarq5Td5kEyOZQPrM5sIVXlLGVjmQo2HKEWSrIjQvOGSC+JJuTqootbYU+5PhPw70r
peSzOjJCySGyySYFf509kd2/UZSsZNTOhoA3Ne6YFHyckqslOCQOt91eEhE2eX5iWg5czi4XvKHS
bKoxdMDZUS/PGgwFehitQvN7KawE+Lxuj5sH+N9A3ftlt5tzxdLUrh3iK+U1QLHcbrWPHEHovWet
2VFNkmVLtAPxG8ZqLFwRQdvBIvnMKJXyezZFJX1tkQDn7r/jGZN5fXi8m9I+5rdq1i1XojmMmlyZ
qccGpEuUcqJMMJX5YFtV64NAgShM6zq4SoYCXN3v9IS20etrbpQVd6IZMUesPkNPSZCP0oeHdORb
I8BTsjT41cbhMezekwVo+TPIQlc/Go10zlbQD+VKY+5WVeJzR2tt25brVangZ0yXn7kegYFDyLJJ
YiyloysPqQOvTfM6xus9E1CXxv7DvcxF4h66OVWJugmtIGEA/QszpE85jNUzTpF3xnpW9dgjkcML
9fium+iC2POSN6QrhcpXfpzcAR9b0GnDTApJ25+bVBzbwPwq1lHFs4AgHJftq3vKkZBez5mbNt1K
5USO0DmvExGIxmEQxQV1a10KEkBLPm4WqBtbvWR9o6F2wckmM55t/QDxVAVNZTARDstHqBb7S8wb
aim8qsjBLouIjZVDD+9srLgb26k/BhW7vn9VjSCLzYKK5hN5ba7V/aoebDABWiyFSmX+1pFxpcWC
KuGagqo1EUBRNhcnkbFHgatAzRAYdnkZafacT2ywkGAVQvJ5W95yEYFfsSIWATHY8whjyoTx4nVA
rcCLS0tjbDrKkvY6HEPmOPwezPSN9j6wPsOhP+wQgWJbHbb2gE6V1kXUBCSLIXdgkjUZOXK+a3jo
+jHbIZqHweFPROQlUdHWLX3XY3EAYgRToXvVt2fmgWhW7owx45A7TUhJfVrwJlA4DHVp4UXdAALq
SJYbAjRVHcJFXT3TACfI0WzZMogbmVXJQ91w013J61JhbPLce0MPiKZYMOB8BTT9lHohTMCODxcV
EPwSziQ2m03y7JN14Lc4Tz2Bu5wNaLK4TX4+CVjS8hzvY11GF/LoiW78A2m7bKl3yNgcGzy4tXRS
X1KhIZWtrPD4uztzhmIoiVMLTUQl8mtJ1hCEcwiaC4ISucbFHOhxclJvTMSXIjeWc14D1+Vct/q6
gDMFW9w6Z82m41Tqzkn78s7n9Pe83vFZnULAiVb/kelVNoQsaL1O0HMXzMAcYPhYnPdVfkhZim6R
IkfZVvI8m3b794EUrETaT3/5M5DPtnrNxZKKqnme3vi4mimyW9Oc0fRS3dGfZ01KjDgnsNcmcXx2
IKk0tDamcO3lVrKdVDlswEzyaBy4RgY2qCYOQ2spcCR+BYEoZiYAXHSV8Nfd75xQwST+jvf04B8q
6wvp1uzXUbbYLO1UcE9dCBOKmlcV5aUr5KnsZVY1rRFGezJwJ8eTP332qI8O16sRg1BSdwvoH3FD
5dLNOSBny9SSEMcnkE5o6uns4xuXNr/XXDGo3LqYSVP8t1gbNg79o4tg3Cv8b/c74VuksjklMSeZ
BggFjTxEpTJLgO3vcCiUOmGH8V+d3hqE4XBWpl3LCjDJWRX6wZnP4+oPFurACQi3ZumGPtKyA3LE
O5inx19ShYaEGSv1eHDTiIvAJ2V2lxRDujueuiJD/WXiS5GWlW+BciLbLvTblP2xEIiG0HqoIbt1
i2B1PG1WikDeoS11FPXcCx5jqySbsOJWWb9G4IN6OmiSkZ1rfGfV+VZd9kU9QUQu5yC9X3Vu4VQc
uqsJFBZt2q5TSsNXRzbvrUGvVMgxfhBRaO6/C3U1O4+g8HeXFsS89zMozFdEidc9kUaUPgD+8ic6
qJUsOiEstBjIlMXzuOqFXgMTNdjyKUyA8Q2ZY+K/5hNsk1Y3qQd+Wjo7y1fqeOaWB7k7RSLc+UUq
GBT2VN+uGeP/JYcRzHgqRi4ZI/jNMaxF1VJPBK86p5sbn0e1yXo7fuCzX/ydawWor49J3brr+uyI
ov/xnRqmyh83Ev8r8rgmEX4NGj/AVyVizAYGOJ3mARMeBbamDDMwi2mnPBty+I0BQQSVsXpPs3Tv
jSeum105MNLOaS5sXn1bH11n+4JxY89N9tQoBvu+3XwgiV5Qch/5VkBY5lmDcMKyPmAXgJQoMUkK
GUw5Uy8tPKAORG+cdL1BBa983qXBTJHvh1EGlo+CSbCWiuLxG8wEFr6gLpJpULB5zetTVXwTYlyg
SU2h7wHWd3xBXbL03/q2dz1wX/cQrLdqsf/EmdQuvWkqk47QzSZpMDuoFuYbDAwZOjUUrVjSe5aO
bGsE2DWIJyzGzbZAc+FK+kaMgvvs2bTHB/bd3TgZJgYbU9kyPNoxNitXhAXJ7LHf2YF+NqhtfZQZ
At0mfiSLAAbBH5NKp/GVafKu6vT6qROtb/rQ2lLi2GfQotL4+ksISfCdqhShcYuofGjZE1h39mY2
/fswGg5eloMGTHYYGQ2Sl8HIfb53Ew5SzXM2mAultzFVWeJH6jwO0cFGWJ+HhgFbLI8OEtAbJNWY
Wv+DIpYXCgckwT3A0l8OHwKjP8fOGXrwhWrIDoF3C2ZDToo8vpk5QdRYCd7D6D6KLJOLGvY5gQII
sVwGbHhDXbi/WPAUF2/55zhlIGqbPDYzeB+5dHT8XP00TlX8U4RkzfnuVHhPlOKJNPw7gAv6aOj+
GIL7aDXsWGyw+eBjMFkttuq0iP1OYLlM45QzfbbrkYro9pxDAGPO8FIdUUXC5Lv4YK/Wad0APX/U
giroyWyZZkRHrYSb9v9BfrbqCZ+9ps3YZBWPpIKyB5CwBryOqkS8AYD8TdkLKJuIBLSK/Fw4lbMM
gOqHNAcKPVKhvfsqciyvRHOfLBEciyMYv8pcKrDkUMXUJKby7AOgoH12GJduMOKb6vME55bsKxja
OUkDzRimDXBFBXXET/jGoKFybSfbv7ekxYvmu0erZDiR0JV7J1619qvESJucYZDJZxrKDiGMaqF8
sMNWpthXAdgihL0hDxOeZ5uPsDUa6SYjzJekOR7YElZxlb69h/bgVZnFqw45216XpX0xp+sXA1BH
z2ecVr4pKQyVJlcE+CK3chsPrCnf/QYYG+2+SxNBcJ5CoXVNX88PS0i57gDJfdbRI8Irc2lurtbJ
GaNpjCUnNTnRpReJXSVXwE3Jpu4hkarmWvbo/1Sr7T4ovSpdKhFkm5NuP8EOcZdA0NleKe82bsgY
rnEjPGSq53t+jAqSzeDBPs222QJAmJLnjZGAB40M38Y6VtpXx+Ocxtp8gt5BZtkSkUK++nslbU+A
r+zCSuZ0fj4dUbv54CJelynoac8srbict+Rvjm4W0GIhz+bzBbmWzfhHKo4/Y6AEFo1cY+Un39MG
ruHgtfnMwgOQjeOpffMk9GM/VfToC3Nt0ZRofWyCaNMvVIWpsTdjDk5TcNri9FxE1q7osnMxXG3m
Io2n1dhDI7aVRSjfLev0iV2q/sG1R+67HaeYfCqvmhf7F4DwwFhYEQul1Alolite3KeP3Bn3RyM+
ADUSSoPntuPgvvob+ObgG1u9DiNBk5U7hrneCjyc5Udx75KoiX6cGIOHaYMsXxNI699xJC3+Ddar
UHWILFTG/GcNHnSrjN0Xt6LrxIM784+h5T4wi7AU+ycz5hsPHWsFi1M8ku38V2okcpQTgo0BkwTZ
+yzE8aYP72TNd5U+nmt2pOTW1EzZxTfFJmJHQKH2269sOW2ZrOD+NDIGSZHcIM3NYt+qWrMPIEkd
+4vnKZD81thSS30LhkPW531lMWWhrH8K0tb7OzW1Aa4REf5mPo3mPD+dlz4v1T61dU6tOa+42Es2
8C58xKddm94MoVLCFOVel0UKYeEpWCGPbEk2kM8Q2pP63GAjGKbWEhrKkiN8rp0dH/A2wwmYq2vf
K5gMqtV0PJU6uW5dGTsq+pBF76giOcFKEZG9khiEu3rnFs29FqHH1Pgow5NfoZmqRRvgDmX0uYbS
RPR6UuBfuNZziZCqqJM/te+l3bFvQddRc7hij0WCQybU0Atdjt7eG2anxcfnf5OotbsUnvMVLpf5
LJGU9Yy3c1HNmDyandq5SdXTRm5f+dSwehm1y3goKRYiKwnGxeD9E86y6vDZu3MlrSKIWM5xcZCv
WU9y4XAAPZXi9eGoLJiZM/UgYJ9QwftibPmkp1vFIziOI0MyEHp3nw4Y04GTScYv1nGv/XV2Y2sb
HU0GNZ3mWyrsHrzG2/RpEK04/Ogx/bvDsG5VA9zwXjt1j64cIybVgCGpiVJ1dAXTinDdWJJQAMjP
ZjOe94VLOI33Ato/S8pvdK2eeyaRobrqwJmW1MTeqgWuKR4CAVLUk5IUKsbkx53hNKtHqiYuGpnG
n1ieIV1lZIOAoMW90hXV6CaENk2vltgLqLJJbhJWCucbvbTZw5G5YIcdB+NHHV/VnAx3llLZRmrY
cTn92XW7mUBIh/32t1EBcaw9cjYAbsHBFkR/jbwbNNxi4liuy+or1tgpjc7SBriOHF90rBOfgl8j
4Xk9TzHdosLRuD1oi0cz6FPlJKcYoW+szFQQq+2zc4V+FBhunTDf+xrHmZ1SYvx9Y3BPgL1lcXiQ
eBsQq9zD94FDzh2eX8IiaVplwvHZyjn/Yosy1dOJ71VK4wZcaG9PaMbvnKgEKR8bYJ5Tesh+V9uV
fmEjorM3Yb/WR61s6pJlhhMrYvMfZCDk1UwHpW+b1AZ1Birj8wr1kECUwkzbIZxklqZ2LruYnHfh
Ac8m5XVBby6hOvIgtHbcFgnVozdmFQxUTgzVYiZzc+98Cs+KhwZoR+abBKzDhloyjRAPRPZZr8ZW
1Ubc/RKb16mGwrFuk7tPfhXmdwZqTuiZV5rfiqKNVaWc2/j33c83EOxZgDFxUF6tjO3JF574hf0T
VyYdtyl1MUQD7MH7ytKH1S3Pbe3lUJMi5xOo/nF2HgtvWjGIwDrcwFsb0VS3ZFRyyJLogCyVhKf5
yNWfirqMBnU0qjTHtkStNiSShoRg0P44gZlk4ybXtGFM0Ag13GGKhsVxFPLdgjIBBbdafI7GLcnh
IQFyKT4NPrzdN6yfNDe2HsIPEKjDgSGm6rVDZD44K85xE/ZeJSo269p+bbMd90fIVLO/pSNiCii1
+F0hMhLqXuKI0bFOh8tbtz2oreoLoJ12SXusBysSxdkU/eUMAmt/YePgp5ehyVzRKq4kMNIxqHV/
NSBX8pP8DapZ/vHgCIjnjHXwUU1yNo28lePtSD6mBRamRsdoV81BQTFL3c6QPSu9MuIKN720Xa+m
RofNFMfUOkigrqdchQN5doHe3hmOK7ohLD83rf60K0XvexHi1cOOskNPabh5tVGIRPCsj2298PqV
Ev9zm3m9yB7kxfxxwDQ37hCubZyvFvauyE3uXaPI9oL+3BXAU771/IioVo+tya8wzuxtr/iBif2D
gY+MWUvAfgPrL4b3xY5mRQwlBuVKYdHd6GvYfxVSja906BqnU6hKbnhcVUcoLLiPHQn8NShivRm6
JMR17iapBFNYdxUJIEiV6y6L0QdJLnqUUlPK7gRbFwvKJWaarLf5dyFm8gIwC4ChGeW3Htkrxz4T
QMzJUXp/BP6JUo0LV8D8TgTdkLz8/+4dokqlL1A7iS4AU0BwpahIa9+dERobJfFMPN+GnPeNGnGN
bJuaFHZCvUudwpt4nyZBD493MpWTiPdOmEj5EjZCpC4D744E4FmqqvRnjPH0uIQH/Ydls968+bNr
L+29Lql8S8V4/jY1tD6wzLDjrBgdSbuDQLfUARxZOQzsYR5YhZHfvGKjfF1WdAWuzbSrs4Ufu4Fu
cCObZWBYFEfrGrHmHVko54QtOYvU5eaBmLIzGyxPqJeVOTVfGdPXD+9fIcWUg+pt5ns8U5THb4Bh
R49SwGrkTf3FzPf3u1nuFG7BaTU6Vmo2iFFkT4bvCpIwdTx6U748tnP5Ct9rSbWQZZKER5BqXCho
WbEc8QUUsZih4DxqxIidG58h9yW8sHdo3YEdguiUxT/MhwscXqV5f0MQ72Nwty4u+3LCV+aV/1ih
1fsTrHTcQRG7hbq2GtgTxCYGGovZZ9o2nQaYKyBVx2r884Z3BWWIeaWvJPKcmnwolpjpHjC1RtKP
P0XBAmBtQofUJxqDcZWkZA+cpbQnIigd2v4ERavV98/6Z6zsJ1AshzoNw+Ueuu4lrNeei5Wm4nXu
bFEzw5Dsq0uR80o7t+/gPDxeIC3MYs5Ca/W5QOosvRuowb0S4xcjzgi+Z2pr3RsKEy4p7qls7Vlf
6yhzLF93V0zfEyjIjSSZ9GBbK7qDyxGjUmTVqq0EfHM+xXR5UTdXpmY04zDe5XrY1uLXHKHDSpzz
83iBVt6HgpLPWJtU2y1QA0SeAL+FkgkahINJZtXmtqgmCDXUSw1P6vzw5mvULZm3qnqbFOUg+VPD
lH/KbQNP4k7JjaQZ+CFAAWsbpw+owwHFIOf6EG1YVJKfxUBkjh0m+jCCwyboaLXu3vBCQpPjMua2
SHhfkxose5bTcFN23fj6c5t7ly3+bXsaAVn0U2DYY33rhE/jGePFPOH/4wylV2C9pvif1oVxI6PG
5/NZgKwkwyTSUrAExsaYRjrM5kRMZ6XEAFYEMGY7RP9DiOLiMfGSgRUx6MBJMD9c6xDGZu+tpwHW
8AW+OZh1VIFE5hqpYIe5clDTjAu3R8P828SAw0jq1E0b5bRsde1olBP3MpC7NeKQhvB5t5M0vYjs
F05kowe4Yn6UzAsbmEDaJPuV7r7sUgHRPJVh2SMduxvZ/+Ps5UEYdxPRx9tpmKO//ZA4M9UVafYf
U3TZHPx4F44KJjhgQtJJrxlcF5VoomBLv5jbEpivnYeIDyEUR6LURxX1bRG63Gqx1sJEFS5ECSfP
iYrfRbr1OJ2WKwavawPgePAHK8x9mnXrNjpyHS387Ft6UjNE3p4whFVuvrYc1YicfmjfPbZlbf/C
hFA2h4T0faphdAGd4Vfg0KOlPgRGiYc2g6QUWv9py7T4moVGRvyvpeFpvQrOXDelIEQMV1Xbh9q2
9WQSzJn9QakkuJnXCkhfP2UVVLEZOFvi4yna9BMDF6u+clZ5k07tE2uI/uTHAdzOHBeDYupg5ZsS
sCA7vJaQ/E0VMc3R7p18A2BnV/BqPB7+x6ykX4CsGcDRhynmGR9gQ4oautLT6pgqnbts+AsheX6r
5aW4SWM2gBdbOHPYHYvWpZFqYSv7B3OXCzXfsSfGEFhwU7Wd2su07aC6w3Ml7IkJ5y3lPsxSdYyf
ftVMWZAx1YhAKG6qdOgbEsS5gmda1iY8Gqn5E9Q2ISybREFQyLz2DhuEJhmEsd3m/GKP0FZ5EdBr
I5/ciQiQiU7FXvfFqPpesls6lEdfpiI9hzHou1jz6/GnCX0BkeW13E9tWghNOwEC0UvlJ6ny3nJG
ySj+1GJkPgQduFWcXBxJmQLciec4AHlN23w6ns0eN32zQaowUitWMmp8ASVT4AA8OYo5osNb5Wya
+48uNlZHh86YcXdjiE4D1gyQ0LUTEXmNUEMkfwdHvdLI52iu0HZicF2HcbToq2uj5J7WKJwUheEo
J+7XvOG4242nuSr+ryZC5HbjfESbx2Zb2kVrjTMmHZ5fac7wUwg1N6RHTfVCIJzcwuamc/GQyx+A
E39PslylJLH3SEatqK2F4icG/zrvNYaWns0PIzon92PP/HIP9z9X6a/A8AVr4HnFm1qEloucIoJA
4rmgWXiFc4/IoXLG1tMzFUf7rGND1yJI0cc5W0kAIXdGf3Q7odx59LtKtvgEBPcnjy0wQP6K+hFW
xCcuvEG7t7qdb0Q1qyFPGVhm6u/8scQB54SBvNeDsEIcIhuOs4U9aUb3F/CS1rj62cU/gl/IqvuT
GUudGoOEtN6mCZryZR5uz6Uhci/mTkwuuj5grd5y4jykexQFG+SlL1YVI0+hJmwU2NHdlbPrVGsd
6C+OIDo7rrs3URim+xVBeMOglAv1s/2CtP7EOpos4OxeUbECgIqhKRTvbYfD7sK61JzI4JDqz6ds
2e1oAv0jYJ0PeCgGNk5PBT4EG0etQzrHpx8wVweVBCocrD72vi/l7F0mxYWkOqShaiZLFMD5r7eT
ZctP3bILqXPOkp+/iSfnskgI7iDf/XJiBRkr6y1QcNtJb27r/on/t+Xd1J4gcKoxO4gzEJAk3zTU
laJ3UZ7nNGPBLEztICBxKOa2yT4cOfWDcIidy+3m0savlaDKg+eURUt9FC5d+QL42RzTZ5K/TisX
/9i0z1JS5v0ZXSZwKx5ZJUeWeLZe88hW6AdkUHixCHZdN60bs6bOEt038+qMqvGkQir2p7ZquU9T
8/DQULhDchaOp49k4DOjeHyaZ5OP+2tOEN/3lXIcTBIMdXmriKOaq2cgjQdxTqSwMugKqmqe3xA1
d5841g9KDXoZ+GbZlDYWcFSFCrEW+C8Rme0BqeO3tQyITphgYP/VVpQIwgIPM21pytzgrbuLRvU1
R+Vu19auYVi0j14JnHGtb+u9FD6eSLWxtmNqPVU2jaDqUODrHgN+1q5imLutI6XjAN6Hbvh7yRMH
/gmgCiedg4lqvpNO2cCVAiVszCjwnlPE+mIHZSHp2JvmSvYnrvIukjbF6hXcpyQDwRjO8uAdS+vL
ynghX30Sh2HlUDs8bnoNPYRDDwxgRTWgiQA/5eWVAq1pUMydehJ1Q2/dkMmQ6ysEfbC5t5cLtcaZ
HNykFnwHtchPfm+ksjIyRQDSi4bt4FtSkyMdVTYbi8i3BS6fSlvnQP3Fl6n/KLv06HPNa2kVhiI4
P/GWmZlTEMKJ1c6CwGvkZcv+big81YNXKcM69GxcY4lQrOaZ0aCnjQWPu757NV78FoBep/5K+37B
MfVqimDoKf+O+tuP8FiYVCo+/vGmdvzQ+n63uC96XxbQaAHz2M0ax+M7nKIqCTRbqbxxf1tx0Fbv
h8IDLSHkXQYvDq4GA+xwuOfndn9FzWCsyOf7kmRVBl0pddPccSzxm3ZJKOrK6974qqhEksZz/xGr
4fgvR8kCApSuqI7x7MYOi1wqOEFuIQkCSQqA9CB2TcOaeEU1gVYv0HVJ4Bz/0A9/Z2CFtLktK9MU
VEosaCiqx/Vy+ycUgC5YthswCnTcFEh8LvaTZFrVEdv1IeuDi3pnodpw3oQgZuM/BtrX33W1yoeV
pXa0igjOQLaYroQ+0DzkCttxBu9E6fRLBT1U6g9Yss3OcBa7tCnOjqwks+fEHVasuG0sJkZOvVTc
wxjrnh8Cnw0kXkDmSqURQMGmtvOuFUmvuLb7WymPtTe1DAV8RWPFA9Ty5tqOt3Fpy7p6aRPpDfHK
5ZS/pfYQa56vdylOMYVNqkkla9FNEWafaX7KrO+AoYxtK0sepJTKWecAl+zvO0I+jTKlUdtmklxw
hOwLnHS9U9xqRD6x3VfBKFgZuNpBBnxqGLE0OSZ2Y6UIkhZN3PIEXGoDJOZaLIgRPbT9r7poBYX8
kGC3J69LkGp6T4EwMqYlQ32r5gRIrKjvwJ9qUvFR/kAMkBjqJYeJLwsZENV3J9kr40o8564WyOyP
dyYqqV+3NmA1d4wXe+0dA7pidh1/0pkGA1YWalYTXFamAwuVGnseuvd7ceUpJ3YfVoW+9F6MCvQN
8vMvobhYGsXrFti2ej70GKCEtm5swTiT6tsKOU+4d3514aiqqxkte63SO7AN6awlkSsHQdhvtANe
idf0RaHZ861rwmHisqqzpwpni5LnZfPZIvZILIPs9cuTjT22uBT89RQl4jVLYcZJYWAgKWsRbVIi
hgBOdgogVEKuwv8kE1dSlLm2uOtS16xrs7VAHNtD4Y/SiurPC1UfN4HfI4MYBdTC7Vb+lmGw0B9J
BALPfINH3u1tAn+8X6+DTTuXxrzRYjjb7Tspc+BLOaWO56x/M8ip9dKA+Ou/RNzedpAzdhx2Y610
ft6vdfMGqSZT/PkYXJt701KdKLJriBRdReGcVlSiFIWEwk1ehqHLPy/s3xKY9pvg4veeFA0AfEbB
8IASSl6CvqZuU5JBrF4X7Zo25mpg9XXPb2eHmKLBJbWeFWBYpTPXIKP5CtdIO0zg5F07IbNK5J+d
70GrU35vsNHrHUD5vLApxdUC55vIc1EQC/QQXrA3E2qJ0v39DzIjO0AIn3kfTDB5oIowLAN1EAxq
LeiSgu7dwJpMwMNS/naVhzqBfGwNuUFtwtKW8FgdHDoOiANfbUqJ+dIAFtJ9qyaM3Dp/m/yPKMgU
pmbs6r7NqlArBwMyrM5/84EpMPg9yu/i5fhRZZigQoVDZjboltjiD3TTf/LSLhQKswsGLhdZG7NL
IgqlkuhJKsUksZeJjV97Pgi1zsqe5CPUyikbdaBSH4sAqGDouNeADmkw1UkXpOX2uDhljSPR438Y
Yen/YNBkjPkKN+qAOpdFN5ngSQt1LwiBVn2+FRuQ12bTQJ3HTH0I9J+nysrfdqthUwmHkGlTfvXX
pgmKVe0KfWYLDW1W+GIxLn+srYzQqG97QKQb/XsRLE/yw2wvhxKL2M32XHk4250UiNj7p92XYIjU
C9cUj02nGqL7sZdsw9OVpuVEM8Uy9KlEs/qBh8hI0ZhsAiT7S7jlPkmI6AptVGMDNhHYnqJ3BWCg
uJvOotS3pQHMq+IgmJKRLTkaEeDkEq6Z1HXw0K25aVCu+1KyPSMObnyOu+C+PMAautKrZQpkopr2
dJCIR+LBsjF74nrTau7Yt7dLC0mkHfewuHUhvKF58YvtAv9zaC1aVKXzlYyV+v+cFdHZjVQVXSMZ
y6s/5dy9MfkQu8fZaCP0cJXnDQX/caym/33Sx+KhX1Fo/fpDs0JKBrkjHhJytxfxOjL2bG44Uyr+
qCuPHoS/9OE6XzPPLacnVq9Vk/FBDqDEGNZW3goNuVE7X4EWu2FceiB7n0Vy2PjSOIWU6yIMLETN
PNbEiPEhFef+bitGIVz2Rj4Satg+51jGSTCHroHNjXm8DIqRqGblgpT38TiPFGWyNnAMB8w26E2u
bHuj3ljgAj3eGSxZzPlXAxeZMBs+NOk7R7+FZuKCKGXW30hFapJV9RUnqAIn08QmZRMfGyGVYLjm
/SETynx1/niMitvgJHdbiqHHI/c09gQl+0b76GiW3/W9rq2uZW0l0ds2Tk9t0p7TAj6uPwjtaupP
Su8XhsEzhI4ivhooiJ6bY1vi2cm4eyU+Ws2SI1nOIFoZyQaNICt7HtCIxSs5M3XdHN/g8LVip9vP
IQbImmy5xisDqU/Q1NzruirFw3N7wQaOzKlgmCXoNLO+eLpI345xqYY6jgwZ4JsXq2vm9+ffBscW
+VC2F3exF6l2o8pm44LarR/Y8oUXmaVzL5+hqZucOAe+NETRqTVa/PwIUsOcoc6J8pUPwO0y+2x9
q4fB5o9857KJN2o8li2B/GOKUyTq0CMtXIdwTngIEfyM4ikMpS7PPHifeceUvRlqId2X6gLNZWrL
rrobTRtvhqNZdJuopVXRbGRpxDfh8pKapMkWl5izGcyPC3lKB0OchXKVd3/qskdD0FJznO7l06rF
lGtbc3546bIW+toIWaNB7BWqDUi7Z/UzZEs/sk/Dpx7Xd+N2cUb5jPdskSFSmK9QvZWO9Vvqn7fL
eSCdk+F7OFD9tnNEXp2GQcrCTgXqJi4scHogFt6+j6vxavyhI9aMVAvvy7RuD9RKZyosgGFC7O/B
2ISJgJa2JNcmNrRX8xIsnBp0T6dAFqjGlRFIyv9Cq2RDgW+qnzQouekFp5wpS29UxYDEpYdDeQMB
7gQISkmuG/SrWC3RkeKvcEHOFcF8izyr6JaPb9bcr8tZenM7oEtuhPjL60I8ANdzdKTnHV/UF22s
hEUbE1KQudl+QqREcGVxfTKNu15hpVwngvVnnFdWyun/iVojQSTxJheoJUO709pQQjucU62VjVam
unl8yi29kcl4c//U7U52XA/+GaWYXQRjXHuN4Ue7wWQDz1NhhcbRN+srbzj+qFbNoNXpk2RO4Bw5
Pm+3ViqYeIyrv/w4jfW1OGOuLk0h59fX/QgtYQsBertFO96dbwTn2PKKRR+sLqiaddkNF7ZEfxxJ
PN5m8sbyTNvk+TY2gdXjXpI3uj3ZmZ6B2l/qUzC0/sRpPGUYkUxIrED+1aO+TvgTM6TH+dJaWmp4
HMnUMvJMGrKFnSFykHROPVmJTdgD8wTttyqNBtyKyka2+i4c4yMC9pLU8/gEszetxWZcGCHcYJXV
XgSK6BV+MO9dqWW/efsOfrvtQDl6ryOXT3ceB8j7WAz3Mn98cCQKgmwQivNjKKTIZhFi5uG3EERy
DIxT9R7ddjCKvMax+7R542zKZFw3png/qWIldcUKESeTqT3dI3hWCxulmBqsFKWKQzseJxE0LexY
fanby2JsjKiHZW5pNA7ZJX3mqfjdL2h8Jjry1xh3C3bQ3AtHjmoVjj3cx1yjQ8Q/W5XOYxgg6t8p
MRoFrCdkris5mMas9QcmuDadV3XUZmGzUD8fH7j6I5zl1U/xNVmXP556pHw7u3AJUEBsub2Zzn8q
H/TlaPoZuxnwvK5ddHzN9DTisc7UIIGdcOD8bb7SpF1o3F/dDIiGTYS0wkaU4Qz2EXAZfJ3MbDqU
BxSsdcPs1KK1o/pC/d4PgUoQzWUlVhwHH8FrR38ApMak2iyxokHPy+xCQC5GFgZz366FfOyxa7O/
l6+PsXRI5s7wxQQWB25LUyix07uHwvh7IpVvOKqwDIHAEGYFxbfpnhV6/NZOpZm9ott/+yKjlCs+
7gBGaz30FnaIp4kc1rzy+/tR6rtxRxX5SpYHMiZ2Sosm8HPLZdSAPBv+LVU+gYaEXGrfVdobjHmj
GKQPRQOJIXe0fR1XmJBXhFodZ253jG0g+mlAQ+1WjUzlM5x7mz3vChByLSoRNpbrXgl33ZcNMRft
TJSrGUWqxFAgESm+mxaVv9kkB4FSz1h/581I8lbUrnGR1vbt23JDLN6XKbW9VeRzu0FzqOblFmFn
rt7oocv7gZuan/UwXaWi9F0YcYeIiIQlJE4D2/ei+M1Ncn70I/7u3WYDc9FIEWr4TW0rysWRkrL5
Hl68SmBEszfw+ngP9mQuo9Y9pzNGLz32ztx1yjpI8QmECDrtqMhU3fFEEk4jK+B/n/M09JW8V0KV
Y5V6HZ35gNT5SLLJqvzxA+VHyKAYYMuYwABMELRIuocn7+jedgEWU3yA9koXYUryul3V6N68gfBx
/OqJMiSp3E8opXHMvHjcdB7OuYXtuZ/NXC5+ySdaHOJ4wmi3kRElQYuOy596f0i4Iewg1Vkv9P78
F9v+EfMZyz5YMj/1pUouddMThtI2A/aJbo3Y4dS4rAuPwTK5LoxFc1nkV3PWHHqwnlApiwzCtTex
b3SUBUYIC8xtJp/UBK6e+vd5Amt0bTlWvOLvO5yr65p+d5KgN6tjCNrSCtnIg8BUxIFTVmG9DOue
0VnfD0Pi2d8tN1zvNESei9QIznD2DlBei2T3X6ay7U4QKG4kaswRA+TIbVmy2ifrpXPDi1ANa8um
Mr6mfviriqHovGWhc88MB+wXTFgc/bkj1ShZ64z43p/EH4icQ+3pIbbiQ9wAOTM88DMG6HYF8WBV
CqdhnKufU4QcchlEsHR2w6eJGe+sF9rDQUlLy2NWuKhHweCn3EK6zyiSlPBr+VGz/+T/r11J4oV2
I3I1Fd8ARSc8dBLaQGepRnBTCwe0myNTSlo077BwOJTr/8E9FdtR/s60if0/4mgDH2OKpd9DYNC4
6TPQGkJUZn7Y4XQH460rDp5Sjpej7CwtevpDV6mAjomlL1Av6aAd6oS/F4AiX19ELziMLQ96c1MX
ipjzVifpsIemZxl3A2oX0wNaM8fbBAcNe99a0R7sQsDk1cBVoPBujt27xpC4eKrPBV/FgFA1RWw0
+8FsP/Z0rQSVIpSXoM7SjmkQVwgTHqlzgLZVGDSqpCeH0gsyovbgYLxtpup4I52vmnWPiKQ/C3nA
PI1p7mrkT7BZiJ1Dkr8kO18NWLu95IJDmw2UOAw6f5CVWe9PODPBoVNop6SNjJwbrTcJ3nL2rs8I
x3/W+IiGDYmg6K7FGD3WLRwbbn8hJ+h9d5jKjb4zpD5qHbFYXDTWFGtzpp+7Su4wZTtmIOBrOFqX
SZVa7hi3S7YiCR3yHaI5HdN0IBtFFu/KWu8feQNnBrAXuno4z/uovS8jpe5A3S4EMrFFIv53jim8
G4FEFlKl23E2xXzpUd17EN/DNwRPwhkXnKMv+XoYXt979OpMk6ErLUGX1T2xQ3y2Jzwlmvw8ZybO
eHIGqvSaR7iVRgte7EILcUBy12z6NwMD92qmy9pwIS8MiOFibaQfBFxNrizUPz5bcr974VF7J5gk
U47rLg5n39hNOpSsZPYyTjdxi4khHFJVLqNNo49w6HRDG8ckSCgNWfZtTQw2pJykjhW4dbvgVBtM
FqfU6XWnoEGIUOCJIYAWvBsHXgeyj5BuTENtOnQ7cfYqR3BnmaAgpBYhvbcspFyzLicJo18I09nN
GDMuLXZ5vSyD1IaWzC+kNvwZC8VyZe6JslvCNm0nOlEryHuaQ3lS7HPnnTpASfUiihoq76DQ2Yzp
Hw6aVs+vPlLU5aHTg75bVJhFYFsadwdQoRTmEU87QWwtl5la3KxKY72/kCXOtVOz4cU2JlNZriCb
6RHEFV9kmSolH9CQaZFnw9jO5//Ovl/dNZMmSoNlhwz53k0HQH10+3YYf6pR8A8oF86OEZVZAtNN
IkOwjeCnhdT9i0oazCJrrf2pSq1Om6X2iaDNXZMYnmosZcshDodwiRcjFIT9I0L+J8wjczlnQgkL
DwQRo2GrEezzDZy6gN8/VvW8CnWVDHZ8Ytg7a8IOFV6Rqv0L4ruuFan/5p/k2YBbh6ZM1VWT2JKA
NYkb7NHn/70t3q1PhlRPbke4lOneQFRa+9qdaIPDRTMC52ZSOg8i4+yH+oBOAOVJV4epe+dlQYkA
EivTCnxBmm2ofCAhHvaN5iIqXMTBCwy8GayVa8sVKMHj+rBKGqxgCQC4wwarEOyMlWag6gykH6re
vfcBG1nRxfSXC7joctOHm0kI7aU/LFelLtnF+QP5EaathlF9U46B+7doV6sxHxCTYVGvfZkTECNx
rDUZYsBKp3keo4rxy1pmDXgxt9qEQnxZDcpcnWhPXW2T+EWIW78/T/RanG2bb6iANEsywJ35gOK8
fiDao47xIXt+DOBzCMFuMxD5N9JL9PJaGrvcLJlJXKD5gpSh3i17+2DqkpEtQhVfcLCJnTTEcysQ
YpqzL0W6v+U9IImUJ4va1TiQkCsdyrWCGu89V/zR79aUkUuUemmUYriG7EWALRWkY5cJCo0IFT3I
oDCdp7zFxlcLItepMCkMkMMLIjLEKwilFOpMkgab4anSU+OMRoHsiJyn4sulupT8XtujEtzVYuoX
jukcTIPg2ADgdEZonbZ6xN/mWUiDHEaoO/HamW9+qTuHjVCWPO1ClfUzGnoVNFZRnxuw9kMDr05c
w84PBpY1chuYrirzvtZH02Pdld2RQ3bXPTnNvHl++MKUxMBBEwdRMoh72d8TrVSlJ5DYy0Gny6FX
/DMhA+WsY645uzCAY/YtfFv8ChiTYEkeg/PSPnDkNr4BgUstA+gp+nwzihsoE77AIMNFgUhS/XSs
Jvp42zepdchVgaqhCPeIXBREN3mzq/UUOPkwSCxVIqzLGx3vwT3mwtxFEAezaYE9cVeFGT1EXjNY
yELnitDDWKv8G6Wvl9Y/eOIZBSBDeqL9chAYlWxy6pL/NxTAcWA64B5T93w784rjqU/JS3dLnLbY
EnU33LwDs8UBiJzUs2Szo45tlGVIoM7CTLNNS6IsMGkp+y1F+c6C4rbs+Vy3AecX/911Vg+K2mCn
sPIDen479CE66iCFYV7WN+xNhtXUXoyPcqR1zoI50e8ekOdOf1BJm9bB7Kff2k4PPv2nCvhe+98n
Bq+GTzCUEIxxpI2BtN9CNi6EqoLyd/7Jw7vBMmrtp+/AqEk/tZX9dIXXbyELErzSWJS8MUO5BKy2
MMPOmpnKPoYNshh53QflLSiOPINd87EKTPvLKxSSNBDRpJ/uPpbWc4Nx07xVEBHeNsmxnsz5fj8F
/PB7ETwjpkFEbl4pZs9PnWH0HZzJ6aTqKTjSqpz2HoMwfEjexNky6C8syNLVQwZMQwuYH7ZrWIkI
diX6lY1eKqoULiCCH6h0jzzWJ0efj05Ro7kF4NAJXiJm9LmOvqnEBHIX0WzsMoJpC8i4SlKgS9pI
G47U5K50siWh094XVU/8q7AdKXDr05Kmkp4ttB9FjadGOVUavqb1vwFMboRP+4JpRTQpXOdKgbrT
0IaSHt3iU48XvTs8ogTDtNKTnZmUK2Iz4MDV17LSXRr2kjG+2zaB7ImxEkFpWiEomGhZ7ojQhC04
XFZA9wblmT9H1ADqRzE2Fj+gN/Y6CndIX8ushFqK3I5ssn14V4HuUsjlrf3N4gRiW7ADBSnsPbvd
Ejc9nd5/EOBDIBDbfUXYkOIdzZ6EGvYEquLuc681no+pHqLH3riCl4cvOXI6LgytsSksAo1zJG3K
7rA9JCC52viEGXB5PPg4NTSdIcyEHZJZ+TtqBcuojkkBoKSi1ajk3U75+69E9gLcFeEcqr0qKHi1
lNUCl984LtNvJZPDyo1g0YxhFMBTzU7nedoqn3VzLHkuI1lO7LhYx4fjkHNdtWO/dE4h5kEsy0jl
1HvD4D4WWIc9FBq5Q2H1RvdGWWG+p2S/SgU9QTTIyG2qr63DjN4os2JYI/1UyMJ1MOfzuW6POt9y
H/kUZIisf2c5Mn8m5PPTrt/I8lXAd4hDLzVuY/yIpLiSavB3O65gxOng7QyhMJ6HQhwJWUa7LA16
olDXUVMjinimDnJPiELEcv0PkUVT3M9sTffbCwqHmXcjicjLvYL5kjeoGSRHrGdDLDg2BhWtyxwP
HY2sDRAj4FksqmFhskk59V6s1NYt8wTplSYBJD3Ek2BsLp230Qitqk/BdyYOZCe/Nj1F0m9JwoAc
QC9R3J4by1WGeBSlLVZQV0Ghfy4DccnXLO5UAPTgNMVOYw2+ZTObwZZTVBnBWgJZ9g0/lsGm0uWX
A0O8V370u3rRsydD7b5FYottKgTlqPm8WwKToTiNH5mtac+6cWUytV5JQyjfPtqRbg/khJU3zqKW
Xor7mJuqXSG+CbIdbRQHuac4g6DtC1OxCfI9848LDcAVPJbODK+8k5aYVVgdiHm228+ANjU/hWvp
uefjXapYpfu7obmD+RZob+lASO2a0O3x+I5gGT0dH3FoEfyaM8yPzaE4KHXXOO7FO8BexrCVV0fD
1slpQBJGUURBWxEr1bJWNwEiwZxICV7SjQcM6jGrDy15rSJI0VghGIPR3yJxIDyZrLTJkEcNMKST
Q4Gzjswf/jYTscUWBhm5v5yc81SzIc+ERqvjfnJo3QZgD+DE6q8geO3XLPq6NYtVzJlDV2AGrSoY
3/AV+AOZvOt6gbK5GJLqwz7obKGMpuWyzdprmNEIQ3dx73EXclonVxST3gP8lByuVvG0PA2a87a9
/2PLsy2H0SxgHJ+D6C0Ql7FxKkqIuMfpRcsdYiyDyiKBmdUvU2Wrbh/4XHGbZU0vjLnaCc+eycil
ghfIFrEdeY8sFi2NM3dpy/G71T7cTkFX7/5iPzNJN22QXpLBpMw+VhBdPE80rqleYJJTJgJIppzJ
76f5LVnuaxTr94WZh9VTCO/R7DXJjcCHUTnpQ859Z0anFNHK5TUJw4ffTxCMsefqlQspFWVUsJ/G
pxIHWAKND1MCAXofy3l/+0dZhaixuLIYOwS4ZbAQTJoLDZhp93uTiadcqeZevnStE+aU/qEtnKfn
pBmo/fTOVrN44qj1VRP4OBCrSbONVLfynyko2ilHL2kJ+TGW3T3Wr6JsxiBzIyBaxNS5DlvssCKs
2slD+TiLOCx+RH3mvz9aDRgbNNXkSqvOl0SccHd8yLEffMZqMt4agivzZkAw7vfjD5oKO4iJf8Br
pFaK5Sdn23kcucKb15mgy2oMw7DY8h4Uk1IkrkpVZC0aU6ynKFqVBU8Sm7kKAQJbM8m5aSuUHEPy
9fPglQ+p9EwOUsG2AEXZKZYRRPhbYyjLGrHtiOCJkUiwF6K0e+39XQ5TtZ/9nSxlUIalBZ1zMv/0
JlQMYLASaiAbfT+vT1KuNvhp4L05d42/sVaZYEHvkuY3bn4bnT2xnJJXeBRZP41cIw/qMjc7cpy7
gNEhmsOTkQDJst1rpoIVixYhLlL38MwKd8eadJKO234OC2isdezpn0q5E0D+qmW6S9OblfFyzNxJ
UObA0a9CFLe+J593F/aMAJ/uqJHgvR6nLqaiPsj4edUKZw1E1sjC7Gl+H0Lm+X9Q92cXWr1MhpDZ
e7kv8/01mHCZHo8brJ0YPZHbP9MTo+f4TSwAPLw+qTxZCbk37MetAMPxgjS5uoY58ZYFJfZpzOiS
HXOYSrdYksWCz5su+A4j3I1LA8AwnTTrjB6Is0zDJ+JExTeFohRd5M9efvSw9rSc/WlRdRuMojUV
H5B7543hYLWE4x67iLCJ1oUdMDXwAflNOOxp4zBhkwpuRRtqXnil0qBOLEmb9yGYsXI+8KEhOnhR
Re0odDTIbcyXv5sVwr8st7WP+Dcg+78MM37bRbUA4tJamWrE20sAf+ZsprIFwo40HldvifHxDl7T
v/rV+BUZudplPj3p2+1+5EeQvFpCg3mdtJUBTtmQrWAlrfFLWyPDEuO0rIJ2hOF0Bwp3AKTlW3AN
SNLRIFiFgIp6eum9VCI+jfQ9LXFBFSG0DfNBVCLFZp0aologb+JqgsyS/6ujXfBlfvaP6eNYBbY5
/e8fmtvzPMJB+0xgRrq2Es0DCdT+mWxweNY+94dekQLjQ0CknyyAT3hPhPUxF3wiEndjgVn+22Cv
U/q1OSwUz8irkdOhIeEjqL21hw2nakQtvZkpniYm3VHEadf41vFK+K6d7TAX+fi5i1qcEZfTpMMM
JTEjX3DTLp1OO9fxiPbeWF+vlt4FsT6okhI8DfZwlMnYykh0VG5DFnBJaL0m0DPOo868DVdqlbVF
rwle3nqvyrjncveCdjzhgwJcRZjCZmIZUythMB8qVhUmKGLWKYt+7rAqHVVnEhmYHs6WP9ie7B0D
ey8Nsn+qvUCBPf5AdG8W4dGrquIRpcjtvAGWb58Fr6ZDC1yfuQ9oqCvomp1m5ohYzSIly8gn6WpG
lm7pfY2NmMYaVVY77iN903hA9RTIeyIdE753F7U545pL3BynmUQ0V9WSifvSo/9O32o8qjtZenTc
sWP2DCJWJCakYXO8e5y/Mr22h7yYuWz1G15cfNwqzu7y+dUrR7veiEXf3VNlzhv+uSZvpw2DD41T
vl/eW+GzvN9q7ec30Qw+yiDwq/hG/i7BJQjqS7xdS9jU4w8MzNAfKqHIqrThYHreB8sm2gJ47ffK
TfIaG8CgTwMp/HH0hwglQ3S9Zqeot1jt+Vm48rkd+x2+fLtwu/QquJgHU99yh04Ga0FTscFWshJE
5g19zPrcLS+YYjYlDhDIJCY/gIJO9sLu8mNklPV+6DbRi90CQ6UWBhnjuJwCk5Pwol0gl1awvr/T
tGYZDBr/bGdopSD8f/p2Dq7arUf+2Ai0vvB3jYiQUpRf1MsnNvIgAPXRRXdU0rzE6rtxQmuX7D7d
+gjsjYviUrO8RPewu3nF9Ao1mw7Fqrp5caojgLJRXwOzb4n3kSbyGdSyOf2szJuf3/E0/YHsNd5o
1XlG+8zARTd7FZ1Hv/DqE+trvdvhmmaFvLBz/3gBkTWIyJRK/9swQArg0utedWVNVKz4Es0LWms5
pBYuh84UIqjLPB1s+LVgcJUZUK0XD0l7QsDgq3l0ZrwVt2CMZrWVr7JSzYZnf8WXM+4bOz1Pa6dn
vbGMpCHjaCFIwBKFfBhlyK1DJV7aaX8ky95a5gUJ/AP16kW3Mu4fn4ixB8JDrNIPoOKs6CPxi+vP
5NQ/x43YBDMyHHnBPmDDEQ5VUpfMXMAFehVYDB/2Bkb6GHhFr2LIhXeC6zkIVtVyOqMd2mSOJAJb
mooUitxsdtcY+HyefL9yehvOXLc1UOJO+1Rza6gSG7v35+lb6Tme7nfdPIwRu6y6OjYcQKZfewTo
Q4HiW/qggz4MWPYx/2fiYdBGgO4sNwCoV0gsFppmLs1xUAGvoq4Da6jhH31ydoTHuR4Gjk6P78Up
srCSnEZyCrvrKHOrYUtCbHniQeAcMFb0Eq21bMxxxACBMkzgoBEqw1gcq3WiSxhinKztbq1a4K2y
V4cqQwXGPDAYoj4ottNdWUdxgXRqthqA/tvX0+TRL/1onTMC+uBlYAn5LBRDehoUyjENCH/gdFue
ejh0ib5JhLNflz1sk830+6vogvHCp3aOGiuYueNCz2LddS7zpsZiysy/Q8JxZ0a7eHETJVV30JnL
6A2VIvT3A99Cmq3sVD1wiTdBzXW16lGysWCkEK6bM22AaxCVHRCXHvYjtp/+nzz5MZlzu1RZsFPe
N3f8d611oHXD8eSlmNZKmUWePbJN/EAD8v5ULtHYzyo+1/JXAjJDuG0VoAkt/XPEgVqnVNeKJA4w
oi7SEzipWmOrbXRDh9njcofdE5jmbmrdkLgwl8KoY7yofghMdomu7bahqVDqFfR3j3E2Bf0X3I53
0QMkfZiMLOF9cWkp2awMWQ0SuHEzDrTdWemJSLZP0/DmwpnhwIvi5m9/8LLP4foP1Ef+lzPwKBAs
KlTW9KudARzghQrNb3tzP8wkD7SD7O+sC5jlyGRI0RIw6q/SHAiaoGb7PNccXk34/RwG+6UGI2sG
jRSDWm6gl+hGLywWyLkDKWu1HS8Xyx+Cnt66TRi02vA2lfTYCl1JoOeDgwxOYAI7EIqC+vG/4rLN
jpOs9YUpvotRRqnq9IwVFjfuENTrD6JLJ60mOCMTHFnbNNQHRe0qJfmi/FfoAoJILnJoqfyAZP/T
sNVwxKUffJ3PK1pkjLZSn7uZazpC9oWeDbXEQwknJPHKr7uMBpPGEKatN0Bkf1SScp1NTXmmTp4l
i9ZOPrXCmvHNUSCKrQYeWgTvTrZNZ14wdOdPcxQ1fwGleSR13FAyxmEMi36HuPi2FRuz/T+UTJuX
jRh3lgHkn3tsoZuo4hlbdcRI+umotURAtB79a+6hJIJvaHMCkxXEAZbcWoQcD+YRm8C3ABDfE7au
voCsl5hvGAxUZ4GQ8DSvwQNPfA6ETWh9EdXpsnMtrdvx0A8GQD1dSAjpyhX0BpH2SLz8/BLas0NF
K0HQyc0gwfMipzFTAbYuTV0jGElKZRcu3aGsaaGDpWb52BTA/r4aYHOHYrCTxeBA4Aq6uIOVUR2m
lsyvnjNyGrbqKii45CNYc4HNuPk0mrDNuTDeLSk3MF6q0Lpx3fd+BeyYQQOuv7R3gerG4G8+tSUp
+nbikJMgSC/O2NM5jz3X1PWkmPMLLwXeKoirpcXuTVf421O6R8njkPiwNwKmyLqzj4cM3tKRrhAd
nLCxYT4uL5y7DXar9vscTINtBXbPrcwAHoayr6hFPeCwL9V6yMTHOEjgRwIxxLaCwlGp0OAgjmU5
/1UHaC64eTvRIbcuFIUSL764VA+9szBHKjrmwqNtnw9WvJCY77uEcMiBEF/+c9dnGTFs1dneAQ6R
HQjg/WBUIw7pJEyt+ZjeHaNDdHLqqD+gu8Wz2Q5eBGZ1qvaPEiJY1Qy8JKFJO7j2dywXjtfEawKH
kII4IyUacyRtkyWJK00T6UjB14EPS5S15cjONNF5c0AJ+YzEXs2XYbSsOClQ2soMeZComiAXAe4m
SSKTvnNfQ97ct119gQDz1CnXhUUIaeOZxFtst/qJv49F+vdeCEO0j9AwVfLHQWwokHl3khxPHUBU
vJwxPjuTFQ1bIBQu5pGbR2MOKn/mjyKYaIMNSY3BqB4XBWKuSfu20vVsiwv2wj1GWp/Rgy9XFc5J
7AMkH4wWtp4wNR4cjGUMvZ2E9a6FknJ+Nq7UUTtyXNpSzLaJUUzm5LLP7sAjsOCzqXff5AH6gGmk
2h6r7hfs/VggCw8JA2acu/Fa9T2yjHzNuDRSDi2ASkGbxg/HZ7okfpvZl4UFUr3diJCJR4K4xcl2
TPiK5uEyJ+ll3SZTXarJl0k+C6B22aRlLuVkGjhbIxzrlfK5mmY9y9zbJ+1MDAfFjJmKCXvHdRGb
FEsYsq8gLwp1eYo4+WfIgl5nr9EZ9lReqZxskVDXK/a0Zwj9cRZHp8OUr91siz2Csa7a3z2v/NzB
DgKChiDjs5XTHk6qWxbtvi8jm0ePQMnXrDB/gfi5d2RsIINi739HPXYb5XegRo8eBF1mQLY3y51H
ye4etNtz5jWW/ORy8xvi6JdHtvTnSlQMQQ2vBmruFC5RDl8NUHhdlCCik+6ZZ+2R9VNUgOWyHix4
uffwRPSiUuasGHSx+1orJzK7xfFPX6mSWWN2eqmDAkIfCaoLpbIbUnnA3tQr7xHOByh3rpjV5/AP
ZD6u1sH8XvC3tju+T2MK8uZVcC6jLgD0TNFasnZrPtEWEP6hhd9ZsBS5LbuA+sLP1s3JwkKIRezw
gO/4IzqnPBFmwwWn80X85eK0U8cm+H+rED5cx3CEdzbIk9gY5ZU8We6WQt+k9mIB46rs+SqBCM7N
cjOh65PiiZOZu6fb/FPXrjbTb7Ul9TBg1aol3CvShQDZnPIUVBb+NP6Qk7RuPv4DFpOp4vEXQ87F
g8uVmGXVfQHEhyXD2OV44dhTXrSe91lWMUcuf5deWYCnANLc25RT3mu8V4p2bYzb5S9iyWRhy8La
Pu2pYiNYbU6XHM9ZtrAq4/pE6ucyTY/zbw5dDnl+StE5VaF/wyiSZSexh2+b+mULUaURijFXNLH9
tsDMzcdKm9GULe+kRcG9tKPa/SFhQRV+9HMnHHcMkiP/7YYRWqQ1grwHF1CmAqZEH6CRpF+7y9B6
yWg1wWDvB0m7XtwmDxXgLwDelwhVDT9XC8uAtKopKVGXlUBN2k0P+M179iMiTXDJbm7R5XYsw+Ws
IVaUAL3Z0Zg7fdEb6xOtyzI42RuPHGeB0X28VTkLC36nR++jch88OuZToN/Tfc4iogv+NxNs1RhK
4nc+Ezhx+eRwjxFP5peKol952B6uCtiM5QYuqLFfyP/IFS0LA6MIXrZ+ITYPUwn7zbpUpNnHbUQZ
8XxmrVTscbPizBftXHCjPNazu3xqFVaFrgxv5ySEbqG3d+cNg+lMc5utaPr6pm+UX3wDj9hmveYg
ixuDDdHp77YphEgkAVpCi7O5+dv+yKSXm6zk1q0HEpcGHme6hwzSVXDn/PGE5Ctb6K8ubILzbGy+
ORC/mlwxFyrwMJQf7d70GUkkcARb/fn+EknKJr8TNogTRLpSnIsFVg7Z6aektFMbD75NPggOt+Xs
9q9JtD5D5OmAh+MLL3alBcdQoL7gpvW9LAzNRHtWwzD/fqsDEnLPstWASn0Brua3M2PaPtjrClkn
+xvKWSuvX8MgwoD3p002JWQax+ppcuBsHj0K4MVDi6JfuVb3ejvFK42EobtI4VSeu3Kcg0mPOe6l
EyGchqYpdv7/UOdveYCjz8uWZh2XFOqJOQ/VuihcLiqnoBnZgvMTF7kd7Lhg5k0jZ6gLCZLZ7Zjw
/BCwENIiapqg7HawEkJ1IXKMsnr6tL99x7sEQKlvd0SrULs2RrBVNsJmY3FkiXCmxcAFHG/h+fV0
gNeXkNlc1V4ccbHusVf5w4JG/vq8kLquO4tH4QCIyh50x/MvwV0I/JeUa2vetH3FIgcM38rxnKDR
x5lEDwPOOU16Z0sf62xTgYSpukGIME3khJyvHcBgJugVwU6kPixvwSGj9K56GV0NmUGHWds5Ry2v
vpEHQDtP18RHHzaD6OTmN+Wn+9BJXHoF4quvGk49QOKG/W6+valtPOyquCnaJ8f1GmGcSGONhPRQ
ShyV6CRbDpMlQWuFsnTvXWL7/EC0NN+YdC5vcDNICFgUkcWnDOyOWAFQZO6M7HNI05RvCrpRXDUk
HgwXDB2DnMKv+zP+YxhWmWERFEjJ2129jSQHnLmc/rIDB58YYIQbwg6Px2zwvmBP0aAlD5na+M+P
AbfMalfWRupmlFks7rfeVY6s0Jj3+w89/ZwoDBuUVFCBMoDuJioCeuHNQPhUiwxdE7+icA/Hl12G
RHBpnstEV2Q6SyXOuVKaRHAklYdaIJH0VNYz5duT3RmH/5THbwp0/sbfxLazZImqP0ogVVaZ0SwW
eyGBCaGYB82WH1wLKA4nh+/qV75PoqK/kujN10RbKS8aZx/TaBIS5ZKKenA/De5uKYp6x/dbEvTf
RDtSkRFvSloVJW53CfL5gRnoKulZdO/pOO55L4DFT2Ra5vGhrdebU0rBh08PHlREmNUpxDzVoBNu
tZyHVZ0nSinvSKPa/sMUuZpLzgWmbVPjFR0BdSrld5cJNMNHrPEdmFyUpBvU8KdM/q0GQWvdEs6V
I7/W1ueTjKkJCpA1SJwtT3q7ZRURpqMEalcIpYi8efEiux47jZxEMCsKh+aJgNmtk5Dcj3J8ipz0
xzHps1YXVsYORaKCZbL37QMGFDB146BUoS/D52+R/oQk0qDPn1F7W803dVA5chQcjE3Ltsm4vZ58
3McAcNeG0eOH++LsCnND5UuTEe754x496tckB1N3iuhP6tG5BFaXWeXXVvXwvJsVP0O45k8kxgt6
ful5z4K+wkDc1Vd0jNQWx99/E3dB/BGMK4Ad9aiJJ5B/B+J6BBF32ZCXAtRMH2yaVl9lBqplXtEp
Sl5IKg0evz6t+7LsK0lUx5OmCDu/vRI4IIre76NFgYzVyM+UlGqEr93r26ExkJb+PwTrZNQ0LyeF
j+pSIbZXu8g/UUEF+LGENcAQPzS+Iw6oSqofDIGKJlNkiWsJGEld3FmJfUlIlrnCbS5jWJeBBUO9
3/WBqieECy9KVzV2ZiCH515e6M53LndN6NuS/f32pLl1Zl8FbJfclpwgyM0wEUH9/hyaAO6WfUv2
PStedCE4nB2CG/KKv1i58/SzPKZw8qtxlmLvnmmaDsCZc1VwfYFdjqRwfusz3h8GQR0ZpB7aEsqe
VO5Oo8GZzNySnOrPhnKkdtEjs3nAcdtqV+t3D/MD6BFUsLX0ISyE2yAE3IUbKsaW+KkWn3U4hiTE
5PTmmbIyGudcOz+/uQ3V+AdzMbxagj+edZQ1mjd9P+pzwdCp4EP9nz8wzmK8cVbQc7eU7WshP7mN
dhToJ0DICJ9Ls6JhBa8XXucVWwDSBuMm9BK/n/PuFiaIRpEi47dEYZFB8KVHirvLjqp7yV0t5Ozf
cnkuxJn8LjDt9eL/zN0ZRUmVVwPRkw94KX2O3vvJbo8BLPcj+Jje5nze1BLIwSQ3cnbGIUE7Prey
sqJRh8KS7w/SaPZoC9PA/HDjOHzICF/Yi4uxwFi2utAP7O4shF1PuhfOge1kl9zw4IM0hHSByBJm
FFqPepMyx08LwLiN+GCj/bjVIBStd5ushdBIh95vA/WorheC2rAqi1O/fVAtbwZHaiJAIOJevfCZ
xMz9FrYMbYxAVh1Ir5RFq74tYNCKeQcmvSInL2GsBk3cOcXQglyoQy8rqYNnl1KYdA5GRvF16i2j
chtg9cQjdR65EZHHqLEAj/yVywFdoWmgC8DK+Jcw7bFs40GHTR2Uvg0KxufYtQRgdLd1Wtdkd09G
bVZ3uRRjAJcUHYWFDpAAm8NAKteE2PFP/ZizfGL27xQgA7gmc8gAj5hf5IsKEawUjvhh5A6Zu57W
Eong6KepRHYosJ5nOwJ7UtezRL9bocjMZk8A/sEaKTJmYtfhGFzD4T0v/LSYvRn/XS/C39ocMx5q
QCv3rfLXeiRux1Bwc86yTm5WOwl9iKJKEDFbdg3NH42jUAVkRA77Em+m5yRfjsLqEaR2QnOY3DL3
ThW7Cjks1sj2NLMBKP8KVDRpyoa/qsNh6x2ZvUa7fYDbBhYADciAwsPov9Uxf5MvnM9MyBQqlQip
REdn4K70p6rYWGmdSYcbXwb5zsoxqL7B22CLnnK76ikilSyRrMg1kkm+BVGns7xw0rqd39n2iyag
ic0K5reWekJNLkhAyLz+ITG5JwRo1V3yWdoysgh2bAdkKDc1o6RcS/kA/RShibMozcbVS+2v8w2d
DIqf1jo7Dd2u+0XT7AveoyG61Wcdfj0SBj5fxrb1ImsMUFt4/bIjaFm/raI1X0uK2dJGrZX/X80s
4NMm2dh8kXzHABafKNKHV2vunL+tvt//OfrT/qjzgYaW7CsFqC8+Z7Pf1YL8nldpSki1W/fAD7SM
W2huDLnrAa9X/KqQknn8zsPrD1rt1mDgQW8gxLGKwCwsOdrwV7k+h2O7ZdudEvODdUh3NYI7da3J
6qamk518YU/+DmHZPNdJ0qeCHOBe2dfpvdRnfvcVk6YocfVcRV5rPawPxh+rdIerz8q4hjqDRlCJ
YGwIilcnykWW0bZGQZPz7HsveKtx/f0jb49Cx1VUER0Cw7TInHcBq77/BjblGpzNycdeiDG7vvA/
nn1pqdRWd2MJKeILMh+RMAbjavfmoNIW6xjQKQnJu7ecJ9z7IjJ+647p/J6yet7j4nePWiLHNINa
Et0FoisV3pR6Cf8rNW56dBRHieMm/ZzOBYbBnfezz/RyQa33ffb6zFYKxMtm61uHXijaADUdxCQT
ACyvRGKQUZh7yIDeV+941ovubPBX0yOrt01KfeS1Zn1aa53QjSBaAN+i6b8VPCdy6pk0ocs0TY23
gw/w9f/bolqXeCun9+NeUliYGVzADwYOjH8k+tIABtHyJ6vUMYTZZF/DVs3zH7gqAVxnfd1Aa5av
UyoMVrRoC2LmSsMndrhfymvvLR6CySeuROK3nwBHsAdi/ifeEDHJGZwiE8kVok4oXdAuVtaWFt0h
DQVGFPl3biGF8LCpcRh920Ne/fJNoBX8UG2VZYw4oUNJSRHcFaFRvpuMvf2BL+anSUg2IH7mPpk8
CoC1bn7vZ4m896lONCkFaW2fUAAtUmcdPV61lCxxAMHcyMcnRI7e7PHdZ5Ni2sKkNB9uJqpgsu3u
8SySIcvsOu+DX1I32wwfhvitHlDthQ6dGoG0pgrEJuTQKw5Y4wpsBtOky/49zQrY0FyfkilQCsC8
lr2/hc/AyDBrBwQxpArMPUf6TZkw5L6zjiFCXtatToHhvwiUkC9KsOLHaUunn15uyfiYlJNnsfDA
UFJ6UQ+rHJNOmUAb7kyWWKHh4rdqps9cwoW4iAF1lJtc0E5p6M9F+FcVL3lnP+wF2tGz/zzezgt/
iuhEPvhn6moBlCPM0OkeBCUkn0BcabKMcSPx7tT652vVRQxwQhNfhNHhnaxyeeB/p2nwE1xtH9HT
XzRCyzDg4XlNwKdf4zOsNT+wf3RqCoRuXukLR3Ob8Y5DfKZLJPk1PoY6y5FA5/KZjOX34YuRcpDY
kLUmjDlVblSGP5gpGvhP0VYLx08cJSpkGJ6gA9L6734oosx6kTkaGNfUh/JSgYelT3Oyp1DQrZFB
99/8ZM0heY4FaJRRM3XrdRQjAdJfIjfhRI29OyBeMExjLAfllXO2n5He/9eemSFGiyLkMFfue67s
WuB1d84yA7birHeNTEbjQpmws9FL84ZdtHsZn7MuiCpcvtyo50mzmCAP9cndmtb8JUngvnh9EC60
XaG2P8WFNhhE2kJ3jFoFL02MIOudBpcFEFo8uANO9dPOWqIOJySuA17XRgj68af+O7o3rO2UnaTr
LH3NqTJgI1FnhqYIPZTYo2VEzKef5Q+SXSp4/8ajrT3d9rOaYLdG+iNSfrLj07CzbH1EKq6IRhz1
d45D+Jl62TJu1FexbmzI1qdyurbJrus+J8mP16Ag4X9dFURX+mGSOFp4q9wZ5QRPEOdG+edG7ZBn
csM/oaGzxo6jq2nMVw3eXet917tM3xFKwdDhjyKy1URCzGeRw7auDFyHLfI1qQnBhw1eOGVfc17G
H8GeET7bCubjLlw7nlwgAZUjKe9SDxF3kmKtlhYnccJFBbYDdzctw8Lf9Z9clRrlKn+DeL5Qg32/
s2F0/SvPrwecm4Qju5+I40B731AT5hMZ/lh6h0oC39C2X2zIYAXYFbszuQ0bgmF1KAXaIB/2G2ob
eYe0m1qLfQoNPnUVzYen9Y1no4UDBw0EitkWyhERa++tHKbiwuTY7NAFvcf28oVKVjcmGSV2iE7i
se52KYRAzpoNIis1zex7be9EIJranbV3nxx0RRVbrqkNBZMPZPDJyoKfUCeJFUsL9LuaTjRT0PIE
k2ImuajEdeIHr0bV9E8h5fn0OZbbmdbjnjQ0ieCnA7J9vNK+ckd0D2nqf4MtG22oFA/DYapkExjk
i41Enc3I1tslfD3jZyMCmCI2LcP8MUhz8/4Wbg8xGz2Z1FBcWdsKDOkX/uGRTsax7KVEruqVbn5J
r8oh2u21XfcxuW8uAkIJUZxB8qziHOuI+okzeOqxcX/9pZPTfgTwlR1K5wISo1wjafIv50TQizlb
ZCtjUlDmIBImLzEoGQrIiz0KpDZtCiwafDwEVlU13CG3tOnUbId6EFamLD/KJXuvD83cRXQsLgeu
4eVMvijprmKpqU5ezFYQkqPJ3ER4CFKTygRQRKcICIZE+onEgAur4mjNs8T7d7RT0vaYwFQ42mId
Yr3SVXTPaJAgT1+WJOFHhi5I+TVrrV+hhQ9YmwgAoi0yNwtRh08BEB2y6YwhNBc9+/m4IhGjdjWW
k2PkXes+a3iB8QQhtdk+c36HUFsqoUOKDsRCEripNGmoemm/KcZxMFZAr+EU9OojF1JpqI/EwAw5
oKwk5cDvKnOBXtDAUOmt0fd0lGgt4ZaBLiir0f8L8Hhmnut00gm4rSBEUpDHuZ+rgKPMAU0mwCEv
LlAOpySvrmi/Ft9Gm8X4ZN6m8HCzCgexptRT81Q0REIGwg032ufqjAip95ONhk9aEfzhyiU3uHsy
NH/6RxDw2RENmmWGblpQ4IOZi9KyzgDlN6t8EunO095FNWnKd6TnC2mfBFtyXZ0VJCF719Ok2ugD
xK+f3bwVUNdx6tOcFU9PsvNHYvEzLHxlqkp9yHmAt7cZ2TfFKEdOVRNGZY8/6SdekKNxcTELu+/p
X3J6Poqgwpozs/ydz0hNWU/QrCFTDOUQlimmQmBNasXarTUfHBnIZRq6PhiVMOezZdh/Ji6+GeWA
2Cb/b3G3vU8JlUoXZPpwpRmbHDjxRYzL+sCuTX4M71SWzUXcJAGhg6VnJ/gPP47YdUtDBS8QI7+W
H2rktQYtjHOy1u4+6TIgkTEPVrMPCy3hrgge08HOU+dF7wM7konL1TW2DMgx1o1DID9Y1nRU1tD6
wXOGgXKf99T4zShzriZ4rhJ4QyMBQA7in7ZZwx4cPqcK6cpi70dtxOBrCCrgmbQ0CVtyXtKF6wv/
eMQjoSE77ejulkxFLLx0PDCu/p3WPpHLXqQXjx4a0TLuF8A7EsQ6O+5QM3Lr889OsO60PW5gstLy
afJ4JedMTBWENWMXniucQU7RgMXSrlyUvgAFPJW6cFZwhKZJbO+1WfV47DUaJUlhYIiU1STtqC2D
GstdF9/31ABhWPt6aZWHbEHsl8Z3tpsy/LzyjWV6GHSQAK+iN9TCU9cT8aIEgCVbsN2eYhhlOGHm
ckGvKEb8upZNTbl2R3okvaqjxzMbIIe+8qRw4muDXdXa8LsZshe/g3c9TwPqfsCtHb37ZVjscxJK
45OARVhOJgKvMGftYV9AGKDpgUym9RbngoDzlVfXaOwOQtgVy9MH0v5/rMbBwS890xoyC49ro90q
sFu5FkUAjnc6uX58QLObW4Ky/7zBJT/mxfplaZEwATUrya6Bzg5u3tErj74joYgqYMYdFVDXWALf
x0aUbocOjybTzDOH9tGjij9zt//YXds3vbxguWj6Ez2/+jEJAJSj/iDHQrjJnX9HqiLHS0kT+py0
Jp5rrvY0nYbCXQ0KK+SLySYaYKfem2sGkljQK8YIyUNi2tbo8vbVBcYc0bCiTuKcgfqzWXI1nv9c
O2PVv0cYfR1vbQvmd22kWwck/j+iXWQavsXjpj2DoKto5cEZre7QJQcv8cl3V3lfln+/rDM4Iqy/
L5WlBPYcnKTMWheOZ75UK+blqjDDwnq0k2JaDz4t1p1lUPMe32D9mZDehrFkFab7ua4GoS1O/PSp
5NY071zTLxEErB+Q41xd+CAQrdfgO3QQtoHoUg2rC61thsZ0dLNkeEvV/5VfIVNZ5mi/8BNwx6TZ
wDvAKDxFHxUwGX4jCc4PjhPYO+wMDAxyodxPNgWnhvqN5WRw6KBGRmy/Wwu9WBKLlxf0kZLYquFv
6Z9rcklD+l/FV8GnpxQ5T2n00MVV2wdNYDsm3LltCSIYhlZDCUI6UveVdZU7pPeGRSY51Wo4F4on
FuxCuxYxZgR08qyYN5eMtRw8e7r3QQv1LFBzgniOMjOvM2aFuyrbzVm0xrT3j1/ER8+OZZm5OhV6
U8fVygXeZ1lG2RCwIPKeW8sTK2D1gREmBrCTAqmqLUjN7/x+N+UNjQ+MKMusp20oWor/P3koSaGs
FtHEDncdWC6tBya4iI7bvyoUD0dwjjTCPgW9Sz3/nfvfbOGJLf9yNp8/WsAYW0qhG5jScMtaOYQI
ay0SamDqYFSnciVXni55y2ZyXOWFVfXbK4mnSUOdT36HvgrkMzHMB/ujxUjU22dkkh/1jmSTa8eQ
aUZfz+tBEg9qeYvzD++4QB8JBrc7UStHf504R1Ae0esTdxycVCLZvh9hvs/quAkKbD9UqqyEmfEu
KCk8feZZL8zXcrt5/Qw+C7YswT2FdTWT1+5S3w+Tr4UjBCGYfMukEqYMm6F7xtUMs4oHa8Oisxt7
LEEDlybx7uHisxzTHLPy3DgLRDXfx2S8tgqP4PRkzwBv70cd8K5VWx87jFkiWcjUzyQmzxH0zHJb
wF4tUFXDU76UspLTSuCFdAFAFtEn8U31MgyX200hdicY+BmT/7M1uZS1UBtG75b19EQV9fwbgW8I
i1OQj3gF0EJ3FToupH6IgO987tfAEgCBv+FZDWkwB5w1BTKj/VVASviuZ2ggd9+wH+e/jm0CTHQM
Yl77TvvQwL1NPnuF8PfCPsm5pSJtt4hxQQpjtu/dWk7rmWULVGmEgfWwSW4VjMgojONBPyT/thqN
iea579MW0ZL7km6fFNN50sarNvAkziOucRgubQDFChwOV8F77jdVVUu83usG6GkOuYwR3MxNGXpL
dpQPilhpR5K3B0NWktEr4ZsL9pN4WEYamrVHyiXwJJ4KRiopNiQRbNHUuP72phDhSYcqsCdJ8+9w
0WKf+BDfsSHmsK/HVSFYZnMZwtvamzUd8vAp5C1wKoRW6gm6/bwWqkHLGNQ2jWSN4utf6Zd6zAd+
qKJ+4pC4jiHkG/ebV4QGGEOyZj0OGB/4++C7qK3dc0OHqUd3/Jyue2KS0xzpmAJFO/MWVhGMM6F+
JD/r6IJwGzIC5CVIMAh639deT+VhHLe3eY4yDWleNZ3pMBQLVfBFTEB2kx/djUCjcpZKvMYkFx4q
iTlFbTnRYF/pl4u4cGsvROEVa9ZAgKotMQY4J7QoCh+SwjHSI4JqHXUxA4Z/IzcKSDNgQ2i56jRB
NC4HfXK3APi8wCcievswuaYXgHVlg47Op5JewXXK13jz21bVtwXH5I5QBIbCb3zpj5Oe/Zqe0BWq
RR/t/zTTJcsH5nDku1P/X6FrxNHWtUB6MnzJ6AuX3XgtYEnmVvqsQGpBAiGfI+aTL76FaD1dMC+I
CgMtZlYkv3qufXlyokgslCFYJrEmf2DdoN3inGJpvj/CeOpk/hXljgvFv4R+vkexTdxJbesE+tPz
Q3I1ftorHsLDET0RcHDsfC6cV8rXrVDuF0IR7WUV9k0vzgHl+Em+6wpwy2oIGcKD2wMSbKLJQl48
UNBXI6bi1feyzs22yYYQ8c2P0gKMyH9JIL+cpWqTUz6GhEOkO6fZuMsuSBZTwfEGnfqNqaywnj0I
Sd6tBtkSaB+s6FeitKvjVYh7UX1l8EWPcBLsJbpw015U9JXAT6pWmuiyYIcntuMWR1VxN3vHlrdC
cuOuaEkwDmkZLGalhG0yVMiR87VaJGC2wtvr4OJzXXOZo6Lt3C6bYI0NQmrdNHmNtCRURq/3OSrW
SqSpuH40z1mR3+gU1vTJJtcPX30Kct3CRlt9xNaFMArHFXwAM+4bbGvj3YzegieWaXy+ija96mxQ
tfVGcokmWQq1t2EdVwcSznzH26ve5OD7Jtk9Y6htZvZysUAMhGwv53qfkA6bqC64AU7EGNTcHhY5
gXh/gjzHhUK8aTxm7h8tDHQamgoP1B+faqE2hChJIelR+H7VyGGJojmwa3UMICPlyxBuB0zDycmI
YaD0soMgbFimGKCVqhKzRn4WTOzLA9Nc1q712AxrT48+102yNw51bT0NiRzfpaG5bc3e/ZhAFAW+
17V/6Jy38ktHHk4efE2UAdQbUFHW2M6C2ds9lQ1+e+PKKOiWctCgqOjI91+jKgEr1gZJjclmoWc5
OuKWge0JcAO5BGQveUGhnivTQ5IPlA4A2ZKsRdSr8puNbrvDB5PUiHYZjF3XSoTs1+o62cLUXWIq
DYVPYJqQeMoLq6zsM0gWv3jnE+gvoufrDk6Qv8NYXHiQmmyHQFb1rfS275cuGDm7m8lZ8DWzidXf
Nrnfc5I0xEjQojA/0hBoxkwbTuv+oKiOYG9iYNWMYyex1HB5hR0Vs0K9Cm7Bsawmvm0c7uA9z+sx
VBJdm03Sxg1LVV6TDBR9BC3MI8qIMiwNH6xE0BRwwJ1oswnS1fwNjI+syz2Ayba2IJxAvj0i2zu1
2VlxjgM1DXGwBxyFFvjfHJCyT0nQ597rz6YmopT8rWerbGjfY/n/Wy4gFYAmvRg180rvaG2sqdhi
JXe7KBXgEshGY/M8te03aBSL1gWysUvPKh+YJkGw6A9p9yh7k/L8IBxDksmvqXZvNzY7ykPzUXA9
ujBt6ie7Hilzk5xTPTfsdlMmi/4LQSBNTozzuK5kGPhXQC22WE/vUnHWTtjnIB9T2sIRQSy/gREH
hhq9b9eB10oI2DTtjTGxh0zLn01msWrd8mySN6u+HDP4yY3XBcJ4IXX5fcx2OhNFDLE/9w0fPGtm
/tf0ni0MxLsNpiea0aXwt0YZZOPbNb0KPFXO/0HV5jJVjLxGyrGhPQsgbsvyftxY3qoyke8eIEjI
XCNQ4BBG5VDG6ckdpw9SNyd2RzkAFuY1bO/PhQsy+HFnS1zKh+Tt6Ax1HKBDlo7Y0G3veu75vPE9
/CQueyAZz8W43Kz0PHKxTuktvPfr9nNhzTPZuDtacOTi9eLH/0Z5j3z1MmbsC+wi4X/OL/yBbZIr
vtY3BEpIk45pGTrV0HWj5+k78idJxVbsctvufU1CScbSwE+8lg7hoH8ggywqNcgUl/+fBY9ObNbj
xoJwuXsWQLqE/MfDqbFe4H2okw6HOZWC02wFslLiLGXXWmgthqjHGl2qv84ej62hnjGehZf2wnQC
weR6T7U+CSjBoVanwi3yOe5wlYDRYUobHr8J68u2YEQljxlvuQAlQ8xRVnzAgiTailjEre/r0QKM
sIeXJhPMmCqSxuN15pjz3mT30B6zFYutf31CrUJWMRVnIKyKQvFs99alooXNpDJccmhh5vv5RwqR
x/QzPfr+tqlyicVB1tQcbRB+xjRWpJY+Xj7qF9X+zMc0dwsuifhNILn9Gv7d1ddRVf7iKTHmLdHw
oVlTfrJWTkRZ4ESZoHbeGibX0sv739xQ1AN2cJQ43HlwW2uobFOYnFgg7kbDmTL+tNSL+p+b0pEY
TvgwYTAedbswxo9To8HtJM84KpM4IVw+kuTmPAKbbPZk4ZT8qEpyfSd0KjfeJ1nDJ+xWKA7AXqTF
gEDXrFX+pyFEQTSeXQV5HIkb5C0k7ickqfEsPEG84Ih75+20QrZb7DNyZ2MeSW+kifoqxN/NCCwZ
R0wX4oZ5LjUDi62cexSFFG9qVM8J1EOOBYx6y8qmi8UCAeXtow13smHMHEywNWOdyBRni3ol46LL
GdDuLr8804KVK2hikpADq+MF4prB3G0u4pUQyKqANNvoEWQfZE7/Yd4xPNXQvhC67Z8YHvLgtR1o
H2zh9T1m7bRsmK0fTZlYBlF+dtQh+dpq4SAtkBqJRydWM4RbgRL2WAmRRtaXKofjr0qZGOQNI7jU
6nxxl8rzgVk4FJZRIcYb34DMQiV3mz2ERD2MUpgm5bbrmnIfVaA2JtNCVEmQ4CQVNWn7/IAT9Jzo
laD5x8mO6YiOhuTeYFaFJ5EAI7M5vaHPX1eK2ECOy7cPqY0KfY/cv8ga5rKQ/F41ZeOHG6eNBP2b
KfPeGEIiJxER+fL0T5ESUd7mBwazEuxhGebMrw3EEFV4/OIUvDzDoua/5MzNGrrUUW4fWe0ZUpm4
t3AWN5MZWrxGSjFZwxu5PH0K5fqGulK2tzD1k/dPZwhgUFNS1UraWOwW5KjJoB0C/n98pQiMSc/b
3ItDvGlq8mx6snQJk6XVgxDt4gtU3Bj9KOf0exljbOUhNn3OGjrtooe7XlsODGTF7gJzYCkb9V6Y
odwkKZKuSsh1WlGfVgem6xDWCK+GusRXI2HztURX/HpQLUg78Bu+cn440XyU7Ki2hVRf69OIYa0V
potpcqX05chHW+fKE9baOoN+r6AAGZSb8QJMOs9BgvoVynzwt+Jq84Ti6MBsNjWaFwYWwosEBdYT
8HTgCDPDYB2RrW4zbLJ6C25DmIv7oDOI1Z6US1ak3whSA0WA/m6CJn0UL6wO/AV6XyJKgjDvaCE5
GY28uAH1FqFOuNxYM3JqCTAW9PjlBIBPS8BhHrIU1V+WX/DxXx28XBWXs1R3hEO7X7+vIyIfxxT5
XGIYHsvYCMpMX9qbwbT719c5wHOX5QZlulzdxWWqD23GbMDQ1TfIFoWVwkw1BFKS7p/mFvz8q56O
i2j6ce+s4Ey05O3TkUaxIs46EnsIQtGlLXHbO4RQ1F6MnY767sA/P7rKZLi3Lq6usZ646UvCJyhg
elEbAKOyBoXatJnJaHbR2HhQETmR7yoSfECp6RffwAJeOGmURONfXk13W/q24llFocmj9i93qwSL
KXveQvdZtpY0iZkEhNBU3GEkVIIaTQZfT74mbYrwQKx+D41YrCAKNXjMiaOJbHaRjzIaKi6uQVDk
/DdImysP1LMvTMcMFelpSF3TiEP22YvUlT2lH4wgCNpazbjzBW977buQRkfObc47hw/JlTCkm7/h
I1pGE0P3xn3z5KZtQt8nhNsku24rTDk4GZ8dYsWAoXqyxju6jSKEIHhm1TdxV+nkqMlDIL7oVf1c
DTYdDogVXA3cITWl+T+NGAlNJYa0fSZY5ry0I4oPULwp+qkIPFwqI1FL6USv5EHtRMoJyCS4CpHw
0SIw9QTqeAjInHw4WJEMqxzp95mijPnCcnce7WmpmKtRXVnnc6rdAy36D72NFnndqa12AXuzBbis
6/exgnaX7dUDRLT6TtW2SsGhIoKvcCnz/edx4EJhfVJAoBQuHKNLouNopHWERgZuTz8fx+SVtaSH
sHjDe1sMYubFpFPSSyBzV/G9L1Q8k5XB6FUo2Ve9xaUG2/bVE0Hj4n3p0o1WSVzS9iGDZUnntxVZ
b4iRAxAKoy8dbQkl9ZqQRuSNuvSY66clyTzBbvWyMHsgkhNaKwhTj1BYybIReaqmaOgdAlRfzdwb
q3jeALIvX3ROFy/MH06XI13AIPzhDtOL3r9tKXFk4UoEPRHUK0FmnxXn89Wx0zFJczqUnbnFB7Bh
9wMgt4JJkc9JB6s/ZdHwQLkevf08WaDAmbTfIsIu3prBBKl0I4BD//WMv2bQwQNwxiSldLAbmg/+
mvxYOrnpBWsa1lP4i0/cNQHvU6zGwbc6Z9JtAD5efDODNjkqa8fVRejXYSEqlxXgX0ihjND/cqro
lHVNLZov+GzBcdcRbAaNkNxul/ee7FfeRPktVzOLdzgf34RzbQcO5/EaLKBmZSekbIGu2MJGcSMd
BlC+T3p7z4ThFhnFklg+WK5LEAfrEwOT/urO/GqcPkjR7tcReBY1zhKL4EjWE4X6pH7frVYNYloL
c08Ikrz4VdXXyQ/vV809pb0cGNbye03pLnks+NacMCTKEY61Ci5JRriaIKcBGfpzrx34BQHegypQ
kOPJ4jj5m9xsPc/robjLiSiyy1C2TvdmSoH8embp9QfoVTyukIDHFeO11X9svrfzywDUFO50dS4+
WmqxLugZv2KhAB43xH+EXxWlStVUCZJrYlTXkF1mxju7e/LJx4jO1hFJvI5ujZmDQ1LiFTNjYhon
DwGYh2ycF/qapAsApOp9XqYqUSb38o4ceWU7jQfri7jifBxmRHsGKbW8C1hGSmMvZeUTLxbIG5SQ
jPlwX0NZizqTnIZ5+oDOmQdecwN/lruXV4Hcmm/fyTu8CW4TDp27wk85cnsiQ5TBTUG/i1b230/N
BEFKkfeZXxongj63J/Wt7HcQmMgIfuYQjw+3suYMS3xFT5jdmMTZQTilRbeszNepquje8MTTxckH
+2Vor+nB40JJRaepfWb9KvQYc5cFpy05L3xy/zBWNKxdHlIRA1wKgD8r2/Th365nGIj6xzKVCzaJ
3CEzReXiYdMUX5xm8dhmAx0lYtRyD+Do1nYyXSrUIVU5f4RtWzcThTAR+0QKGvrHFgLI2cLSgKYd
0tJgq/vqSvS6/xZsT0MtkNAbuWM5TIur/4xI7qTDaVt/6rjOgtbOi43VDAvRwTSf1s6cYyn2SSSq
HmZ6K8aeDHYnmkpqJ763V8rFmzw0xCu5LUDZmu2EZ5XNFCFgfuxjBzFav/zhpZnoiAGWDGBb5c5N
QQvWx0v4fesbdbm+RGCZVDMDxTQUm3GXCaUtlqcZbUzJizPv88OHoOmoxrKcRZkuH1gSW74jnaeN
1V2EnFx4kciaa1wpKLkF52qgvCQjLjFKfPiuL4tq2C4lAMq7BZ0m9fh5UG9F0OvHe6b1gr2nk9a+
wkmi9WRQ1+H9FsemwB5+Ui3TUqm4o8TpGd2fD4D86vxFYsWZRXkYuKxOzE+vgqnHxMjw9QgaCUoW
7FTMg3TOo32il1f5fl8lYoEZTkt+S1Fg/L6OJKc2n3110etgkdWmo8Lg0HOHPtYxrMXEy7J4RI+K
fSaxdCC91LZO8uC1jtIB9SMcsg6tsXWky0OQYadBXx9J8z1ZFSAELYPFlD9ZXVrOyNcooFdSdKz8
wvKoPqMs/pB/ZbEGrQVOKZvHljkhnrkU4dmGNx0SEQMmw/64LX3AR7URr673lQepmTou+LjtEBX4
7QMWci3bffUkNE04G0XrIEKo9o62G60JZm5ae/Xy2XV7T+NNSK88/gB3wFifZy2mE71iqNV3Z9g3
cacDSoFMwNoLdHlKQg6UqOyaAE5uaFX8IhmSE0GiESSw6a53dYEI2EMRWaDD2h0Ssgj5f/GNNETT
QDfwlKVmycOTr5/2YoTWAn5xuUMbtRY5ookZmH4y/RwKHDB6wvofFRnibDklRVp6LZMwJPhXLnlh
58rQA8cjhl7Dhjcedyc647bVSPxmlayeb2hW347+QohbYktPqbQNcKFX5ItdygjkohM1vktI0VHF
6+jFYO9pWkdYotxHudrzxPLkIMuOYgACmAXu/frAF1D/LOTBCGcGDV8onMAUmvJ4wSVMG6S3vwX6
f/g0bhp8chEKpGZQ3y9A2ljcoqbpPLYKxkkM8M+oMWofWSKvQbh20O426fEZky97VCW3FcjpeYxZ
L/QhO1L+ucoM/f49P/K7JKaL9czQpj4Vb8P0pzHqBGTfwVKXmUc6VnrPHrYlBTynE5HFSVGRQ+eP
zgPAJX0vD/nzqGvjQ4xs3f083FzWfjnCGKOIiM3tobXkDCNU3wSVwYovYlwLIxtbS+RspicV5dc0
AZnrZq6XqSSki7v2d74/Skj/Z1PBOEv+5jFK/WXeCyDFmhi0xGin54yK5zYl3au+yQZMRCN101KQ
0/iO804YHaxppg4TnYlBehCy80KsKZKmGdJ3LXiJ7L6XW2NlXM2Es8hvCcLEDAVstWq/l5wLMkUn
6JsCbZNo7REDva2r+vGE3ogNaebbf8q2hJnAvb/keJZbF8KKX8F/oFJc8wf+h92ZT7zdiVxUXQ7q
4kwtfhn8M3b8W63ty4mpXPPTUJKy91Dx8ra2ZH3kZDqXSE/iqo6w+41b+r2fxIsMq8LEmuVuhCWM
1Qh8vbBlZXq1O9tSXOmmsXQMTnRT/OgLE6odbZY6LQW+To7Up2+KkdOOWD8qVDt5B5eXMYh5vjoy
8wENwgx9OvkB57SQ4yICx+bf+SNUP8htj47YyWrV5oqsO8nF3+Owid4aRirDkG5bjCOwtuY30Nsz
G3WQOHSbvzonq27quzGDpn6+bR5es4S3ubx2j+BhDxVddAtl161oOQ71WiWeHT+y3fBYFKbiaPem
eftE2BvtNzHQlOnICgZrgMK0XNL8fWnJMKric8R1pPMpFxoX9ula7TmbErnF7V5dpjRFhgnNZ0tJ
VHP/mKm3mWwhiTdSuUTkKz2dQ8Ucve4c28fYL439z5EwuZaHGRzv4fM1dqiObaQukQH3eICTD1xI
NyWhcELYy3hUJ81c+9fqI5c6GRXEDk54wmP5a+17Fkig/Mdp8FGMchD2gcnBlB1O/0fG/FvDNAYP
Ef88ObcrT9pWOLLs5HY13k6ysSjsHkW7Tmz+isFo5aTVefqFE4uJwf60Y9o63yYfTNch2I/Bp0z6
R92YGsSAEObF/0TJjJDDx91Wx3FXb0mGrNVWO1w/U+W7rj+ExBi7VJ/wB4/n5Q8+04jSdy9HNLYG
kwxXctImX1H4sT0KGwiGogcl7drBvZyW61Q1QsTgIhrkVB5x0RE+YbDn98mAUGnXbU4zzDdQYsoc
2OLaHuI2FqKdI0FrsrT2Oi2ftzIEtjXoz2H4eU7oojNgjDVOn7J9vriZZ/i3Vp6qJ/6U02+MsGNJ
EvGZ0a0om6tm6re0D2YawxSffGZZkR4tfvuV4arJ6bIjiUb3Jao2HEl1zflzDUCScYXu/9ZSm4i2
5yHYBnyeNj/yEOx9o6C3tkq75BpB1TPMr4i0Of6+W73TxA5tzLrDihzuGi8psOHu7gguqmPiJ3vk
dy7/n8b0LxKTPlCQ27z5o5sKXaOaM30yk8vRI5Rw+bjrdJQHIQSLmAFFT2JIcCLWvamKbBQIgFxD
d16AOs6pTGQK+Qe58vIoxTezUgHBVfWjbrEVMQtBtSaev20Sz+45HQUbaeeqsR067Pd9deqLuiz5
2gynZNqcnHvjFX94O2F3BRgbZ9Ueep+0u+0qsYUdytqmbBxFoR+3c+a+TKTY9oB20osid+Zh+bIo
6WbZb2DcUM6jjgOLZN2vOA86sCio29pHpVsBl2Y72YtKdbkjNMn1UleGGpXp1xjtBigJlR7LX2lM
qAgYwDMI5gYoGGJ4jVG3FbynVe6vjPh6q7GYW30NfuLJouYmYiZyoK1G3HQ7HczvLNH/LFSE6z+O
310q8CF4+BIZ3Ts6AoHb9X6MM6cXD9rq/hYsbZEjpE8vxJaog6jL5dSAkhLjcTy/HIDUbkPVGJ/q
Vapa5eouANx9cnWCtmfkOKt8vg70xCemNfeqfSo7SChnS0Ckoo+uxXh/otlRFUoYPVFFO9RYcES0
NlaRTL6T/wUgJsdJNOWPm9qWeuFdHg3cK3hXVxbH6MDnct3ooMwdMQ/FdX+W6S2DERwBDpHTyPJU
tHMvTv35qjOfiBz/SKCsgss9kbpmIGlIg0gABSjwb1e511vHYExtIqFO+gHAoEZ+rhluM9g8Ix/I
GSCZjc9ntMw2J3V9ibx873j+pTQqFplW82m3BV/fiJlbWIN2EPgw9v8FT5Dv/cG3tdkAMHC30CSI
lU5PG1gQ9vDSPgjCBmcnxpd6eMeE5nEJTuteVrprVZDe3AR1M7ZJgId0WlEp4daLTqFpphukCawq
zngkHi9F56LjgfUIa8P+5RksQGFoaDAt8+0FBkXW90RjK9abS95TOCfnvvSSOPEremO+6aTxHQ1b
mPcAJp2m2ByanMYF+6l4z7cfFNr8aOSfxeMHVu2z2V305F7ezoHPq5qnZCnpiLWCiD9rD0GksSje
8+8DURw7t0UK+CMPga5lSHXON0uAIxdsUtq+fjXnM6c8h2+DpR8gIYGoq3qDaqemApzZTg7IQ19D
/aOhkXDdjXE27Qok8/VA0XpikpwCTZbvQJorC4etrLI/R4zBSFfIwNsklsBgqc7ZT5DjUDpahBJo
V6nmKzpJTVlg6T7xHjvXrcWa6bAVZUhrulR/uWbuzyKmyPEsVMnViD78PlYfIEHU6DLix34aeZp3
ba58Z8ha3cKr6DpO1830zLHS7hM2AoqQCR1axffo5d2nvMlMxKGrOkl0ro5wglI8bxtMyQA1yfaU
/CaGPoS5V2RMAlXX1JGU+WLRFmmEfLRSGlharFjsiQ6MIr6Nj4X1tTje7cMpCCCmsfwL0TVTKTKh
HWWVe/CW+GqN/U7vvzJPszIwrIPecr9e+K8YLhiTZ9kEWjYvn9nZaMRLiJYGoIt8zD0L6c0WRZ+0
bTt6DbGUayH0gYtfuUDyl6xX4DJUM1RFjcpjavXT1GaCf2NY0p4TGK/69ICG9fSq3Eb7oOY0HHe2
MCKlRU5+ku0NlPYZ7TP4Es+8Xwhh0D0WkGJPXlWJDRPUkV2nE+Xzm6HrAF9TMTSGhe3b4Pqy1A10
Q0HT5/QAi90+7dvjBWQDvV7NrAQyGG/mLhYmWSknfPet1HY6VxUY0uKDZhJ6XzScF0xbXxb+rWEn
EYHFNXOga33fvBM5hsfGZsNGcWPQyO3B0kzlCdFJnJ00u2R4YHjvBtfY02lEJdTIu5g0ud9Ejdbo
+mlRfa58/Heqmr1F0qOQxv9FdeiUR0t0DRqVVV2DEmj/xjseclpQGkKkjdmoTI9wsUZOBTCdQpGf
BQ4pjz3xgUqStygoanSUMwKpqmYH2JEW6PbLgZWya3stEbNL0E+Xv1/edP2K85RPplbv0WZAsHDS
6h4/LqfC5WcRSBBB7Ql2jxDNdmKonBltWkGr28C641MHa9pSbjxTOm7zn2uG7IntFWy8VagIZJDy
izoAHhtSu4j3yfImpjOzwJxfChqw+WROILK/4Wj9stVTpUO3j9xLULF2VilLpV8DCF81YWvm3/oF
wUUOGGUhj0VI6WKdSzw5yjXiEV1uPoBQFCqJK1ZGm/+kum302ze8fPBA02iKbAyA3nxIBwTRm6q4
q3hELOxSP/fJ1XOKG7NzaM/Cvs5ohQpfj1sqTQ1kb9XQmV2PTESQbCzcMa8O0K1cVlBo4Ky4zTna
qHIbVpurO+IcrhKxUmwidRgOcs7wQASGPMLo30eOJiztvQZT5vgfcB+wsI21wZd8F+yv32VhUBS9
qycWm0fNjsPHDbYjylvIE4+IHXuxDo7KSzba7IMao7MFnkUZP971LFqT08szBMhx1W30wUiqem4P
K4hMnOx/qp+TgCd/pmAzMyOmCVhYB195qU1DVdk9easLfL5pIFUHW++C9VBBKQXzRy4nS9Vb17zh
VEHIUUnrrKEuyCKc8GGVLzc9kS5tnRnAGugEj98qEWhkzEvqf3T0bsMbFCypTV45fzjx9cNBS8/W
c6etTMjkGnyRGcMHlx10gKIb3l5YPxzhgdtLY1Lde9HGF4EoS0hq9DNKguieBxvpApaE3NqVINIf
TiyV5Kw75D//rre7QNkcb9kJfcIy17tXI0XYiWGjnf2LwM4mYzkZljvKgfvJqx5T4xOs0MeQ/+Y7
ARRNzoHfzLL3333O2tn8lWVIhZbuIJ5EE8zhdhRcTBYt1yO5pOVSILVy2TYDpU5N00eV10XlGMLf
+e+2jpTVGS5IqwFlDMo76w7E2DBPWlCgPpmtKbsjy/4lnH7JK8+o+BQvUVNGgtF9ss0vZYgRYKSW
evR6QjXAfgyl9vHzY4U3SfWU1kU6XVcQ1EzgJ63Ho1OaozNi5YqNgRSYinp7iZyrg6DtpqJlsTIH
7Z+FJ9NzPYmWF4zyab/rEpDfNraJMuPh8gxleLQ1m3CK96DZ0GGECJuFpuI1fwZHXkkAyS4oslR2
FG4AzrIKpmMU5LiJ0Ttc7P3Vc8hhsubRjnWPB6GqkCaDdQ6391AO1n5fkE+xFZTU7Py9yWQ8RSNv
h89GyY0KSab23Kqldtjh5MUkeYCEQPZpJWH6PuHrhiRNWuKgteyu2WqAEK4jNOmZ7wdXuksYhT2Q
xh4EJtwLKc19tJVA2CpB+5lUBw3gk1CHT+L+MZFhzd1kP+/5VROdhIcr4kelITkBJGTW8lT5R+8p
y/pYjgjpBqUgssQiEEKfcBrOSL8itY0SBh9gK6NtvpmcIKYeFPbOTQhU/P528ZYoX/M01m8db8EO
OrSY5nI+na24yDby1AYGnKX2icgA1Mf5dTluaSY+k9rwATyuwOA/ER/hMiJK+NZ4pae4H8TTqOzV
1ImQf4dwRA7aEp6c+XiQnFeuvq0X8j/nFBhTBMMqJ92k59W31A5miIXdhKG/4K5rcCDAzJsNzpOD
jfWAEgKsi/26SkwwINJ4bZl0dZ5ory3LPoeli62hyISKI2S5TIlOgEwkwf3qyU+4Yzlb4a+IrmUQ
0zeE0YAIY/mf60/Rd8n8hFL5CpxH79qeA+KfjjAQVwKmq/ZIEAcnYmj0JtnSsI+c5jceXiQ2IGWZ
Sgud6H0hd+gHXwHSm2B4UwgFXeyBaIc3FDna2WIi2daF20IfVlS5iGl7Rhs3KND1cG+txny0TiRl
UZG4t0Jk1UzflDDnBj6D+SIAdEeZOdF19FTphUUwfo2tfwbjAOH17G9HiCW0R/usW1Y+i2Ss1g1c
+FlmXaHUoPWGzBKx/ipi1S6ziLEW2Abwv6mV9nctl6o2AMRCuP//qWiFT9QzojBbzOgOMrzAO7sO
NbxfASg4PKr60GOu3zZrROnBACHopr0JC8QBwri4u56KvIG360bWvxDBSWeeRIOovis5j2rsjEyd
Oi5735532Hw6ZzjugVvdgMAJk3cbhyFMQ/tSCaymRi1njjQBAKMmnziJJC8Q/0p2TX5oWdRRKa4W
G0rQcJhwUPn5nVBMAjbUv9olLCDZ4V15q9IejrA/yDywsMiSvYyOyDW+tMsdPQsIrPfTFFuDpQ+2
2R+8MCIE3QyTo0pq9yM2nNMUheqhoxCjPgJJSaHeMN0tUdirnBSNgczpHMzB1SELPDgZWUwVCKaS
CW6gIglb+Cv460SQtViVnlSCRXcFKUvaql1csyQiOY6bJvKg8lIZUUg6X60sSTRewBLGiuVQ95fz
FGP1YrTNAldu8gQtaecX0JOCc0ZLCaaJmnbJezU6otITV1a9UXuv5n339alu7ADTbB0oFBJ2KaTd
kR3rCe84PIsc4bQCLOOvG+vbCn/SOnzXOEDbQjx3OhszwWPSujoF9tu47/0U2/Bb+Eyh8pvf7K+x
PjsCG7EM6O3U9H3AQhf5hptOVMD2OWkI4h84/oZgGgyNQzC2W9RCbz8tJQ8KfgTZvrsX9aA45U1Y
gb/FAImHo4qrHeRHo8Bjl/YL39z18Q6a4dSB+42wa0MTNvckQnxnAtVLjuyzj03W1tkZzjmQW3Ca
p/NPczUBTS+SirDuTepjRWG1gXxc64NQSQeiDsTIkZgrjrLtuHtLeXf8wuJ7rk42/URdxorjUw4r
7pOze8bsWdUxTOg8/ommAmFumenEjE0YQbX7PjZv6Mrn9OLrC0EgkZWCIKqUArTL6ppFkfUQIjbj
JpDDAAHorT6eu6iCJzxdUu4hmkKMDDLz1T/gvKZTR0rDEQzfLRYUJiMzIZEB3t0izhzNz3CzDyy5
KVDU8j4RLqotYbd6hb6xf6hAFRK4aTVm5povg8LDrOddXFbivZhT+e3Vy1LSIU+aCgaomw4YdBFu
m9VmgvwV4PFIrYOY166cJWohXv+6a8cjn4xhicaB24k4Phs76tu3Vf40KFlGbePichbjJMt2jn7i
fef5szKbRTjEpOcW2g/Pjg7MN9ovGyYWIGnQ3DdwlkEnc5cWUlV3BGpsMdzxw04kflVCtjFj6871
ZXmvi6SZCvjPCZXlwBrRhakpOqliUO8uhcFHrbGkRKfQBQgPby6Gks/QSJ8bL7fUCgsUUQxg5SN9
NzUdSDh4MC86lK/ZFFQGdSa4LYBHjuMp0UayoFb8mgKp3MjLr4NUlzWTigL4G86mIKZa8Ka/S0fb
1ofih3+SI12i08GlDWA7tgoqJy3htBi8OwvU9gec03zRUu8h8l0Wgrmu+d5cpCiSCrtW5t3PayE3
0RALxNpjGJy0R0KWwWTeqXrwzkETsmngJr0R+nJ/sURRCDiGOEfa5xyDuEQtV70zQWQdZyEnsDpu
8Q+sK9MUuosrzwEMfe/xUIotOCJRfJ/iUpc9rr839EKTaUykGsllvb53JW/dwffPbFKRHdsMrIlo
M9x1SLCOEu0fvbUQW7dDv+zeiuutTUC+DPzvKUZeO/lU+1zUhLtxoOOpRiKne2FPyWf5sJUH3tyl
2mw+Uc9xRQ+yPesYkcwitjMkMTjvcvaB8cYA/8RCPjVrkU7nRGTUwMHfDd3rKN8pc0vKcykzd+z+
fG7fLdn2xZ1n6y5NXYWN9OVxMozCh5IEGAsUvdDhIV/8MQB4AbTrbcQ6aI5ijWirNcIIvYdV84K2
twNb1X69BSNyygzs3fSAIAfIZCH4gCVy6J8FuCZO+pkoPo6EIGRm8RwLnQ/xvCNjcSHzGX80LPVZ
W4U382HG2+zc9i+n+WN1UuAosrzCOA94aPDI1V9FeCrjtyAQwMKriOfU3NYOZxMjEVJZwRdSYhVW
0Gj0VIjKYI4qsv/CW86mj7VNXR9sO4m5cw6u5XbVq9HXcv0oSWmZROe1ssX3t0ub3vlnYbKdy40D
yO5dbvWdMF9wdUP556tTuMWyBULuR2Igm7887EzOi9RUEum6h8dEc4t37hEF754QmF447Unew6dx
yEs85QPW7R5GLLooJbeEvw1IgHay4Gmxn0uxejDcTnh9E5+ECbV3JkKazazFgOI9rVuaShc2su/e
VagctZjjwU26ub7BuZJNJytB0a1yEVPKFlXGkcc1/TE5F+jJHwFx1T8Qm9Eox/gwv9GRbltBUB9x
rUWLXgPqKDtAFMSpkjIbj4HoYgCiXZPaB67rvhAGu0lNWTc5+msWBIch7h8FgAjva7lrIuVz7oe0
z/GNMTfPB8e5Vuuj0xpMZjq7+uIRxjL+BNBOb3Fh1jKSrhd5LMmyip6KbdLOSiLylAYG650hm9z2
eDsRglZNhPUWzTA6wK9Q3JyXzuyOZJ5N1tBx0v72k40vczg0Jz7yP0K0VLaeGEbqtANhMsCxCc6x
rXtKeEoPWEPkABf0K2i8abVw/+oN9h93C7zYpKTfpS9jc3RzG3Z4AiBlUlz+lNLKGZ94BsqApRVo
v3uyjkVQ9KGtxRndfIzZDCfdT4OTkJICDe25F0Cc48JumrkRnSIO9uBHDu0hpXM/WUOWUej8w/Hv
RKlrVAUVpukE8Unyy7QS/EmtRP4gKS6yarHu0A5Io4rluv+nCisKhE4tNVhEnGMgM1PmUNaR4d+n
UQLpbFXsJgG+j0xDjdwkDJatbf/5Z20pFFLndr4vXaT7rLwtN5o1v+YgVBW4UPe/fUdejfAgDXoD
8VHcWFbtkiGtagoN+NkXmtzh22aTVV5PVH3lQiU1wC8EVjpv3SATOqgs/Bk5efiijLmGjdxlIESl
buxFyTWqEBf4GphJ1zJ9LuJqqyg8zk/rV9eYiPepHPymce1vwtFxuMfRZSwFQtSAflhoaFK/1Ui3
fIMAyL/g43LAYAk2vsm8rW7+LiW1wqKE81KzSD2LxYM3zdgFG+HHC+FLAH+mYgmqok5ediLDy+29
BGMYUTUgbd5xs4h77UmC0Hqq2Typnaqn/wnlGfHDd9zvtDiA8f+4G4rPE101btulg2yqJKxhfFIh
Q6hgsDOmCO1ZUkeeZG6AFCttBWby2bDobmbs540WR0IpIv28fZq4jSJJgYmmFWXFiAUXl6W7xq0/
s4X80ahxaUu75jgJ708sqL3nMjVNxAhj6Fcl5/eVIliAb2sNdxnl2Da1mQNpvRvp95qrXA5/R7Pt
exIYqEsSOmW+0Q2NrvP/v74aEHJ8A1suhS7DTkTlL3QCw/ryiFU+0uTZePZXf+9oTHj65LG6gZux
E3XqVn7tsjLtukJerYCKZeV1oRFnrhbktfFF8SOlVxZ+/sGSi4gIgWQsDMKL9+fKhvrWWKcy10QQ
PXJP9PM6ugmA2lNG6EvBCa5cUf7IipTc6itnIDFyCznrKo2YR3OllFZHI4sAMEsKWmvcLw864BT6
M7MOYr9zU9HRSSwUrCo01kD/7iAgya9DDfWhkZ29YokdSTqScJo+lc2E8B/RcUJKUC25/V+OuYaW
LuGz1WDAD7lB3dzJvfIcKU5Eu5pfxYMuS5bGTvLYg39MzA5QNYPvTsGQWyNCAwcSwwwR4D9i+sbn
XIgPFrQ579mbCjRFrz7Ckx5kKg1mrrn2HHSkzILuH3BX/sN5w6bQATCcRH2xiEt+4JzHdyd3tIRD
DcZVcxCadem9GXKCzJRoZqBdDphMuNzrSvNms+/WRLoq+/8VFD52Z17bu31HT8mmGBAU6WXa24Vn
dQeliWnckwHzyW4T8BrI9V5odroMQRINa3AWRlFmeYczfSnun5nqwbxLEDwpvMgb5lAj9XknJntz
4YlYhVtaElcCKiTmWnGYlKmQb+3Fx0Oxv2/eGubzx1mCFfKWJI94uQNGmTdeqAGBzUZJTgbGSto9
DWi8/+nu9bLVNq9f1X9NRW/PThBDDajBv6NsGZLYItFlT/OzLhzYnfxIJ0jQErNWq56k2ZyZIMFd
LbCuOU1fgmI9op6MSWRUKfEBpbdi6dBdmTV5bdQnSU9TpyTG1oTSWxPl2U34k0p/S4aMLQ7MToum
S7OWIBgvAQNTZh8hR+T87xkKsTwM+IZ2TcJgkFYxVvrIKZHD6dFFfWpo1O9j4zyIO+d9s+hfNDs7
G7Fx1/BmQ93LpLjk6AVGUlXMZRXwzjNVO09EW0SmhUwFqpwlRd43LlkipdpB65s1xrFh1uaeaWt+
Ac04qY4xWKTDZIxRvQVd7M11EsxrLtHxjYYlIDtfUbCYirrNtujlOm6/b+qRluavDF3+y3zpKWEx
cEu0VTCTP3LubeA3xk6FhEACkOjeKAZEDD0sl29+ZKkglTLZiM3i+ZR2AE9uo227uNTkQlQJnpBY
1m51avPFGx1P24OpRTI8C5zVLB/nWPGbpmIeCF3HvY4hDDHUSDqh34GxXk8VGnuD4ZjRTUH5QZMq
f/zj1AQTyHXO86wrwuxFHaAlxcwLsOxsCNmfiWPWGquW3tcv8sU4voOlo58QSabTe0+81ygktfS1
FOBtndZ50RhHERTlOJ5peVGWwLaM45jlp5JCGSapYPBgU8h9qH75ej1eC83KpPkPvbOlowB+5GX/
UnoaLYhbzzhdEuyeGvJ7miHeuJq/rONlDbbZpmtT06GlFk05L5NrVpUZDx8RO24aAaKbJsoHbufG
ZTOVkPbs2ToyinT9cJwTZaa0zuLBUU0k2g/pEI295SzA80Ehee4UihoSxIQeF4R73oNzNsa7LqWy
8+TyidNob4E2uzgZs7MUw4gBQVBBRMU8wrxwAfa1u0G49CqjYReobAh5oH+mPCqa//ktdIRQcOae
5OuNTLqLKbjx+9dW7irbc5hqN5tM/Ud+qCg7Tyfo0PqtapsiVLkTkOwiBBu7DrskGpxVixeU9ZdC
F7YZgMImuckareSjE2CE+3EEBceSQDLlTzh9qiyCZk1fmzuzzELTJ04L3UCO3nTx0K4RkfW1X4DY
AjuVdUCvNjE8CKfxkxlCHBPQhVa2/MaBh0wN/vqzEg76N9MQ1S9vHWOjLHbu34lsLE1f4q9Lq57p
XMxG6qXoxlme30Sq+A6VDN+Z9Ak4g5JG/8X2PeJVLQHrRs7sIKPxRoIaJIk3MPSxMrrFdNVeaAhd
l2wJT3nz/vfdKrPY7TJTLl2fawQdqZj3KILVvcsSQ4vYWRQZ8TCcAhd1b7UQxOvOs33btmvyxj1n
oJmyVpM16epXWszBU/bEJNCDngSEMtIrl7JvzOtuRIyeTSP+8JXg4SbNqXdfDDSiv3xzfq+d2wpA
tf5RB20ossvbsPhVEs7Q3tE7W6eeZmibCGb3biGrqwYOkh4Sp55M6vktClFM9ZBYueuoXqeEmLS/
naYdrdSTaPv3nR/zttm8wN+CUBbIIGcJSrGnARF/ceEeC+HMQRg+K2b9ExzXUhs6ZjlDZjeMmykc
L95DteupjfkZualWe/qsEI1vdjjb+fbxVEw5YXCqUgHFRjVI4x1+qDEZCPuZuu1qbXWL0cc3OmiR
r0neS38RwB2rT7bB2+FXG1sdgiNQedH2c4oAaAEAEM9eDVDgaSAkdSKWNRL7ooH7r5cO6NOn4lgt
/lZCm5jGGWK4uSflRgSy68hEX/y2dsXzU4/Z+4e4rblCbytYYeR5K3EQudCo0ktd2eAWCq2lkGk2
N0czSD+fSPxyMqnPO/E35sz5yG66Ksxf9UiCyUKOmvC+I8vi8vbbB13E9IXBHpMFQI4Z3qH463Jj
gWPv3/9mVM3T4vK/JH43WWO8vXB5mJ3vjTdhAsxvOyY73uRGEJ3w9HJ7cNwmpAgQKlEPd68RSCKH
a5aK3DVIjuZ/tPO9pWKGldIL5iOYUGxAR6chrlmm8PXIryfg6bmes7NNecusxzZQfyHCrikGu4ag
qoyzRBkSSMS/qHWk7raAoM91nTjq2ivKmLPJwEKRNNzcQjA4Ke4gK76DtkPnf7R8S7hXsnVFvAJt
vdxVyiAV324sKNHOxXQ4lgW7VJnHEBeijdte3l6HcYqzETEEWn2hTFXGYK6Zhv/BSj2+dq/OwJUu
YMpLfytAglNMrEaOp6wXCLY3jDVSP1s2v7ADqRObD+VbRT1bBlvz1ZLktwUfWxHOazA7DcgrtWtc
LjxxBfBfU2J+PLyfubE4NmddweXhRNfa+U3hPvFKLH/SbdZAhrmD5WyQTFJyGlMA9wPFxAhkqksS
UYwSCIn0smqgILWLBvBd+gmaitM1k36EBBObxce2u3V7OYUu12tbJYvoaxfy7sJ7XrEQwrHidjod
cjezTecH7Dvc7wkZt8OxQgHUqf6gfxsyPqNuYdRZ4rqeiQn2WORQBbpoj+aYRTOA+SZVIXBbL6FC
oQMdwxw6+ZmLy2kQICjgCAti6jRFLEnVzSM9NCTQtOCZHkcJKCzqys1LIu0HrpxKJOPC2MkPS4rY
g+P4w0Ti1I55R3sNTc4St3l6xHsTsot/EQFtACoYIEZ8VVWUW281L8s5IXrrObiaBrbeUTZ+ex1s
0OwojXeubmwgGL5R/kVR3UouQVyW6WrCF5y49r5ymQq/+ncLLpqvx8u2viFiTcEixfR6UIgP7Pri
pjtt5Qme1hkn0TUpA7wVJ7CwKzaIj0G8NyhFYlSIZO8t5vhl5RelmcQsWW+FFcC2432F2igVdwFP
zccJLmXdw56MAvppjeudG5NlPOOzA+TA89kUtCwif2RVx5eC0dRM6kh85iqBvlpjsPAH2HJtiprw
rdZ6XoRIs6jf7C8HrNa04by+pkcojzw6Ism4/7AsDRB7KCKjAEBqzJMy3NP/8JGiRA5F6NLomNLy
x2dnX73nP9v5+rKiEZskMh4gh0TG8g1o3OG4I9DrHSdqD85r816nQ1owN7G5L+RNpfWPt/frBuh5
Z/zFUv30qKIcXAKpIGh7M7WnQzLQr54EMjCdpTcMR2hWa0ld1otCgcwH/CRQOL8UraYEFmgQzk6v
88bFVvdx87cT01HCytkaoNFvfsh0YjOglgLiN6JKiwjQAReOUTlhfMoRAynjPBw411/D6b7wixUn
/rigXmsRBvfZugeGWEoHRihI81v5FvsTp4a1l5XdaKSScjZs7nyY2v2M0bKfq0/x1+5RfZVgw/YO
G0W9R6zhjQsbVDslUPekF3WZq/Bhc3Y3bjNbXPFZAx7EP9TDVkxAW8Kdm+RtlBW4BHLvA9K07FRt
jbvayaJNDfUeTYqRj5b8zY5khvU7tDT1hyErJqC1JfhaOnYmaU6KnV5b1YN1NwlwIEGTMgQJL0Ad
tsPBuyL5zWrNGfid1QvXuBbY+K14SnmEeL1KxN6xUCq9jZGdX6odvwR3Py2dDPcKws8Ze+nL/SaO
FE2nh4bLQetCQL+H5VXs5eljlT4d6HqXObFDzXaoHLR8uQCbqJfVczb7Jl02TOKelvRb6YS28dRc
H+R0XXzjA2KDhcnSCkCL7Otkz5OftOww20O/sz9weoSX6p7t0VXCA8PgJL7Q9SwXUbA9EF3yQhPT
zHeTzTO290LOGQYy50CZzu958/uUWWKLOCEVZVbOMyvSUOIIAanPQRNJc3IVbQCYfaIhrLWwHsPd
/lPLYF/v2e1HQFzjXpSgjqgEcSMGrZPRPPgFQsna+nN2oRkiATBXaUbIgsYtKDqTJ7UzGkYOKchj
ExT0N83YJzbQb8JiZV6DegqYJMDiNICPcll9frvYPyGr+iqiki/NH7HW5jJ8fH90/yy/AOX0p/uI
BLsJSKrd3N7oy7n614tECxvkvsu7usKaFfl0YOqXkL6tl6do1ohZsZneMAbSlLzm1cOoqZEX7Woo
7eqZ1sgvwR+WZfcK9V2WQHFfTQ6nZ653hTY+zHqWWzmE53CsDpdihN6aEA2u+eje+02HzmQ5zjQA
KwU2WLci/m2gBet7UPsyQycNkSwjcNy5XVALbu0TrobTRd8b2gywGBoFmPcyyzyS7eu2cZ3dj/ia
TMMFyDaul58FldBoSRsCzVRe23+02RMajmHcOhlAnk8YQKenUruZVpqNWp71d1tCdxLQOyucrKTi
NM+spGuyrcb4w4gKPkmDuMB2lg0GDf0au4reQL1esFkWfpnIyzRri19pb+RqvYVBIEsweU7Dg3fI
nf+eISu2pTYHajiBPm+rb9M2KjWivnZqnJ/2Cb6Yck8Nv1shh9bxxpXlzlOL6aRbYaeG5YhKAsQp
Ak7dKGmdTH6oCn89WRyVj/zzv8gln5G7BX3raN3u+aKtA5vQvh/B0mv1T+15VlKKt0OO0WOUt3HO
8shE97/bxNb6XM+1xX4YMjb9NPyM7YA4SE7uTme+vIzhqrdBwrxaxzlIZvQ//J3X4E8Px5bv7TqA
UQ3R886tTWPdJnLhtL19179jhZFyMTo51CEKe6Wn/KlbuWdPWPgEeSugyoIMq3joF2ymeOs7l3x7
seYEGd5wsK76TdwWfZPrTD75bk60AZdZwPiQ5Jn5X5rM9R5okctabUwKh+pw5LsB5n7RymbNvLcC
7H2UcOjg7gilKQ1uvhfLZPgleCWXf4dzkooGemM+PBQq1QFJOZgg6OiQe5GvPWDypWy977Mihg/I
nC59Zh+lYseDJNWab4bx0jfGgRovYnZFp55DZghVkNInv+SSa+zm3cX3cYZh54NdmTJXQvBBt4GO
yKmFupmed8gKzXKwx83nCRlur/MJCHq48BjexIMGDrNt9TBZtQN5R9GcoYyTFHsli03Nh99KuFMS
1dAdlqJh4S5sWwzoEFGyXwl/VCqnodpAMxQ04n/yYpkGBKG+BqFARPGZGVkgg5jB5NtHBflLGSEC
ZYIn02SvCHCqRBsDeyor6yl2UKWZJ1lVhe/DfKabPaGk93Psouq44eP9qRcpmz5YeH1JeFH6568G
lqVfb1KwkPkyHWi62VIoJ7VcmMsgDO/HwcIYb71mpUmHLpEEfyTHyeOhazjsEbcL0z6r0s7I5z5t
z1hvLKzGGIjcMIQ+QeMnVwjYwxYM1xFC8ZH7f4a8v3OIZa0xsNWLmss/1nspGbCZBCC1FVw3ZWEr
AtexdiKCOta5flfJXz4g3RjU3eAnEWBhiB68jAbT+GCkZ00C2VFgmXOx6WT4XV467ZqD+OOAZaMI
sAu+tbco/o5lrtfm7qdHLlAZgImhNxDNXJYgrV8E6W/jW3bh5cOJKNLqhUC7AtWHPemwOhar2GlC
14WasFjiWNB8JMLthTBSqHFcFImgp7ZbO7YhV5gPRzYmGpBkA6jby3xiUH79t6OVHTy1HUZN2Fyp
vv8JONoMzTx/IBYagBhL8ofAuT0pBG1aTLdul0cDbMQO158OzQRcikVOwkbHdpEmZYhSd8GqMs4z
m7pR0fEP9xB4wDwQy5d/RgNZ/Kz7tQ2NbnXi0BgOSiE4hav86v8lJm8nvMPsPEkumy931WRq+zEl
pMdyKnycifKL0I2t2AlIcDvkI9+vuaApmTP9PQibhRBJ3ds4eQ875TIHPdQG2+O7HMcTYaDe5NYu
c0uvf/K5uCrNgWOoZMgVVr4k49FzAuX1xWSFFZk+znaF3FzBCruJ1OknqwOVWF83VTGB6CVO7NZH
xzOgbTxlT4N0BkkWxxTt1b7jSskrMdO4nhg+R/9yQzYRV6bxDFvRSAbH6kXImTpJ9RTVzPD6QGdi
s/1Z3Yoj7eZ7p/hREW62Ix/xcBjfy5MjlxngNYmjcD8k/7TSGzmSRvYucp5HhWNIAd2avrG03adS
FIz8l6LHOk/nsZy11gyevI4WuZ0BtfwexiS/OBCnWf6uIwxuMrXY1zaGe6ietQaBF8f+sqvv1hQX
w5qaYP8UoAqcgocBBAK2juN/zL7K3GuBmNr8EUIZlr4SQ7eFzXJGCEFEF8FoqGruXGCA5h+s/jqp
DBKqvF+9/2ARXCSe++796qyb1r4dpJbvK82utKgjNKmDCTD3ptlFN+pVNjUIAvMayB3NOfUH7NyM
cLqg66A2BIpxIZBL4U+IhpOvxIvJD2OEiMvxEAcKEuEQFdMfq0cQfhGIlz2AI7BslwB9n4G2z7PR
YazFmhRwV4+47pYcyVRwOTXjyw8QwGylc7uSckG7ltpzcoiaK+U7ibBEp45dbNgrB5JFIRIwzXxF
LpF9TZQq7dZwqpVOGua3mTVBIJeBGIDtbCLfgMIIL1BmI+ZPmqDebhmSby7kTNV2zYBQt1yLajfu
cHy/KhFoWBL+9vsnHjehLtMm+yp40vESDcpD4GNYWkzdTGOEDj66NDyAp1djqBLiyxTCDKsMLtUH
r95WjVjGDt1kcxuR7/ttjz+TfMmaGCorxeOwYT4IT8MUEDoIA8qtts9a2/l5HXx55MHofFjbKAWC
PYOxC66FxMP7A3AWlqlDr9B2kQ0ZMvEiG7qo7kTezrIgdzOJ1WLt7VI2HGTyBBkjZIkx9SI5AbYz
1GCXxuDUUKszzZYopRCDT2TxtH6HKtL7YaKSreW3AQqS9RO7cM7FyGEFFSPM2nJC3fgfKanDoLwg
RzWqdoj5PksO1A2Wk6GjWpp1azyhh4Z129tt2WiX61FZb/8VwORvJzSRKrDibDVVuOHLUUD5Yg5d
7TJZigIQyQeMI6feZfWc+Cx4OJt6ncf/z6CZt2t7hYZjS5UxIwxa8KgQth/eMiWLfDWxZWfcLqrL
BSFbAdbVqQCZNaTrVrX3t+ajO1UFc9XFHtNUZ4R0fP+jgyxOqQgxjfpBi+qz4aSlwgrQjz+dEEeD
jyu7w/BHAAoKQergThPsgViHaIQswmTm1iu5RaDIMhhnt9FyMPGZACMYHheugkYhgN9gsn+A8H/z
hLUgGzNTI0OJkgYrSygLtFpCeZY01AN0omgVbFVXESv7e4/Emv5ds7ixGgcJoXS87cSNR8TnSUyM
Jtn0vMhDRs0Trm9hJXOHUxPX4U+189dtptoSsG8P/gOOVsntZeiA0AQauKZQKwJYhzmxZI0fjoGG
sCfwd4GldG8vbwiSLbKyd6v9HF+xJ14D/RzLHJRR81tWHsLS1ai9RCUjV601ikux67F68CFwJ+x+
t/46hy2QDc7DExAj5BCIJPNI6HOPt/y5vqOs0jvUBdMUDv9uBnLWErmOzxowbWPtaYI5M7Yv3scj
99jfBCBbfCP7DP4zhNmDYVVJ1aAE4gBPpqvtdLv9EqklbSDZl7lE3BdMDR6J34QaU6S/l7j9yRa0
WcbhAzO0fV5MUF7vc1Qk1ePcXBE4z/6TiXwOM5dJ+T7pV14RV7JsFTH4Z4wxKIA1QOiBQLkk72zV
4W3J0vcKB4AL98Bt8tYO1mSBsPJSZQK/Sm3DEbJaQdr+8HGOJB+LfnKrAFvkLkxtDJqNq28UOu3Z
4ivoS+hiOmOcGxS2muPYpKFLXqCzJBSAaphy1IB9cXcrPlBmYzt9hM0zEsl+bwpBh0A+eJE+3Tn3
Q65AS2yUMOAytDr6ahU2EX8m93QjddnNhV982IZ9stq7uIj72GjboQUHjIIrNOv2a0jDvIZQReBM
NWQsdjQjYf7QB2w4W1R0ogfVWfl8i7S+e2+70JqJdxAWh7a8PuwmTLLwyFcMpUDYJObO9zgQGspP
+ZPhsuziMO/eEfyOgpXsCDsxaolyS4n4XdGLMoI0YdCmOJ7sfg6nLa+lvxAYOgMK/IvEWfu2mbdu
eOsdljeIrWiDyFMaJi5AmcgFfUIkG8P5uxo8hUA8138XuATMsa3qxLjBlraqGcZGXV0oNuR6DInk
t30Neu0Yxi0qS3vwWnpTLZyU8sq3kMum86qCrA13oPBfR+Ip5eUyQBYUtmTgsPbHmFqavZv+Kno9
MgZ3r6ZUcBrC21vsEMzCV2lBcMCuWhWPGGaPRCOs42bXU1xuqSociqQ9YVfpieZ5bTjkgz5l5J9g
uYd4bExbT9unTdnBqJPjPk8wATNNLVaIX32KSfZ1OBWErhL6gqp91weFCMRGH8TTLJF0VghWtgtN
gLO6UeSJRP+x73eE4zMLFqhsrMgJU24S0Wamkc6jKeM93dkpBKT+PfOl3A1UIppADi0gggFjoWI6
XrSsHz6iERBU4006g6vbqhC8QBdCGIi1bQhk1bYTh728LwrhCTQJWm6PxrtQJXA3I2ZmyDlMspUn
k7RHUBpKvL6rwX6irkjCpCk9bGM3J+mTxIXSTgw2ajY3M04OgtRSX4iCWYs7s3Wop95lE91VeHsG
SKnVnB6pPa3l8ZOnGQ9b5gLcO/DqeOqoasNJoxct9RvRFe9TZ/G7QXAcpRYcXZ0Ah4l6+0j9Bv5G
H8HN4nJWGtU8ZzP4bZNIyRTQ18d0Z5dpfMizGyulhizQTqL8xrWaqBMnrVDasz50GOI4N1RpVyVv
QfBSQmYJl8F/Cj2zvjGGgqQd5zg5UHXTc/OFwJtqdT3+7tQir+LSZaOAG4nmqLHR+qoKPnN6+bbP
Prb9b6SPC0+L+R8DkBb7ErnqUK/xZyl4viVbVziCUfstSGswGnYgF84GJ3JTTveFUg4avC5iPWE8
QtbqTGQA6bEWViUb7NOzTJBhKJhKAQ52s/sJsT09gu0o0FAxyavwXXovWo3gnL2mbv5SIh02OtfV
tTf5rL7wIeGmbj/wIzsQz2LFKfdbC3RMnvpImHFW1cm0c7e0K77H/3d9eoEULNI3eW7UDwipGEKq
mvWs7XAeQxjfeMS9LyFZiFJTg7CzRyh6pBqZwswigKpHIQ7rGKidNaDmfGXs+fFoZTImtLvuP6Kh
eBqpMaRA7cEk8kQewPvrb9Qq3j27uTwx/KRlveevXjRZyELmPN746VVyyji18KiQhVA+8dEQFXXu
q3euDYs72+sk2P/A8VSwmOkYS5jtkrnjUnA8E6zKSjxogagFW933lhA2/fcnfsQnTJbYrUcefRl2
Gb0DMIdxxitqO0VI5DiKzBAKqCnvED+81E6VWCHrYJEo7wLwnGHqd2eatv6l7XtFMod7gxvXsjE9
U88KWNa5iZktzozIZiaLZqWBQ+e5hPAWlw4rEkoaGcyip+BNMxR1YQTQcLKop1Hhg3JMsZfGncw6
Kqi8ET2b42N+mi55uiT/nESdJSymfDa4G79yy4TsJfW44MCwkXF1xQJDZJoAVMx6XhmMNK5zepMw
TTqn6s1Tg+jlTp7OPS47FL0lA4+kfZrLu3LaqW+nXk3WiutAX9dWhZbobZulMMrhRL+/XGps5CbF
bR1t0Y2+nm5x0iMTWy0dIpQNhA0rklqir2XMeY9whuNsBCNhwXIofIDZB0WS9pr20eLatOqrVLTj
/kVNVZK3wtkakgxAj0iBrIka5fskPHm6A/DqZWBZJgDOlRsPMi8lL56oN9lT5l/9oljBuiwb1QAq
96YsL/WF9DiMlTUYqLc7RGWm0zNk7Z0thDBHCTFBV8FuCgIk0OqY4e807MU0z3npf9eFTJMOxkrv
NvDe7KZPdwzbwy2dhQ0fcPmQ+xYIkcG54pExdJtnbyf8wM1qvTjrpkh7GFbQPPmAfNQ1VsobPEHn
Fg0miBLHo0udQDdiLxegFPshDJqJ3XxYoFwlNJkOBjUpLP8j/o4jKLi3ZwAKDZL7y+1vm6BgYd31
ZykVUE4Cn59VieFUVjyOmVmD6KedgINXzpf2VTHXIv/K5+Xp+AQfKPmUzr6Oz4dLvVufUYNCrehH
fu6bjfiYhzfq5LL2huk2qDHr1NYHvylWjxP3U0RwHm8XxJJtY0JjaBi1PfZMqpwR3AvLY6V+8otS
E2rfJkQMq87C8xO+ap5dcLmfF1ZfIn5vjwRlYHVcImncBO+3Cjt/xNsKzS02fpXdVe3t31/84x9w
+n1miwpkVL9pQBYUikHdPXywREox2EU826QV5xqj1Odfc5KRGzSuNFjI7mGHb3/AJybjygTHTOTo
ZAg5hJLcwoHViF0FUxGrBPCoi0k8zGjSdNHuqLwIHBEzAgJ4yvQR98Hn0MgOmNO9kR/qkDVx5Qar
BHVfqChqeYxLpwf6BXf6qEynxAr3gGUZtXERLdJ9zYd/pINHUlj+s/Ymq8ujWoqZGvkUsDQxNlsf
eZj/NI9y7NYLxnaC3o+r/880+sXUnG+fcmREQhS59uEImzDyUPJxSpNfgIpso3a1ulbXjM0z4ih2
tN7/ILiQ3ae1ZorhkJ18BcoibdN9XGL4cHG6k4W1aGGTp7yOViW7sg8TSJzXV6wthFh7otnR42oa
xmmliHm3bJ33ipwaLD2dfal7yBUt+QMXWALu76ga3bqz10+Dhd8twH8sokGVbox0EUkk5T3vyuYh
vqqCkOU3fX4PPJBqPchCpLz5nhfpFtDsbKZwZ5H4rfD1p5qX9jhv03g4Vd7sRMa+z5EhFholaR0c
6uZ4CbOInGlqO02CMgDVmJQ0FZmXJkH3PE0TWskYaKxU+vVaxfCtChnquleEEQ5aZ+sxXaluZYfZ
Tq3ndsxHucERaUV1IImJWhgFsziv4qhTGS57ZrgKCG4uvjfvuzcuduroglax4F3AidPLpnsh3EkF
ozHS4m6qMxWxY4RckY/SNTuLHorkqXohuMlH0WwW+re1i5l2E98TUnP4oWubjDJVBJcKn5GkB5cH
SZxE3chdMrHRF9JGKMq4SdyaHwR1IrDWHsQ0eHnfanyJtGkI0F5MHrglopTFIZcYBQ9Z5mE5F57o
M920RfqnbrLdXYN/0E1hqdBg6LA6Dz4pPGoLAVfOrBF/E0qnYIgKDm/JtG2PotKt4bBnIZ+tfnt2
8CRVVNty7GUVfHBrsYvLzTeTWKct5DuVdpThJTb5t27P16Ztsyty4EJG6FBca/YH9obIc7GIOBiL
FaZbC6+Xs+Df6dCeb4BdKmRAQKtp+1qKcN8E6F0yUcAFREXkWmKtNAIqPhcHTdBGEJjT/D4pq/rG
Vx/iSCUd3DrdqyUwFoAsGZWX8M+I0JcscpRIUX/0HfCj9xPFO09xDFNUWDLpXmhSMDBxx+EZSvA+
Yw98fVyPPgYXbgHVNGO48mszL+POfToJlyR4TYQgJd9um1Gq65dQhGl/pmzDb4H6eEgbXDRwUwYM
t1YUuA/ykmFazfmAzduYDt+PNxgkIvdubSHrhNr7ETvrEY9di3Z3P2AaZviRVIFZRsbA0whmgd1M
LOFWqbSJBBDkGu0x3hne+AjI36jUUeJZx4NRAqtMaSuMY5cI0t/jIBc9Oyt51pRDXKi1ugl/lz2X
YGMcR0FASGsvgaDjxD0PsR2rbpmsq1l+ooV2tp1jyiScQzs0kn89SRZVisnnZ7U27KRXt9knFt/E
+S3+a7KhGsdeP/MuLFDn0vGIns+gKL28aYHHVXqpso/Nxi8W2wSx61TiFxKkHdSxnIbqNKwX3qrB
zA2U9rARg5zP3ejT59h6IKLWpFvVnnBmAuWJ8UUwEdSSq5M+Va1J9eHUs9dGrNNl57iuwvTZwSJb
73gTearVQ/qSAZUIgckVfbMbnYMWcgFOnMYOYy926j7GgvdrKpfirBf2A8KbB1hO3/fOKU6M74ma
xZb47GUuHVRzEfGycddaUSGqci1QfjT2ZMP1dJgsNI4eHBjhpHy3Qi9kItG1dceAEXyx7lDkhvIS
a142BK6TbQ4LokZH+YnSgUcnFMeBkUkXfmJJo0jNIfC42m9NqC9NNVD1Num4BYtUIPOJEGFgpywa
5RSyfI1wptJThsA+4Am/7ZasXKNn/eOsBPtOrppe0JrmINhp8X45Jb0ugKSnwdhjGD7tNtew233n
+uZklBKVGOiT0rdPbwupNbv6PT64PeqAWwikIfkfjMeYRZVlyIW7NAFdyvCBuXW8oG0gbNPmsg/z
F7mLgon0whseaXY9g3e8+CCGQ6VGHoC/4/TdYQ+hTrvl9E4E351FSz2KzUEmzmb9xV8ph+NiaxUm
KqzuXAmp4wQGP9abqY30PyU8E1jrht5+4DpowUccuuQEiXr2bFz5SxMSEpwwlbiDtAjCrvoAM6u4
qlS7u2Wd4lM6yOZ/dlEODpsYEX7NNgTEWJsiJJWcPX8aMLobcbnPyUh9QirD/Iu7MyFPq486aSq/
0hI2DYh+O0jx8PVxXK07Dmp8D1oSrMrNX7UUAQJoD7ycsp50JReyFI0zUO2Ej90/eQub9YafkSIx
q6cFym/7AHw+SqwiUzSC/rbYD23wkt9W0adgFiM1rigeCXQr7yHnqYm1VNL+WA5kNZ/DqC2PUfoE
MYdAu0tuAnY/OpgF6YmK4wMVbtmgi+8aLr0ubrlcx7vukaRWBK6hkrzoo48//9pP3F9luozwC5Yr
vS5tEwk4K3/WFjKjFVqeUVtpuW5laU5sVJi6rhrScF4NE5HSR8bLpxYGEkYCXukKUIxzO1f2TZzN
e0pM1fZcy7A1F5Hia6X5VdPDDM2CodjCllODUhc/jjtkr5MPXk/zNTOeZ6MkMU3HwfOSMw2JT5Gt
iU5cmzCgTJqFlx20A+uxN7KzJlgBjzS5245py8wcPRuVLFX+GcW+ksrbrbmVRtHQL5FmN9co/weE
D0BJPOn0aHZ/qdfY4H3MC+GRG7JdR/gettFbEHaIxXljZ4nUF7VTdsncWCnFehDxNgtOcBShVGZs
5QQbLoHwxLe3Lx+rsvzvGwQd6Fyk6Mm1r6dtNYqjU5AYiGaCUUwLsRquKxDWai1hMGgm+SV6BC8u
WTdoYG0+cAsLW48yJn4tJK2u7B+2zTYiqjmQJHYWxqAh+DhxHgp7M6pCgtfvwZ/d/g6Jet7wIsU/
nSfSWoiBVCPJZXitBZCbwXy2zur21L185e3cdWgZsJ3l7LOd+CQ0pqiYilSXfnNrXHzTZ+t59nXu
USnVW9EdO9KJY4owxJVthOND63QfSii82SCKMWGA6Mzi75dJYxQvXouXgZ2NzTFwjnzYtV18Kc6Z
U0sQSFg8ELLviJHW75q8fEjWAo6I49trYyZ2gOe20uk0PaZBVd4zHqxXxoXB+k6vLpWs+QydCWL2
3uGUs6yvqu66cLg60/2NjsjxiYkvUJHW3efMj5+OjDYTpmOpiUtgYZE7Ctjlyrc/Jg03ZrVOuEjz
943DPkC9WuMy5/EJCVHNZhLHXmF4FYTwDm0h1TlbYE6ZMkgqI8uzzMNXn/7GtdVaEsNZUxOHMNf7
Nve4dqNOiV1xAd/JvAZA+7dsOezz2xu1gBUmQHfc+TIKGAN7v60nvCZRY5dxVwcjND6UuOMP4gf6
qTYdYHIHUmFy/qV5nVSWQt6Bz4j2jGzjeg4xumCSe0/CUTy3JkA0UMkNza7qT3ttq7mejkeqsQ7W
Ana+eS+dJaju1oFcQkhv/y9veTyYlG/kSto8DcyDqLDijOw9E3M1LhWgDndZkhf1tBtCZdzF3hst
Giqzbyt7nGk7emWZr33MJe1DinBZtu1QSjY3XgIVf/jpkKcLs2khswuAfiIahyVUH3G+vjAI5dtI
LLm8msEL33cU5mEH0wQzdatVAb2SkzS9N0TkdB6T2GOm3S6gD2k1v2AkOwhmz58Zq/5dDa4HFsym
9uuWkORnrpavYmtnLIVmQIV7dqjOwbfdaoU6H/i3dxxq/MIxUl7QC2paaTiNnxw7et8/hdrXTEYa
kdj+M8+lvSELLQBPyRdF5re6u3RFH2aKqNJhkVfCuzkWp9wPCQi5mosMxwfiCxDh67ux3l4OATVv
jHt2QaxE9LoZ5JBUqpq8F6MrRMYWnCQML45pyI1pzGvuWMDR53VA6x7KgwEhOQd/VPPUP06y22tg
l2RlHTKynGLnXviU1WoGYQkczjZEnPvGOx9WV57srlc5wWNOnfELyyAfYCsLHuFFijZmHjkqSycR
pI/IOihi2aJwEa7vw1dx5XteOqpJrhtvFL1GG0/PPo1oTXF9sD9Xjz//gEKEaf0PiX9mQL+A0bPM
8lrFWveKfm7elUBJKd5QRPQMvxZXy7iZGSAlQmK2Aj5vbz7m7a7bZvuUxi9QP1DOvK9zygX2cZbL
Hfr9uhYqcxvonPyl98t7vpMZEZ32SqQ8j9hNr33cYQ2tftvPdMro9Q9zLq5h63U9X8ipF9bd/TCE
lLotspEmE6x0vAZr0n44xgzGH8yD8aylUCtHoALabKOxo38uq7jMa6k05hTdsjkNPphukqV/esnZ
YSzUQTc1kx/I4ItkPnhKB+P48FvikiOPZ/mSA4fNGdTyoYzkpWrrXXbKNwTVmTZGBdCL8uaCRhhm
AwFN5ZQl1odG3FWmVmMA+1ILOtqZs+UQFkpKzTAaEnOhmG6zrEizDt9jm4e4Lr4q7V5fYCr9Zxxc
omP7hbKmzd9gZS4xzjXIz/SZtnbCAQDCnNHFp+f9uIihespxcTSM0MypP4q+kISTLqZF72AzxjNl
O2cgCfbXrNnie5CP+cNT0vkTQocXzLWM2SRG9CtjeHDWFvW+pjIdOCHgssB65x4KpLwHghhL0fjZ
XeFVzBGTd6I3agMibjf21U0nUfrHFeNKOF/8XX9DfIugIjq8MAHyKLs74lAzFiq9uueijBzGhY2s
K9a/aSJ/30e0qRTwkyhrPPpskwXyVyYl2rN3oOuoL8fVCExy/lYSyQI9QSZq7y9oUdXRP9uuzjch
5cCYcfwtW+ZJWj2jGRtm/eHegOWnA+vjXKWSNXSGMWArnW45/JZEYoHGb3OOHsyvNOlnF+BniFRp
FCSb/bUgLWrVMwqByQLfGPGux9Nx5+M0FHK8nwGGZodpiL6KiEkmnp7yJLGoN8v/EQLumCJFQ2lF
mwIwnMmowRphOrhwu2yIrgZ0xCM2S+4pjQ13ttXly2VFHWWCJtCPIP9A3g/eRxvK4KCZLRrBRTyd
BAcrX/ZxlcrYcf2gXlAn2M6jp3C4xK4ktcjlQZ9BWYrItlEDcd/PQ/3VAKlgwiUeRzVSc6Qtejt/
6LXC8Z7dVUJ9QcjSXZ0q/BqJT0AEXVxQhPpau8NNzNgpnNhpWnpZksmrvtT/uSd9Ecihen41qr5D
Ag6KUffql21V+2WrLecJvZZ3m0J0No/4RIIp9idrLkaFU8DbAvEH7VAPAiPHVsZvZrcAADTUrbxV
giILbgKJBy4HdC3JXxjxQd8ImEnAovyzW02utbGHPfPvBCFE1uAimQBq97WxlY24MsKU288DIsJ6
47SsGY1uhGJIBxVIRJySg8kqS78LIkSPPvYTFFjOuTdBeloURhL2o867f+iFFfB3fYvul98oOdY0
AAmuoCiLCqqB7ofHVLXQf7iQ9ksBfjLuWHirY8ddiRbbMQpMZpc+MMnsMR6kOaCxrAy9D19FI/8e
4XH1fLiDP1RQs2uMAKxCOfSsBmap55IMFaycfZgfEZHICpYKY/Nj5p9vmr82j4w55fvtrNi7yg1U
7WLRrShbr+o/xr4GLLQKtWZvhjgN7RWSjw1oK9R4LAz8P8XsjYwaaO/Rio193hGGNzKb0xHUTO/9
JyxuQuYXlEq5QlSBUnDfsR+tpDOsvZiDTfyFylHFWs64quy6V2nVm4Xk7r/m1XNGDUvj6M6xkAW2
QgBulykkNc2i/D9Gw+SsZJIeiQ3Tk0v1rL2vbRnbd42yhYgmKO/L9faDaO2gWB4Y9d6mh18YtIpE
vhz7ct3oYIkt5qfN2eIUX7zz0i85ABRj3ZTBV3daQhvOwp00I7pXLwjpsBOCUmlpBVu9Df7mPFJn
DeWfgWKXNgf5nDbYAbZdIXg7i7RourJu+XiZnIcRHQ7brOZXABglKxeKbcOZcCICkyFRMkvDBSs+
Hhq0xQb4y8OzJjlCZflmcgGAfnZNTONct27XPXepQVvoyUjIexhuIwVG4ICI5XqIl9MoaWI+gCFP
zLaqyOIEWoyO1hroNEX1R/HSL/1XQafMVkItpkgC+qoZRjLk7xzpHZetWeCn+2YEQ+IqVK4aJZZP
H1R6rdpTqfesV/1C9TRkEDIWTV+mwmUroZIAs1tlv8ZjKddlm73Y0oycwTFZwvvJYd5V4WVbPVQn
Dx18nwsVthYIrtwDAAZARHzI3Yr78x5oq51bw3NHo2vQmgELVkwG9C2Senb+ViTjRi7diXbybRQ6
QGNTHtRlRUOCljhsOxZom7ouBM7V4K7qToCML7FuoB7oXNQeWtizeFzdNmNJ/NHJkxSg66KaAZxL
vCNYRPX63XYumOeyiGN8nveaW4a47NZby9rmXegT+lzmkEk75VYfsIY4l9JGiw2uIGMUPlzfS8cG
q//QfgnXy65eZKHbHBmBOUyXCOnsKU6Wy2deZAgIcyiXBybbXGrZqAXuiTHsjCaj0VWLSDUAUlYF
HaqfbqRRpWMTeYlEeihHeAoQfDjVkW8rHOYAqfmmeGuJcKzKYNtAaQAT9aJGGw/idfna2E0Vl6Ne
jXDrmlyOXJLqpavfrCRjBFH0qif7Lp3xAhpLKTkYZ7ipnq9pT8gW3YSL6QsPH4Qy4UwN0PjVeCIU
UkmPerCE2u76GgbulnEPCW4RWuzqm1UaD/r60f2VS74LFu6DdR1e+BJzsavbxwt3j/2g0yGs1b49
4ioQLnJrKFlGE6O7o1RmJoUrMrVCkp8WeyEn5LgRVekAZMX9M14lwroiC3q63X9ufaZv/Td/3dG+
bPAn8IqPyYOwlV5+zAIy9mAbalWJTOdS55RvhidJ8spe7Ja5MD0hMPU2legQq1hJPA1cZiOzgsEL
C37ktSqNgJF2vGX8zzX221xW4IJRK/jLp1cSL0uAfvu7RmesSiw8Lf6UXbR7qYxv5DUt2U2SASf+
0EWk6yePs9Kj05RkUDbFUv2uawyKsxRN/R+mZkE6ORIuxrxF+G/H0dJRzebElEOqIiLPKR5rd2+k
27FSLK90OxKAGa8NiyOQ8XVNQU46DuhApQV64/afL9wWfPdsQ8aGYSWzy+DGfi+gbGAOyshV+Pbs
nuaWpDeHfuDlg3zkZHgr8v4/uKoKvE83ezbqUmqFf2Vs6FLStr8HZhmuPqqr1d4X2qQDbiZH0GNC
07+Pt4P3fyYsXfYfGBpz5aZAPOzLmk5/OnjnmPatsj3WTGRsTFdjAiKFDc/fzJ6uPIJMMzKesMfe
7BYthe41T++/Cg+uiPjOYIlqh5FXpQ/KsprOKM8x/GZabJQo7lzUYZJ1K5+60fgu9ZyburRoNqMU
yZJk2B2jeSInfIlqXzhTMbEPs3Z1BRSpD+1jEfebdViPHnva59rW2LJWXJ6nAcp0mJtvGk12p/KP
LN9uW8F43HNo+I3daafIc978zAgT385FheHL15P06Wp2cc4gwUa3FlG7QkVVAVPYfQnGyjaXr56W
NtlMJwGp5yUcXPtS3BfwoelqA3iVvZyp6uIFcvvxDNish3Eb3VvvCdAw4opsDLqHGT1RLy7/3n4m
ztN8znjg9PQg+7XuQAfm0EMY7j79o4XJpteTomIUP1mCKQHUek4KSUZbxaAZaGD5LwVvbGF1poDz
luWIVZglaVvoKhOwc3Xm/pmA5+AGsW6uCjAodP46+uhgSQ+2PJQj1ygJIPhviiepx1AfaVbhty2T
Fh2vF65FOceyEo36+/D4LgKRutdzP1Tz35da43/4CO4dgVTXMHMasTZIBSEO7sP5mxSlfts2vBZe
Rb9aq5NwPJCkesbzdm2lPCC1aJmDmobby2zjx6qFlS160GzZOdOb52eqPwvxqWy79+uNPpIOzYRT
XmSc5LG4Yki6OZoAJtwbcaijO4zJWn/Uc5WEVegugcx7u7jWNO/us4tP7sC4qkYMshtTQchx1f0H
R9COVWGA0wC2hFiMghr94/V/PYNk0AWEYfOMmA3BA6Ol2wmM4nvGV8ITmkPSg5dM1U08j6hzONSW
MZ81+hCrVGG2KmdFax6hMoNTvW+gTrtppQN2r1YmSF7FrlOcpaahNo5zq3BzNCkiMHgwA3/SxhFr
x5ZSrMMRob4SXL8gbFkvxv0fgHa+t9zUFpvukkQaosDSCsjnvQuFQPxpLh8SCQnEovSJy8VUZTJq
cT2OQ38nP8oXyiLgqLn/9kUx3NHTGDaG6OTl1E+mG7KxGzztVPDUqWoRcqDuZWRmz0NEDXUbe898
Lrf2Gep/1O6983+frn8CSAAGt1t5ou00AxoRq26jQiylFFreKVxU9usPzGNAupN3ana84iObitW7
RWItR5hzJ1z97pUIHUgL2TNvuESWiqSAm11+Y2HhCy/mfLU70sRDPCYGUaARqHEFfNLXRt5+a3aZ
Nz4YL/Ft0olJO+RAvS/larHnUj/OhJQfRBBFLQwHowT8m0/kRWXHXxjpnQZql/JnctaSxNZEx+46
UG9dQXuzf4duS2tYTOZyufg66YOz4LiwZ6aQ0JFKgO8BJ82OxYB9Zj1XQxelbvEXUNtJJqG/fchw
TrayZU1IUGk7rmSS23gSw6cVaAwQL+J5VbbZNCuPSq6qu3un3yRq4LdmPZL2bkZv4swpHVXjnHav
MZJT84YKHcJEPT8xEv3MpAf4Q1dgZazl0j++eSEKahy2FfQypO2KwtiXRxJtTx/RDghpE0nyB+YY
EOk/blrlrLYI0j90Q4Jl9qKQTRa9VowzlojNooJQgs0KrVpmH3MUJz0Xup1kuilYjjW0AlZZ9Mzc
hPIUfT2fFqcEkzv6994uwYa64b/tuySXJ8kDMH1HqFcHybIB6QAIa/oh6j6y90PhotDt0xaL51PT
O9thp5O1oYFoPfW023y0/naxyCjguaM1qDJ/48dMGGyWy9cOt4XYoJInLiAJG6ZydX5KDJzT1Ecd
7Nq6gKAkzR2xFYoFb7poHPvc11kgAMb/Iy0aJ44fkyT3LgHbw74gQ8NlF2Nxe4urRqmRQFSXPIQG
3KzrNEX9V7OBN5H9vCJDkmtWaoX9WjdvWJLsCrzwgOepSIblmK2OVif5M48cXi6j8g08CoahB/qX
nDsDueEGyWBDWNXK2cV+AgDbt8nFOQCtl1D3jG++/BkTH5FpD3bN+ShKEmSwuuTVU/sM/Djppd/Y
aKcfcpuWxx/BQF2Qzl59CNMHm1aUCRTnDjFaZHRxv6nXvaKCSYlkkCnLWDzg3FMogRwxL/O4M7kf
hCHuBneqH8s4tJLz3qs5madQMOWuwxX3bts0GEGz66sJOi45eSPUMosINNRU9KBOvPxS/zSlsMIW
f8SFAx69MRWgglTfh1js4hWbBXn4LHyJgqdD/zfMpdYt3H9rdUGaGsgLvuuLNdl8VmH9zWc0pSfm
Lsk6jxvLPebk8Z3qlE1N6KEWzpyrvXIDPj1BInXFnoLWw+2aEHwA6wPCcZd0Jgz7F5vbu46rNl+y
o8cgDHFVpHtY11VofM/B3z+igMl0ZrDTI/leFb1ZaTGKNhWf8zTfio22IvsZFqqtrwcz1evvgFqn
PoOdjHejRJ3lRzZ24ZzfnqsLrlRIsz86ZCjZ+Grk5N+JWojBbr9Dy7pmxMdr6ty2zaV8I+nkTM83
B1us1FOuUOIi4pN3AIhZZpoG+5Njp+1TaLU5ApSxqAOxKPaYbtQOevwKMcj4jLaqaZ7QAiKxod+l
fwXDctALrfPo7DLzCwb+x2ln2AxvzvI0h7voUZkwT1Y/oM0Jp7DXlgffJrCnC6xhziiPorquQd33
Rf11FSz6+apMa3yMSy78Qty4WNtPDhjDUdYfXHTThLO5tpjcSd7Y571Y91o4DiAVjVw6Rnjyik/e
GKNDeWRAMKlscbo7tpmwYjlGnsvA5EKu6creq1sls5HjjpRDkG4006m+Usl3jNUwloAUQt/qtmf+
sifVA+SprRh5unH3BgNJ5dvQhUeudFPBDTADzqyTxF2SFsMQHQ7sCBG9rDXVHsZLtsb3aSvf9IFR
KbJRE+nqLyuXW43e9ubkmREjS5a0QhrVIuhndGCwyS/Rx0bTXF1d55CHNmqGec0gpO02EXwrQvTu
C6Le9b0Ggp57zMyPUdvxHSUZS3yEHmT9cv5Rg6aTVbjQs/sHcEBqajyzh/SRc5PiIk/ngEdhk0NL
zwTZjKsfvr2FfVkpalzNJNNVRHj9PRrsqisLPXGCjvLzfveeSLVQzH1ivMYhZ8/r5i2JtpoNPfPD
FJKgY0algktpR1+CTZoZJxKrma3q2z/udJ8cToto+IZkrNQ8CJnPjeoZyByYcsRX4go2ClROLdFF
mwCNIcnsGQyxwSMkYNRcPZ/vBmiJCg/b1XEqLn+YjPzy0ilf8iWTAy7j6etyP6IB6qucz4iVEVrb
iWdlZUzOED0hjFnZMT+7TuCKs8+h0TTRabOblzb3kbvWAiZOiAmo5tlaSVagH/b/Di/9GBpDRaJS
wofvLI1TTd0f97Whsag9TvluyGd5mnJGonms4qyQlMs9Hm04PhKy/ElyWq0iiF3HN3Vlz2UUSnOR
3TrmjOzV27T0tNEbe9OEOJd3RNhg+MGNFsvfzNCXIkOPHR4ntUhYpY2bpRU/Is2rfuDi7hCkMvwE
zIFQSXFtMX644M+CZbmH/zmfnjZc/ESwi3wM2wrRZeEvO6egIdUvhU/XKA7E2yjX09ve9Qy7Yu6R
dR9qX0pNGUoxphfDTw3E38iXbGObWbeFSo9SHVoDvxt+s403PKU5hkEsLgfSZKYyGUwpGb8dml8p
b8qAV3EeWe42OUYSFhAUfMNoHT0V1Jw96cXosth09stTo7TQBdBpepOuIDNGbvMFCkbrzKmkQ007
nDAnr+eVqmP85JxL2Und9lVIg2c0teX62P+IcQ89Yx6xyCuhXTUJBuDUqORpEIkZzfiL7qRY08i9
th4fToFcbdwgSgLoip1Drbm+Yep4EMTgYWX6kdlRGoXXFYzs8rJyHUjuSNdJjE0MgiIUZnInfFoC
yZulpw2XYF555tIyxmUEawnJeMFLeWJDqpC7MyqWXVTWP8vRFIj528M51HizY544KuXn9rs82/Bz
SdPq1d+fUrsjEMZaw/p6K7ODtFXyTebJZ2txiB4fXQi5H5yJShTdUNGIlsXv1lVtRMViX/eQFKF9
bp1wPPjJks6xhkDJ/cQxoB2p874aoRak4+2UkVwZRaMfS0s/1FfH6ja1IpEfrhLYAWhGLaIV/Ez5
hxFcIGZffMot2z5epILcheDXCZhj109IPCM4DBskdoGJdseKzi+pHIWp7zq0pwqeoybz+wHykiv0
pdpDpMRf2WCUy0cSjGyVZU2A3N7NVkzjXNxc0JLjAmRlquw3z7pJBbAzyAwUI08USRR8HcDpLXC9
HD/Tj6NDrzDXOApdOOQGzzyERer2rRQ5fl++yBIhncRw0/y2/Jmdb6nUIo8+05C803+wkRyO8deY
HqV5pdqlmVu7RSB/mSdxZWhkP6plTEjRqD57BjwDvLSLOML1QISRHy+IB9lSliZ3rasPWTsr7ZEv
RpDfVGFxwabZgptN2lb1VqUdiYWThxoY9trJ3nGyr3bHzTx/MOmkKAnxqwR/jDtDvSuksQlPyejS
2nZ8odRv+0FBut+U7HZk5s9x9Ux4+PE0Q1OFvp6Cd6WSzjHSmp/XK0IDNSm/zIN4ATLcLL61umYU
GJbQHQ0/HT77taQczdOfSe5EXwvQjbOeP2T+7xJ3mo08rOHVkAdlohmjDIxR/RX2omSVUkfqLh00
2Z4ENVh8A/DX7lazKxInww50pvUFlmOIUwK6Y12sIlCEsWfqOthSJpv2TvLsKgUKTci7HLQ/fNeR
Ij5qdr7ZS4VR5NW5fbkzstgZkmGi9m7wEBpBHCSkoVpDeSIESy9qTHbBF9WE0d+MQJZpE4OpgNB+
ni9wqU8LvT2EPtguTmt0K0h+oPbuTp7vXpOh/EfX13Tdfpr9Lv6irGsbtGBgqn5LXA3MR+qA1w6u
h1vOurXmU5gpGGulmkdtAaSZkg42vXL7vnUqZyPPBDvbwmH7W34qKkaQmglpw0DJ1ODxA5DOK9eu
T/y48r2EpyfPvrC9RKyOmhUkcLW2G4m7PBuOdoYvJfs5ChMallI96/jRU7gUIBJnFIZilMBG0CsN
i3qS/joeOd08wjXbhRqAgDB9quf4dqACZAANnqiVTiwnqPSsJdO/7vF+0VG0g+d0FCaErwpULjZ5
SB991UujRYAzD/cgLiW3DKY0Awog3T4C+KXCOCsc0SPpPXmALbpNb1DzlGj1yPXo8gOCE/fTmkQO
JCyE5x+Buc+j3IIsDDqCOZWRuClSf77Y7p8DPoVWVjEZ9jALFpN6pBk0Dl6gnmwmLg1ev04wsBCc
5AocTRRaNbVwM4rqxLro8mXYRG7GB/YnHIvSsBBQcTVU3UR08YmLVN2sf25LsY1M9bo84Kj+apfq
HS90hWX+m8SITYHNPsG+Gcp7vsa+lhXD2+r/KQ24qS1IpWRDaGZFIiJngSrwa+LmVOX57Pav6XPE
y+Ulonlhde9D3dgl/u4i/uK57uHl3CO9txREe5zcqLlZMEVtBZm+sKv1s6kdvAtHSvEUm+hspDE6
QoQBRVsxAJZTEiccFLz8pENQkLdupgafZEMm2GdI9vitYCacB+itgHk8I1Tj8psKLDOdMNVvio3X
tQXedCyMhglLjLo4jYomb45Dow/6JpP14xV689Oso1UWi5u0Wc64ZyfK+lCal+Gf9jivjxHRYO8x
ULvxeLoWVL2NuRpcwmpncDlVCxm0O3QVxrzY4hHEoNNq61ilb3OIRgTQw7xw635yEMcMSYyAO/Ed
0mROJ7B441Iz1SIlwnkKpixh2rKSd4GGJ/NlUcLDmiydfsQvcf9Sm5LfSfaG4ivyEsJNAHB/G2Fx
mHg3rxbwO+b0yc0NLJN0o5op0kAQcl7RNfCKjQkpxsqCFl0iHT2vcJNV9XRDxeU0gO2Zi1r4KmdK
BtZc2MbkrWOr/B6woY597l1XCKcAidcE9z7lQ78wiB4TH8hLuramlyy8rwErxn9RKAXVmwpoPFl+
qlPGerOkDIpAB7cq+2GSSDvxyhvhEIOYIOhQCh/u62H3gXM/TKLYFWTQyuwXbUtb/miXdy829nZv
W86rP8j9JZZUS22Sl9q4H9CqDYkAgI1D9rg72SBMXyUEoUJIrf3QCRWOfGZz56c0rFOdOlffJcgh
+1mHOInOpzBLXoaYp9eFx471rvfmXJsCuZgRTiDO+uGXBY4bVQT3bn8cJKzHPlz7sQc3Z9vGXiN4
LECcbEy+CjWQXGew/sZe1l3gG1p4aCQ04pqpouCK85PbyJfPoK75bh5nBWggICHmLM10Gox4UBcI
00kaAYXJAW+HDyp/HIpKW/qKasdwHmaDfh+DtQyBdmjcHLep1BicWMMRv4+O5MvWoVsTLw3CsoQa
MBNQlHAPo/hIhpMgqZ2OYl5kqrlAMdyKzrHKmvmXiRZd49+VdLVJ9IBYcGqTUoUtJq6Gqm/APhsL
zPxHxLmU2bkKQsDAapEu7YvduHv0n8iDAhlleACLpoRWTW/GvBqnGU3mov3NjQEzm3K4al+9nTxR
NNB+UAJtrhyDFccnOS3KKZoUBczLUzDzz7Zn4uyS80rpzbFi0AF1tSz6PYSr/a0YUjRmyM4M06MO
Aa4KwR3AsrjG9aEkwl/VszK2wJrE5fOc/s8FeOuy63vVIcNGMHv4pBrm9QZ5x9E+HBPtusZ7AHur
GG1luJlR2SYTvxmuA2hqaV5lft6QeD4JrpdHaMapaMg0trLHKs1jhuV5slSd0H+96Mzlpwn16X3F
TDrlAHdd9cJeCBYnAKbkFCJXaG9BDgsRKahg+3r+IgfOqIhjyeriTlXownhPoyNHn4Ba+7e1TEe+
oEdhUvB8Y/MUQcpIpHTIuVfdcH8/bboLYrC+jydVuII4nkTRA288nKKdqAN7gu5dGuOoUnh4bTQD
c6HkLDUTXh+RcTuMyVVwZ74rlY0PoVwxdDwnptZ+jbW/y1gb2ffhA9/leNdNPFsZGLBAYFOXdb2T
hw4mtFXQdXhUVoJ7wjG85mjRnIP3kVTavCbpMzI2JJhIPyheoM2hXfvDG+gIYRMsvrDjbOe0/0ZO
/RsYU/by1fez6sBiCE0rDyL8n2LIRqpnGeZ86oupAewCVtF2p/ya67yEhS27T1BguNvGwuzA5rPM
R2E+E677mCCr3gvRhK3MqWX8RzXnADVdlvR3Jw61kshPp2KcWxZk6To2DZ1I+gQXWeP5aBhTfdWp
di93+PxmUblYWMOYHnN3wk+ROegxJYjReNrv2yH8OnzEcY7kvSZAx9mx9ZIY4+fe2hm0Cx7PmXqs
XGgNh7/yAVYCPfrGHwhe1SwXYYA1J+IEb7OzylAuIW9cpo4jZuoJ+kDUgxiQQZ+XjZCh/asJuUhX
879izYHDTjo2cylfGVoXj0gukZsBdj0rVYywk52ZsSAbt0Cnj+uF8A+jo51GOqX5+8UQqFq6c4yt
Si1JA9prZEEerChXM/ejo2d2rQ4ytU4JCQl7JGmaTbp5isVBfXWG5GVQD5UCn7uDwYF2MVt4Bo3c
zjtR4jXfyT6SPvkDSJATdt7SxkCsoIVemPNpQP8ljX1G0Txpdt6Bwk6hqQktchHKnBSx9IDixxyb
1n5LY7tlnfyW6Y05A6/qEUWC/myZdbjUOHqIjEUyHExTSGTGMdy3bxT24jV+7qrsyWVhprel/nkz
8fegAbBXLUdJ8Fusd/Rl2ZQfLvOpaWWSRbBdjka2zDwnD4lVIQ92Q/9B7Wo8ibE24HsNF3ew7m7B
8WZwrHslEfjJ2oPFPLGSsWW8J2oPB0S/fMYBHxmX9kvM7gcYcPlZ5+HKPt0ox8lFzcNJBuCLQXJP
HUda9TSdL5tyKiHJ1JUAyxcBBGDiTAI+5xNk0gYbPQoDrMemDcmP2K594eP3y/+jDUUQqmKdqae7
Bli4usexzq25gi9G74Cx/CYVtboKlLYx+MQ2FhXXkliWitbEW9SBIQ+ObFIioipCu7XUueWW9B8M
49/QzzCnlMwKS+7xih5/4Jbpt/X4dpMlt8gZQFF56FCNJbt0GFkzcDMsN4NOvu0CZbS6yQ2yCGsH
FwD+rOkpOo8CfiIVzDaDgFtbb+gjIjs2jbeRJaIhwbI7XUiAjzOYWNNZYXmUvuyyUjJn897o2wSo
KgwCzAff+ZCKRDk5e3TwC1LxGzjdc9o/Zt97V/ZPgx0d3po713FTyga0LiOIe80SrvFQlDO/W0/1
+a13TMgDLi9qfn9UsPOddajC6HJayig5Zj9zY91q7jvIpWdPtx3grjZFihLbEa1zUiequQCu49bm
YXnJlSt0ZuMe9SZcAxnJfwJlopvBZalLwIfcDYvY2OpvwqPfnh/H4ziaUYR7Qy4dEBLKi2UNuymM
5J+uKIvVsLRjM+kubhbRpHDnUDedy394pSawNLgSpZmP7010YjCgbKHdB/EYu6CSfr7NwRObZpP9
yZdmF93WsO5x41uo27r8kPbWihDIcl625Bqu4bDCQKp1uZwWNEIzxlVH2AEMJOWpJr169RHBBcp7
vku9+0c/VqexcPjU2RhNIX93eYNjf7Y1icNZAkwF1iYzdrxXvnCn3Xhq/ZE4ZgDoWDv8WKB3rv3D
YMF+tIRQ/zn8c8k15cGZrUauAr7TJmgZHrGa0/yJQOtgFodPVwH3ibOLKs2xuBQzk+JumAoNV+dK
zJyBK0ncPdlyxJJn/lwy5m5sLem9KbqmORwnT+/M7hKHKzQWqpYxzGSDK4m9IsqUdhnZIMN4Fd7J
5Aw8Jt5keH068KfU1DveUj8kTgwfpDes7SviBUwjup1m55vDFYaBkNVl4gaInjt/vmj3q9KtZ9OU
TU7I/ksp1kEPjIH1Tnra1UjAVagVSus/WEhdQ914B4PW3mVDL8n3oSLCk0yYjcKBIepPdfL3FMS1
ZLlhq2tJZpJy1ovnFCOGDeNMm3c6irFClvuv91qXbIKGGa5lpNPj4drwPSHLl9t2U8eG6csOrjSh
I0JmCMVEhNQ/IcjjsaxpAj5Elmry9nNLnLE6ubqUDKY75WMYOEVJ4CV9yz+rHzBmF413BAELUpek
VrxTkA854C/QX+YN+TTIkvL7Hbi0boSc9Y40Sfl9YNTdbUzpZbbexmiqZdWSv3AFHPYSHFmXe+qQ
uR9dsdiceUFPY+ne+FkZlEvUcv7xHhBqDFIocG/wBOlM8inD/mfxs7ORlRP3Px03IKQ3O4IBo+oI
EMxGQricEYHnaaeL9g+w6K1NhGInuJa5XhfKFuNw4LmXsANIZJfiKA7k+Z9SPnIe3XNZGhRDhPdZ
6P4O4zOiX7FGU+80ARXDT0q0lEnEKEtZq5GzBH9uvzxlAQSnGPoyrOCIY9rPFRqZUVq9n0tEPlHx
VID7KbzA9YdTNM36rfmZ8BZNJQ9+2ZdILpNu7BWUdY5MCNqW2VyLJRHtmVGr2SAW46PvbCSujS0g
fHtXIND+KuW4StFYku+Rk5cZQTrl6kjl9Gu835qD5HMxGDkMcI/C89IkyBQvdsy1OOB+d3QDi0EK
WZkhfMbvZCSTNXpffkIDjcY8uaV+fMTl153U1D+rG9EB9jN/0HYlg6Pv+3qDuheHHhDh6NdCh2a6
jl+0JliA7NYNaO5CiTKwV/WlyQfmcWrGzZR43PjbPvtgG5eGSxclIeoAZ1TXtBa/JflQ26hjWsIF
+20zkCCB5pc9iYnSNJGMta2AZhMMw0TqTVwic7zO7Pb+oP0A/jgNL2VaePKlazhW+yQCpnMYE44V
votHjsmUpUDFa/NipIE9O5Vg+RV/biWBT5PZ1N3+PCW+wmrpCYz6UnoQoOkGKCQESX2cULcgUYKi
VW65i2e+QxhliX2tri7j3SE85xAyscvKz8HhZih2judh3DDT2RjCNlgKhMh0CkZ5SZ/1OC6L4Aky
pphoCjlOnkL7tsvVkw/Ampn6hChvHW5DP9FxTAQ9ZwizzSnNYcGs2AFm930rZLscwtkcHSghcZlM
g+zgZJ/u/JnuAqLYbdh+ax3VQUfeu3RmuiKvu2L0Po4tQjVa1RuHJRzCu+kTuE/2AaNsK6Ciqyy3
nQJMWk2VgZlZ+EEgERuVKT1meYZl2E9xQ2KoFhmns0Mu5Y7QPdWWXGrHr2lAA8u7hzbKpB743RQ+
cLWgZXw5eJygN83nUxgLyyXApGq8gYPewhBNnDSrin08tOQXjOSn3/8Pkr7JGAzSl0YEd+kRXKcK
uEglXrVMF26GZLwzr2RUBNCoIr83FNy/oAffnX9Cgc0moVRrdN1LAuqnESoJ6mKDkjMlEHG8dbmW
PY42K+I6f+vXb2xUnQ3jhO0fyuhscEzT+iYXfob35oycUqH1DlwSah77qSY56IOSVD3y0HBc8hjD
N4p8zIdKcM4hCeHxGVnGHPwi8T2NICSkuBvsykRejFj5WPQ0WeE6BBGZqGgB1l9FFn/zkIvatqBy
PWGsD0lnQ3CWODd/K90cPd+yHxW3GEONdYdH8gpXxOoGBQrBNKX/Byq8UW5zag0PYzwRorJAGMRF
wQX9H/8y6yXSrrSUIhCk1nwjfJtvKwWmn40nFL8ZpLxh6lN3Vh7X2fY9A5xBOSRIlL2ZAJpCKQ2Q
BZJGsrCZ6NlcUc2m78zpefcf5I45R8tMBE+6a3GHjOCwvQF/uQ87f+yUuL5h7qHvRO61t+ndehV6
9kaIaJnRWPgRcXe+6wnHXMsrl8Uavaq64pqB4H5hcosjTjeSt10EzAhSpRgLYw4SfOCCmzXn9j4a
UyjyVTA2rH26iPeW+edcBg5V2pumZSkOMBcBIzMfiRafr1Tbo6f85kXBAfiQMFDzD84UbEMEeyex
uvtOlB5VBnbY4kACIZOnB+l57LNn0Knqr7TqCiMFE9f18sabcHzAbBgCO4+A5F1UOwEn20kgLXS6
pklM/cfN4eFMklxXn4QwCzYujuZcUmICfHOtRekGts6FqjucV91DbVUqJQQcS071LzoC8BRnjE1w
XSPLjNrfvqzo8e6y2RePhp2SHtJ3+pU0tWLp6uJTZAPTaLfWUiSIiTXjJPsHBizTegHYv6ZQEcOD
4wJABcOolREipgrS06AMyZLO1HISchipxeUwPg+B/X6n9gXpqHmcqWWEJKRVY3H370zPk8z2UjnC
CnVmQTUAQSAewKl4duy8xvzJI0n4nfmz63DlwbJ6Ap+BtU3K5W3AbgvKvA/BkM14xMJudMVz+uXZ
/NXbqlI2v5YufX7onObMjG3G60ESjwM922pqo/HXJW0xQJffahUiGsxMREqo3zz1sqXqRpGlg9gO
hn1RmKVthd0cVl6byvbH01roaGfpeBg+ZntyZFQ6l/5aHhGniEO2uvQQW9AE3rpZXvC/Fy93Tiw1
LZ9fk8Ldo7cT8ndDfZ62nWmLX0WOv0mGcuDeRCb5/mRrsMEkbQQ+wyR6oMEER1UCr1al1sBIZ71u
bBKBZLLC4CAEsoysJwR/WyX0BaU5ml3zZxLjpjM3UGJrPCeZ4XT+CdB5vCmWW6uzbEvz9c7KMZW6
tO8zhO7rlDcWr7Gg/odfBUzOX3c7tn4jCDU3EbTMdjOT4lcV444Jme3h4PhvaxbizGhUZKsCLpE9
TPQrHvjGoqUmDWyeYfEpEAqqR7yo9T8AhccBLmDdIMZLVxSkxudXO5xI+xt+L/FF+uffoIt+tuOD
APiGIkipfQ/6FL+M+Fn5U4LapGmXhRCLL8KnmrnkNj1lMqGOo8bwrZrRY2FUZC5ZyijyZnoh5jhD
ie4VpOUU6c2fXaG8nCwtNu5SA343MI5qLofG9H1m5WbEgvzRm/rTXhGiVcc6dC/bNsNJJd7t4dI8
ii5wte1wwGGSbUZQ7SF4Asd1w/ZfYoxc2cTaCWp1tYgajymSe25h4dnPwGE/CXLzkBsYyCOkqb6l
NztRBd1STCbR7yBbgBGmcxJBxchyJJovpAk/91XfueCYlAEnUZErbf+Y+BsD/a9ZWMxTJTVqlq4w
fKi0ke80lS5oGTp1om342+ACCTMDJOXJKXAvS1YfM2NseWqeB+uVAxrcVi8r3OVloTN3qRXOOSLi
X9nFD2FeG3JhR31D8Mugg4vtgZvQGtYksW09UsBmDb6XfpGpIlqgGroflI60vqDsdg//dNrXSl9f
DpImTqP9oISEY1AMq0YS/rbiwWCdVRP+vH1Mc6XwxDVcg/ObhhFfv/MYohr+kbWXQgeuE0ZMg+Rg
046YRJbai+PCWYJgEc22ripMQl42DvyFp8Xyu/f2MZTNacn1taakshEufgVkf+O4g4rEvzUBd6sk
CF6GRfQ2hv8RlqmE9Z6KxOreTE4fZXB0Y1iOUVYuNZaoX0yr/oIsC+W1frv1faieqbsAlMg4yBxd
85/A7yO3iiju35jsPV9FX86YNBs0zdphyUKW7+M4icCspV/tTEGw793vNRvZhdWIdhwpbx5pbNg6
e85tp5VQJezfpSSvmg9F9i8DIFvNb99YuRd22xcuuzuE0e6BaKoEteUlZCDjhB+/1Ulg65b6L35t
z8vP9rFbrgkipJIVWGY1JeKjfq7WVnG3oTH9V8pJCLZUEP1Ax18ZM/B/MK3xay9YWDfpdT0s3/bY
NKUTWb6eUbzIVIYt+81kzFHRVcpw3abMGC3c1pStyRKv38GC5R6qPd4UBW7n73RLE1OweSPl8osC
xvF4nCgWCWi9mwBRitVkkEEqAkhMzp4UXH7Fw/DSgK+YYePonxB4l99quh3rD0Lds0aLWWAXwDGz
rYo8LUldlU4F5r4ANvAkCP63jqo6BbQHbHKh15eMJRWhrQa/V+x+H1411+f6QGCwYlBeKbO0dMAh
f+rb8eAMMARe6/UAC3+PxCIyH3EekzC6AhC+meyto8JdpF8/ePQGkew73v8EhbGc7RRVKP5fhaGL
V13u2PuPM3MzAleyI+ysiNIjmDfdxemOlxn1sSQPG2FU5wWIL+4Tn5fNdk/LTkiHOI6YWv6GMzNT
S5OMkkaDxdztWRZZXbhE+paMKwMExn90NZBVRh9MItdLpM+EgI67ChNcc+1OI19R8FzH3qEYB+mZ
zsSbeYBk8qC7HuGuA/XNQuy0bSJvQthHVMLkue5rA2zF5ZKw/BJAzaghoNumhVUYMxrXCa7PnB81
lTXGSsxXgkubVXVMeO1oiUUChrsX8mT3KrgLlqhKdVlQdSfL5fLUDBKLD0aah2gi4iSKfOoc2Lvg
4wKsYuS7aJ7FtQnEH3YDw5vSlQ60Z5EWaNERCL+YjoiPLGOgBOxui/qzMSHD0FbGubsEowUPm3zg
FzBDJlUb68vhSX07LNEkmjJV3zIMx4f31Z9h8z/RIG7moNAvyd84ttigiZhs+J9LNAbduzaX1UVw
K/uvYjXuOx5Q+OxthaKSvK5rCguCFQ+B7HCrSrVc1a1wl79yEN2aklQ9kTun827uyHdjBFVcIEul
5deaOWt0vxvLDqsnuZWaWqE1Fr3A9Yp5d6VpfJbwQUBpahCTNZasHshp1CVPXSZni3+Mh3VTZF8f
4xzBKWjQse0KxIl7ARcDAL9ZyFbAo2zLAUSJkLLBRT05gl7zAgyCpqNvbE+pQW3a+RqfWr335gFG
TC8nrsvOizhdYnuWKJj63EbUHo1LMJDlFdoVH4KrNZS/FM2hwFoLLm+wOcHgIhR97ELYpeCPxWPO
OYBT3Q8TL9244POMlPIonGJ68BRW+oOVVii6ICSqNp60SANgBqOFop1sjdlWlH1I66YBN+R5MFaM
SjwapYGirwsI8UU5BnIk9afaLvrTo2lUVYwy4vq40cMEfp9zji2/l84NVxWYvSHDuEBOfzDJFdj9
Bwb6RJIFdEZBFuTfdZi/a4+tm2TeUB+pWXGUTd5DkgY6zSuosMM7ruXKI2n/jUfOr1zy9lpXi436
3qI1iQTdH3sTD6mAzTpLUsUfMb04UPLu3qXUUNiID3pa5ZNNiSbrEybPyiX76Q5vs3VnFOJKtMx2
5TN3rsUNxY66FbsoDkcCVa3LYFxobZm6m2WtAVfpMAYdlCw6py/rgME6j2dbC1JYBB7kTSV2Pniw
oB7FE1RRDcUbRmFKT6KRYrsIIcUnUTP2bXCJK7CRgsvuL4YipcQN/IJGIhhf7ks1SFrwM5xAILrv
qv6F6wHC2x3CJ+1kZZCbwIGXq2CCPoFNZXStHg8Cc/JJdOT/9Ws27QG32EpIjOWsS4klKqcEmM/U
JRrZ6vRLFrE26LBYttsb278HqdEnc9iUbVoMWW4EY1WeFZH8hkbg/3C03R8yazjY9APNsc/T5Nje
vwLfR3oFABz4nNF5PY1AZ1v9uADboxX8MUaphGC7XFlg7A23CvRhMNT2mWk2hyHeTG4oqrH7wpEN
y9kTaoJ0uHyfPWteuoBc4jO9zwJ8jwwGNNxRuDCzBd7GS3DDB7y93+oJ+fgsjdtZUxW+Nj8ZVTBZ
y12RMrxq2oNoZagE4Jnqc3GGzZCYr9Uoumyp6rF9TEqH/gWHopC1zVkw9EB2dA16lMJjxgtXfDYa
fWBp4aOLeAcvvmaay772FCX/ph6NI3OL9+bAQHocwZaoGHGqHbwHVNxOKyXWQVjENobVWnUXBaVv
pw6Tz9WyAaIuByg5huRWGPqPYvpzAA1Lead7Z9veyh8yOsbPE56CLLzjJ2HnxkENvafJnTmDaJiO
03i5e4tmPy8xJqKQmCNnaSujCG2OSiZvipAbnQjkVRuLjOLhVI+xwvT6AECHLqZLgqnTpbATc+Qb
SsGOKXGda/kJrCHr7fqd40XioeWAbq3BNDHYKD72q2jqpGMlRh9tYpyMAqqn2h/e9GV0S1wVQ1ux
RVOBHeMMpb6OP/dWBNlIRBararaEJ1o5lT2/reO6BT+oiDJ/DN/VfRPvU6E4knrnjX2QCsHjAI+U
64qVwAgF0lmWMrXEKXtrldQiFWrtgRYc42qKb0fx4+Y5fk96EOTLewITfsLLG0mJtyWZilHpM/3T
cNyInvSSfCK9GGOicJ1ZqlvBeG43+8mrPqVmxW+MZNYnLbwFU1+0usdM7ZKmtlsEwKzoR0tvmz3p
tI2P5R1J8XtHZsbEOB1PZUfYDiKp6gnuwK/PJczfBisEistgODkZgrrMvHo3cD9LOiWtJ6FzQNPg
O1ByXAWHoaiIdzP02aDQJTJe93RSES7oRajX7zNBktuuHTz7qkxTMT4cN93/2L72O3vuRcLxQUug
Dgayf2wZnxcM/8qnMPGJp483tfuyrtAmw8jXi+CnHL4woRROScw6BpS1ndZBXKtq7sYbxPfRJevI
bZ1uAaRBN9BDi1Wyi6/nYKoXJt/ZPaxMXREApAZ18KKG2taxHwh2vTwADBZJJ1LgP1IQN147LDaM
CA/vWmVY7tD6tBBkF7VKhF9Dos1UVKPBmVcT5+6Sze6sG+wSMpLLoyx1I5nSk5ZWdfelS0qeAOC0
MhrrNTBaN6pqtEct6yHDeYwPetGhWDO2z11cHKqZbcQJMPjhWpxr6/MjIwZeFPfi0TpnrVC0pyop
i+P+oWDMGQ3GsgRupLI5OjAgSWiRPh9ppo3YYUuHC8NZkZSW3KZatZXVemNErQUmTPUHZmT/fWVL
6ABtupz9WDvxj+fPVS4PqhO2iIS5wdwIMXrH66VytGJycX4hR0bA4IfmHFr4yzgl2c8XK/37gN1p
Jpek7wl+jr7nOt1KMmZOJR+DVrG9kXM7cNswJPPhMuLue5wqPuYUdoYBbrawiB8XKQ2Cr4PIDzuI
HjX7oQ0lj1icP7S9oUyNesWpJKXLaVq8hOaUyhXbzAN2uGw6T27cRwkWKmN8DbPZYq21NpzCZC+N
9YIMPE7kNEnuBqipYzRiyWHnB/qtME1EltFm0h/IXXZB0c1t5RrPaU7kQi6KT20WkVh9C+mAfvqp
k20FnwzCKFKTCt29sRmpMxB+UEPE2DxdhzBBiJ2CXb1Ge3ySbxi4NoWN5ZnT6dUPT439pSbd0kVY
B5WHJ6ASHbzDVBSezQm6qyyq811AA1Wn+n8pSrZp1KxUmLt5HhPN/Qz51q7cceP5numnd+4+AN/X
LBt23fkmgcPZLP1nkVtJ+3Jfu2hf1W0wueOb640pSigcE8WpuafQI2XqZw4RwyCqvtZLJFOKqtYx
H/q+MDY50+T12gJ/IaTLiUdWMiRtXPpAPSmonGpDSqnPf0h3TOhHtEgNd+W+DYcXxiYRTvX65vHe
TIiWMh45Qz5YuIwc7qzipBiC/oSeNKukDfuZnQznVnHEQCK6w/tRV+sJmWjuUbRv4Tb01MxNvCes
9n/N4eZUmSG6gJns9BuV0MoDG9G1X5wDMqyG7UC01j7zHECnMnhZvtgfHyqXUtpJABg1PoUcDL2c
Ef5UVO6c4QqjYLSvqd72M5Y52oF7NxzEIHgfl23df+We/ce21ASg4898iWcPn2dT6lxvrf8ek5g/
wd2c5JpuKNhcXasE4LNQJpqweyV4r8dnyh+Itp9VoixMHnZjH0NaUn600ZIWO7HF4cQyXWVnRlO2
7CdyPOejgubzgMQNdC0pYfAao+qXmyq/8YQrkiVw9c2piiZMvphMYYAcxJ3LTbzfY7Hk2v9UDgXC
8+7CtLtxM+YwjwQuSlorJyF+ZR5TQ1LenFArKWEoWvNEY6IUcXfXvltSHa2d9OohnllaoNOh8HmC
dHPtqVHDkJ9vPcGGF+xZ6bE/NEXkV6LbQ7ksytRmZTWS61/34e9eItK3PfdOF5HSnjbxOQYI/KId
nT8HHNFafYUmBWV/p4Q0QqU7uqMv8Kb5yMuzzl8mW845q9rFVRxMNVl0K2+fM5txm44zu2j5aXv3
VFv8JBTC3psq9BkBMfwUmIXmpa682DFBRcuiIyioaiMVy7bJcjLSpMpWmDlfGh4sn5lsWwdZ6GAo
lKv5oQn6meho7fVNbLhzxDA+8Xk0nZyE1vuV7H92IZc1IbNeuCPBmRizLBGWoMVO1NlaXjRZ2k0r
qwxO01XrnYbkKpihE1sXvnpSjXNB6Cpk5qNw/3+I2CrwXWpfZ3ArJ60wpNzmtEfwIayhJVyAJ/gU
Hd9k3Xbh98lq1CKfTqDWBkLQ1KBs7HxlTta2KDAVyHPVSxydhPYgb8BeSa8uzKyXPGXq4Sm7ZUTp
E5H8wgnnizFZUEn8H7QTfdbgmOq9HoQPT5JOBfCuozK7vEcgPeRBBrBcpxz1HkEaKejTrtLmn2fs
iBfrsq821/aIQ0uNPdCSpp5MPFlWPbXgM9lPd5H03psUZP/MJo4Fme79MfGkpry0MoxzEF8niM80
TIZl6F7wXKk7ZoJZ0Qe8iykeh7NT6IsVwG3Kijpu+qOyZ+lEA3G7GfxuSO/WEeCygZ+lfL8LzRb9
IKKnhyNcfWk/XxWcepYQrGrWwx/QRmivIKJkFHL47vWFQDZMTnjB0tWwod515/i7+sFBtpfid+ML
8lBtkJxYIMgF34jLwSuUIjT5FIfkx3VMJDId4espuoAqRSb6LaGY1Us3vSXba5eRXzM5tS65U3rx
JIsfkkMzIH34FEr2+bZliqQMTqf6zQZ49R1ve2yS+WwgiN0M5HxwRKjf11kuuBmQd+UBZltXfX+P
GYLpqfmJy/RUBihXUUdr7pHTlgUQQOz5p3xMtrdL1sv0R3k4jvDzOkGkdd04w5xUGIwr5FqJPdul
7s5VCLir4Qj2vKnO7ABnPY4U2mrPQcNLwTY26bvhc6suITRPh+51ZsFYrYcm8RqfNCSeK96oKAqs
EmB86y8lOpqr9VrZHuNJVI5pPq14YubcJ4QJ3ju28EGIAn3J2ize8hX5WuBXfe/egjnibYOuWKgM
Z+wVjTYalnBFuh3ujkiTbT/EQCnaTrKU08nE5uLl7WvPC815m6TFP4zvA66COPypfLC9hSHmPToF
j4ENHLDcK0RcUoqonKLPO4SdPXxQLyBigyZPUurv9m5oO7/5fFc7uQqvkk36pxq8J9UA6aqGE59M
HU1M/tJR1BCluuxv3az/7BJv9MvAc/LaOmRHis6+lM2BcERr95WPqvsw72s60WQR5+5IqXcju7hg
BRSQs169VgGo4F7SClIhjQX0gL3+aK343iTXbmh29Kl/dBfJkORFVRoHAa6SQ+mrtj0Qn9guOqJ5
/Nr20PqTNQagFV5dVFTDdva0FEwAL19z9OMTOBCV8kzCiFipY8KH4DO0cjFruEpv4SUELKkK5irI
6ABH6w5Fhn9BBbOGFYrT/UjvS4LrW6cKbHvGmzoJt0vwqQhSKKxkRaVsIcd1q2+nc4f/h1C+Msk/
x5/7BHGLCUmYHx4DDMVgDAkwL8cpG3H7a1mM1Eo5ccigdpPyvCqEZFnsFkf1G3gr21fORK4mm6WQ
5AsFR1Fryp/1tLJrt8y5wSo5mTVkU/nFSEfwOzrJX1jJSjS57WwEBlbskXEgfPGt7nKeXAJ4ldKL
buTxd/B7x1EfswigQsMglefFapA7nxtg8JFpB5cQsNg4YGErVpWoVbegTmYqQ37TdRh98Yrlprf4
GWsCCHHrpEu3g/+a8uO5poIN4WpLtdqIwKZq6+DW+5ytT/yff+3+zhRQOKwHMtBShZFxT2nkyHux
yCejEPK5DNA+m6pBvTt/HWE8LFdOt2Hk7fOGPwKL7ZqMDvFYAjq7GxZI/sEfznR8EabEM/4XOpQQ
p+bYmth622tocEFyPJY/X4T+d1Dq8XPM/CRx8Tr8A3bBv7FEuGhdJMNEsHe56yrsKcuTvCuHszNj
ojOU+U3pwJGNWzYTj6wAFhN5L1uzYF3ILV+lNphDU+LwRsobdz0ucNsf/sD4XQXbs9Fd9crQEVZl
xPH0bLq/JoUyToltTnwpDwrZpfb2F8O4CG1FqQC2NOfSlgnknqE6NwWifrjpCFtXBAOscv6GpYOg
0vQ+r7a5F+XTae8xnXeY3YuKFEDqX+W6h5BsWyJg1watjHiOUGVQeBJJ/ng5S13O37tMwXrOHz9m
TCJpDAwbfgHLZPf9zjCvmt8P+2NZCB3dFO45uj6da2pofcD1ev5HdnEvC8KgG/NN5ym0aux0RTcl
pTiq9tHgDVk/3+lO0aFMUUorprnB/j7SRd/fHyugAKB9ch0tMHXq/CT4T0UMh2IPItrZ/dunRniN
aBlhizR7tW1SwqqO+gq1Zd1GD+QHDsHsWxC4neASOdQKblH1fCoC8G0k15en1jGFxtlwY59ediCI
mwin+BojcCUhzxAS8ypBYpVD0lerrYhZdBvnl/76EFPfgDZ2V7g3p9GocdFLAywYjF6MdywIQl3y
OXRS3hRxw4ERdLeUaQYBB9rgSolOFQL77C/xOg73rWl5jUMjBYUULGVeXKkZqYS5ibaHzPqbmw10
rgS1fd2fUPjH+5gh/Xhw7Bs9PFXjliRKEc12ENDCmEtvg+paj1Zxij4n+EKKmLsAqoWTSR+ChbIR
N8jMiez5ZADFbBaWzYqwz7nTWT2piZ+XNlRfuq2ZG1KO4C0AR/0WksbyVAci8Cjk1xt2miE6+Ug2
pSQwPI7BGp2YRO/2amf8qFGHdG1Gp9CEA6uDtE2V9LTSN2KbW1nCwmpvZ2TF4q2Oe4yc8aikSYUN
Sb3a1CMEDc0vmNvMwNaDgR5FT6q/Mrbi3C+ELuL38svKmag5S29P9e+UCeAS65VNagsSxxLUFeXo
57f1btILbqHfGH1uNd5iUEgQT6v90owA65lh4smt6lIK/XZpe9f14X8vSQHtlxF0+TRcRE8YApDr
VkgB04uXmJ+CTKNFRYi0nghBpouJisSMu6XkQgyHUew5OkepyDjbBmLoNpgXl7kzgNjNGLAW1QoZ
Yz2bvtYObnaKVgsjVXLUhtV51Ov4m1U0CTXkjiG7HfzeGFFvgd/sApnB2F3VW1XKV0oa+IhY4V+l
KATKFbhhDRmOlxN7LHFGkaXNtVFjUKM59qqltRVeuUGAKnOSCItev5LwwC0UeFLn9hXJagVvzSN/
+e8TlzANfmJOeycfH10ym61z6oEQnii0b2lrM9b7iuGTZDZnH2Th01OOe1UHmLi9+HWSBuo6GCaP
WT7kQeJt2qM423FMnrEitPPaT9zQGbYyr/9EZ3aI+rYeK0yeiogmOtRYvPtr3aTb72HmV0JCDT5d
KN1T2TaJ6RM6Rqbbgos17/+ujFnU0Gbj67XjR5ZCm/EJ3urIeWZcDl1Vtwgz6LOgWQI3csucZZXu
x0tT1L2NfwlaCZJOYwjK/pgAxJeAC8NSiiO3T8mI+RXgmeipiRnXHQ2sZrEAPX9Oe9bUSD83yw50
+GmNAiayRpuvfDEQTUhCdKMTxkT45fmV3hablfZJTBepVf5MHcHcnVwyd2Do1gG7RwFOgZruqiJ9
3Jdz3a+0NqcRlkpbN80Dc9QkxQWwzbRWRVsjJX9Hn21WPWA+bSswOC2/KXJFdyC1qPqD1blKjVK6
9kOKnP28flIdDgdEjjUPxZgmMYzZf+6Z2N92Y74vIPoPiciuQ2Ne84ejWktRfbxSjPiw2+aVP4oP
4TYJ0CFUwZbMJeyvmN8etpzOlVKd7/fYQy/AjOi8h3ryC72FYPYHVNZwr0Zz4TWflJrLx5eAwG4O
7SJRXg4bUqtHYPeOoeA59wS1E2GS1qjO1/1oTkSV/Uu2zUVN38pntFUGf/5g82CZngaRZvlu50J1
GjrYd+MANo2sa15Xjv0b4OEme4J2RWQDmweaSTBw6Kccrn+Y4aaNuceQ2NC2Jlm46BH+30n4uSFY
daXu8lC3c3YUWWBwp5gJ/BtEHoJSad728vMhJFDlsaRs7HzPsxASsvlQ3vBdJcsPYnig/CDE6LHx
C0fk61fycxrRzh/kTzEt00hDcni9E7/H1xWaaEFEvBZGJW5jjBHJ9k1unWelzYDavT0j0w1L9gv5
Xw6+/sXTKHQOWkGU66sI1TMIUX7PD62EAZfJbIKIoqnyq3RznRqO1+D5dj4cvq0h3sk1l3nPLHiU
XDXyqDRma5XG2C3iby/6ivrS5rfqwkDa7TQZW6y55jxTOZ4ACwPyXukpU3O3LK8/lO1diNEMUS7C
vpdtGfVzIWN77c9exK+tydl680nRmWjQOBSr7KkPv9ZWHvKboDaoJIufznl7nep5vhjM9fjVgg0V
7kl3RSo2BWRjAXYNZOSBWdlS9GWAk9BJR7Pf84BMKjNylH0Ow0uXzkFK92Fn6AI+EAp3Xtagg/bE
I/ovkOtwfi3m2YO//ma5fAL43Z4OhWNamjEtauJv0iqHXNi9mFvoxFMNGBUhD37yxvCvMoPt7Pot
neI9oXPhMJEcmjB3CT0Rx5Daylp1EIaus3hJW1MU9aTCYlbgFh1NFqK3khLH+kHbXaqEXF6ESJkD
NQPTAncHq5/aEQbdnyr6DyglfyQu/0sMCcve7/h49Iz7+jl1k7cMVa9ez/xWZUPElKPnl9k4yq2S
RIaJ9f0B6D8VvUAH2WH0rK8MUfXgmhB7fS50XwXuleDsWi40WO76J3U3+oiwjGcBDK52RNyrvDzj
o3D/PbIrMMoFTBH8i7n6vEDhNP80Lyw+QTC+H3KzXka2gZiT2tRGANwPAfHNZhwhRpSxzXBmEQ4u
psbruWRlRkSuDrvN1mOBbGxD/IC8LsNPTbQ7Yzlor/CwPBO38Xoyae9+9O2n29mc/Nze0VtubqzV
qktPSdnynnsBal3vqZX+49Tg4+y6xLmcxEfTmkU+XHb7DHI7waDmDa64tEm7OEiPaiebHFaA6M77
gi6uSZK+mmSDzmuh9OoutfCgY6sR4fBTLtKu67LK71n6xRHEnmmaO2UHVAErQc/+KLmeSheMrwBJ
komrZdUeivMBmCdFrb92uK3NQCYBhJrMjj62GaemJ9kGRVUsVffQ6lSKH+FPeBgAoXYdJTW9fn1u
XB9R9n0v4eSDB3lP/vUJyGV6CKOP/UZBLjT4/Uu9s3hVoYB9ljgjTb0eDwm02CTio7wGIggVQdZe
tuH8ctbAzSok657QX126yPqRkpoV2tMG65UcD67HESLo8TRTn6lIiX1wJtLmb58vG6xQ6pLXYP4u
tvdQRciCrkN63LggF7cR050XnYb/OwHRcrpkux8JRU2g/BZTsWk57oL4j6Azu83eu4/0va3cUQ4t
9lc3v+9TXPxINflqKyT566RkbUFvyg/tIdaJPgc2gt7hLnyivsQ31iQnyyOJHloqgiLaP+u7g16a
wG6DkviuyAcKJ9alEzTHgFVAMfZCcyS23idD+sDPhDC7QCuEeWjwuKLwPbW3CmCLOH6DfwyltmZm
S5qMhVjT3WuUVUfupVI4kDSI6jkf/ZVYtBjykFT47kG0sVbFPVRo2auCA09SuJWXbtkiw+6dOQzT
3C+Tb71IHf7bEOSU1xudWG35wePA6a7aIf3u5MySBOvF/PSw2jLR0cudaVI3i6qCFJ0kY8+X7BTM
bmeR+e89qmS3FHJKAVChtw+03C61ny+4rnAA+FeHdE1s43eFx/vi/dXocg3y1omTEoj4k7NPVBTJ
Yaue2hfm07p+6VGzAAR7QgnKoyIQKC/Sm/DkKhi5UhwxMbcPlD864oavzVV1gJh/Hbg3lcqlfur6
LB0q4q40RSQMLuD1Oonjkwa7lmhl1akJPw0lUhJVy7VjVLsKJHf86nE5jhNVG4LdGMYyU5RPfFzS
JXDFqo836VtLEzowW1qF0utHt+u46NE3iW8ozopCpw1NiR5VjAITpMD6CIaYdyzAb21pFxyVKolW
rjJusFPITwjjQKov6joSWPoKz0kGGlTAEVUjPMlDE6SsYgBIHNRkNGDU2lAU2AcdvQcVoJdKAVMR
eCFJhUs1sYwZIsDjJiHUepgkfdQv1WKn7J/B1qwWUdD73xFxyqw6KIAlZquvHq4dr3NahpRoBJK/
JWIEzEBUwFi+ileYz4Fh2rY02X0kN5FsWttS8+O/kQxJkTLxcOQ+bFrg8s9FF3ysyOiaAz9Nniqs
G4Co/qX3z3qqOmUvYSosiZ+2rm7cOoQ5WOqe/qGjwnElGwKN24oxjbI8G1DOP1uQbqeQbJuoKt8v
x2I4iNqySh4/SdEh9Feyn4o2HmJ+AskLQ3gkLj2lkfknvdyPRD9jSsMHqj/GsUi1i7m/VoSa0Bsr
lrU2+XAkVqy/MrR9iWzReR2pZEL9Id16koCNCebf8gRdXmLcgeVruFfdGPE6Io72San80Oic0FSY
PVrV24iX921jurdiJz7uBmXNfWo6+mCBdrYyuuiTafq8nVKObGwmHwIuRUtZzSTVYXrRHYCI4E3+
UjdhTV7NmK/30u0zhMsdUUZRNdQvq0RTj5fhTA+AhLgAvy1ox9ImSi6tbq+U1MamM9c9QK2wYIgY
tSbTSCDm8CzT08MlHhoFawzEUsUmL/TPL3NvTy6l2nTZSUJx6zbpm1Cw7QV6noVCBlv8Z/ToogF4
5c6zgee1LkR5VjrC2U0XiwP4mx0yfWYcuyCJH67xLVWXEmBiHvUvoCnynPTjQk5xClfRbEjkfe4H
jxtKJ1uR36yITsX7FsZupc6e2rNf9Sqzi/iAwDVLFszM/VQgfMjyAjPuWfOHI7wARShhaJYVx2dE
wkyTUlPTT3XRdC+yN8qzdVdA0qgULi06Rr8fl/zCVruI9yxwHT5OvTmkqmYgUOtbEjuqm/ox1wdS
/uj30SwG3FWycBnDRYPihTUr/CTXLYR7nm1lul9dlRrK8o2VTH9j585xlGHDOOD5t7vkQP4lpbLn
mRkpsVwJa0cqhv0fQ3vJCjNuo3TWdWzSwvJD0Y/HR1gb9Nqs7wA7ntfHkHc5/Gx4OLUTztKFr4gV
f47yahujgK/p6GqPtSuEsYwwvvDeM3lc88/pCGg8fXobVPF7laxCu5tW2Sa82TzBtW/TOfHiKXIT
WUfLr+dRX8zEORMbarRkL0//nQHPONvQW6PDcaJMlCCLJQCxH6dAgFMrqtiB5DdgWsJQctDuubro
Bm5u8wRNQq6y47Lnk1T1UbHWCTVgGOJ5vEQGAV3wy/cWA7Wv99uG/NvlGfaMntHwGD1tzXCQksMq
JGGIVswf7USJWghukUyWLG0FTBc5nt/vygmG0wF5ShDFy+Eh7XqbBtXfku2hPhi52xPTEdwaWsp0
RA2w8P+sdKoxtqJvBFYFgo/ZXz9f3bVOn8zHDhacYbJEOhG1efUbuHy99tV3EPeuCJYHiweG4XbO
YlSAFFrsPncjmLMckMrsEDaecVGESeSYF1LNcXE4ZE21sA8ugE8egPCjSHlUeF7QseGo5F5efOJm
LkqbTP3hpVS7vjk/fcC+O792xQJYnXCQdfcgeeoEoF7/hHpxdV0n63/j7OVyWK5K+LIgLBt0Qzda
MU1mFtB5EhImF0IZfnm0Fz1driXeai0T9RCbo0RAup9/V47IXG/t8YS084x77MPKprfGDjbRVM1o
uoqLg1FY3HKQSGDMhG0A/3uGHKnnMZwrFGP2PMOtf04IU7KhuegP4A1qJe6Qqt66uqdGkZdri+aF
jU4c9BmayXexLO/+RreCHbgenXzM2SfIH78iw/MrsUWLPpPAEQQOK1ZYmi/1NdKiTWP3Q546HDtA
/XTzh3Vc8xYpyVxjcaaCUEWojyKWXPCMkK6DH3bj8v/gl3Qt2oJCJthcrttLZUP3Fh27JYbMB7wb
8IaPpHxnsvlFXIAIhtjMJCBiWkNvB06GKBGxSrtJEWrg3OcBxXVskGejwjQWh2iQ23kjn71KDysX
VoV1wNFr1xo8qENPZMCXu6UN2FY//HEDM/PbFSIQRPUnkA29XI2J/mIBdfQRc+Gwm2NY8j1NSVqI
YOdrg8DK1Vc3QOwpKZOE9g2MwJjVNqSsivPxpv6CTfqC1MkaZSgyTnYW7EseqUjjUBm5SHogExFv
umIJ7kOobRec9VUK0GRWaBPU/jTh1XQGLqnuLUTJD27wIUK2IFjMZGhe6qiZ5ME02yFTI6I6Ud00
cY9QNAkxm0hGfOczDI7RQT5n7dx1cUEn4fF4rcF7/ezVdFAN9GWwQXzaf1rwJ14U1I7kHnZ21pFl
n72C5HSipHPkbD9ioc45lWsW27yoaA2aVZCQguUp6Jlqlo43tuDNyN2NfBmRc8j8F9g1vG9hgbze
04PbdBy6fEvnFfEcqv2n/nului7x7GcIUDUosH0WE4VIWoOTXsHO/weALY0M70WMxuC6meQBj6Mp
w3KUSqKY7HomCRBNUdsTT+kwdO//rXsuwb78+BQMsxw7OqBoWuF8bzYpzKJl8BCjnMkQTmyUJfeU
qxsCDF5zN/89AWjxBPJRpIjMEdl3Q3YKHpiaRlJ4jDIDQZcptXp8cyHA5Xubb2gnnm3JNwtRIg7N
qNGH6eN89VGkb0cpsRObTYwOuf4mba2lTl5HoG7kOFd4XSeNC6gqLGHflvOgidF2jI+BX2Ho078g
yNXCf8e4mI6mlyQYtwtQ2yWw9ZpD7DgcBNvn9ShE5JSIDp8p3EsrUp64pgrhq/KXmRTUr1nx7Vgj
MpuozCGBh7GciyYxExr0LsHmjZq/nvOqFElpk73VVjL3ZkpJ/4vWqBouENxxFJRU6QsHtX0jkzOX
HcmrDUvvJ5zIjGp3PQ9X1rzSb2bsMv7qJHvi+B0bcRtbJQJDwEo1cRFT2NYNJRPSwWF+cYg/VWR9
ysOWVyBEcboBFkbXyQfud4o8ifScp7iqqQ/i2zKzjDvejqxbT72gYA/tuXZTePA7edYM2P6xww7m
4m0i9ilJ5q1pHS/Wu2/9ckO3MOs2L5yOajWLFtrjfy4fbhCFEGeABEtJsnA0H2QnZSxN4blnebv6
qhDlcKGZwZxUQrKP01wv6HVHr4wD7+CWr5BYFy8A9k0t7fSHhSILo5fjqmeajP1aDPQ9JAbDHb8I
2TuNMQqWC9kzzUeEjT4pWuqR9CdC7Qa3OwOnIr8z3OT57M8jwjvtJmnN+BuGqv6WwJEJlNfQca8l
1Jy8+CS8mVCCsmsejtuWXx1PG1KljFP8BCQdEU1i3N7xFsg20ZzrmJf6HfA4VqEa0KUQCPuSVEGt
IaKFO6k3ZvgXpJ6nxiIy/XaNdG49VxqXLcjXeke3LO40COZwsTFWB2BcZAEcYlIfriRhGISeIs8z
dg0dZ8RDOXgRI48uGJTWCwlR7risvflxzuGTR7o3liDn/kFVFTG05RIa2EwxhGh3H2yDz6Sdhuvp
TTz/ppSEHu7r98GHeY9TuzRg1rNpVgbtwufmZoXGPMnXxF6g5OjpTQdgTTd7WuTpyDDFCpwujz8l
4qR7isuGL7SrbhAvkb6102lQnKF+Yl5DF3mLXh4vYatJz2ibvHhWSMz+4/Ek8NQkA4zvop5XfGHt
GA0tyKwwFXiObBYoYrRd2hWSTl3uod1O2H/CrUsd1OYWqvFH1fZaZ6cxZbuzigJ76ntXmEpUfWX1
DWIseiPVXz5zmsD2owwR99IRRaFC/KOK1LcfWSMW2GqKZtYIB9R5+kX3rWBbgS1QJPeKyNJmQq+U
mq1ojQ+yhJabBHCOxhb4NCDHMI5I1FRYsGOO834/oid/xtQAwjYAfOEaUvyD7koAmASAzGzNtiem
vFfn2KLFtyN0h3l2E0d3P17Fam9nB8j+qTKJzn6txOdm/i9Y+doFe5DO8ep37gJnoiSolpMgEpva
QVdebKfRR6kSTLnZRfkGIBqud5GTafxpj7Rny37bcq8OuNKwcv4RX4KGFkNufJSUcT9ySVlh+ZVe
duEg3y2pdpGWOG6bS7uGYm0YRe1R5+jij3TDKbDBG6Cl+aab8uIC8L6GPJ29ihNk/aHkHsjl43WC
LqhXhVlZEtDMM/vXyCvPZXyrASbY+s86nK2KCt4ycs6vNSfZaGc+yDUtQ9UR/8qHgLbsHWDC6VrF
Xf5ZlwRs9O6sz6y2xJWDPePkSA8HIsITo7TC6jtAsw7vFB5pHesxPIsDtS0PcvS6GbJF0lwYOSn2
ij3nXqTV2zqGbsHvYAHsoSkQ4SRIL4C2EjuR0OEfdSDpn8GQr7tRN5uuP5H9BNucuJNLM1KtMKdz
j04NY/WcHyLtmO3Y207MXkBvDfoaED6/L1r7AUq8pOBFRjYr4+rmD8NLRdwxekZSiigYE5aQNFiA
/l3V9pAB0L5+MYgB2AafvOaY8xWBgWz07I22sCi0fPHJoDrN7MjQDKHVFrrtlKSm9pVa0YqvBd6Y
bKWoQpGsJtkiOu17w5qSAWItrNhcCtxF1PgHGSv8eIcLYncvlkqbIOmMLTF3tX0sS51WeAjzUhZ6
DWf2KXHpv+p1s65oSC3993HozD2Pod/PmDH6Xq5mWeGXrFMGvKldMp8tm515MOiX6jl+5eFr8wEu
mwiT0b0eAva8abqAdtKlT9WifHRawX5KjabDxFjLkqD9eSqNsyHsiA6NOyAr8sT5dIK/KcXKMvGa
F8PQYa3vM+m+xBVRlyJuZ6qPyiFX62X2fz6U+06AlcXrea9FNrQES4aASYSSP1kNNG6zVlKAtpnm
A8nrLeQHL0irDMGMBEZEqv5dgMqSN2G+Rkokr6gW844hmza+byeOeL5NZQM7c5clFLswi8j2LWHK
RaEuULkw3Ax71Jg+It9OJwaOaxWYVQZqt0r6mnClBj7RlSfoF4fQvCZ6PTl4mAURjGMUmdsKjvi/
6BmLiy1X816NImLA42uRNhrZt6gwHDNxVAvj0krYZIupudcRkA8j3VagQ6IuD6mDV8YhWJAKIeHo
I1zCRcwGcXIRhvKuUUMJtAi0WRNU3EyjE1YPPPexO6d7zlvM6ybBh1abJLW8vSsTF6MV/DDzxMWr
1pUrDoQZcwi5gBsR4z2hZ2R2ypxkkXRxM0KcHEsb0YL/QlV0i0K6LzEeE5H+2Xmb23lUcbo5Ti+A
lsbTuJJhPfLUBYswW1OMp1kKzaZss/Lm854faTsTqtG4krE9oxeB7DJlbsDbGZGOcc5k1ZmBRtxz
4ICw1pPLntYjk9Hbr36WpGiP4yycElKm5cggbUvat7b6uFEtUY7P1znDSz8OaCMGSRg7aAT8UD/0
OoNvjdHXg+1tH5WxiVAJngEvWQGKrFKmKKssWQcLZPg7gpw59nGxAP/NQhLaZkYDHYzQAE6oC0Ty
RC7FWRE5th2V0q7pv1o1+4vpjPH27C4mw+tEhueZeMAeoLW/5P/U9oYdJb/mlD3+8h3LY/B11c9b
VQLBn8orflzz/A7WfoZt6V6lujvHIU67hWogw4ktwjSQIWI2eQ3gNX4DJYefiWnz8gto6jsvx2ea
WBxDUsYhtgL+Q96KqJ6bsdbghr5XUkiIkU2mVkso1C0GGOpN+ovhYhk3YDOA/DF/DUKdM22RmeHZ
YuScy1tquuQeiBruDgI3pHlAymKkSdpwvdm/d0ZodvPqdiSmWQkasYcJnGgH4a5+ZG2QSuSvphdr
CFzmhEyCvUvlXSG/kDJ+0XtSe0VFC0H4CVjluUFkup6GH1421igzLIEeoNcSByAK7iv5/Zvs9ipr
HVIjGq6sCOOZZOYQAZ/GuC5NO4PHy0MualHSp8xwYwNOzUTpvg7yGVV7LRuEByjaH7t6qscTxT2Y
tr26wcAiDYU3xyi3Bv9kjpuNxM8eZBRKoss530lMwMsqSAbaozpULmThb4vryhBi5Jg87K7CVpgO
z5SUNWyTy0feV8T+8ECbPb7FRLw+z4Lly/jJO8BPAHX3pc1P+7h+YJDePfZ92lkt6GqQwpSnXa/9
j/ojpW7iidQyZ82rBOP51Pww3DipaMbWibC1H//gSOGEgNM42x7j+Jm36Me91EQq5Gz+iBG+DVOF
cDx72g17EY/SZTvo5g63aZrf9m3x6b6jQU4QZ/5rFboKZLLqKCFrbK+6lSlTSsggkppgrAz15OrD
H5FAUI7DtHS3EuDk4c2nMZn9lYdHqa644yqPWNMsGbMveRmMKI8Q5uTu4A2OTCao5xxGj7INdA0l
vroURfz/LEwioOSj43YgX1BFptGfYpHdgY7rrCwEsGt0pX6BOY17CImC7BD71dl7o7KiguC20TZU
s5ItrAYR+wUI+WgZHE+m1ntMYzUHJvNyGBu7wfORFcgAu3i1l59aWCuGTyHMPgm4EHe+aV1B6FU3
F/186qmYqNiPSoCxb9WzY73KoXzl1/9mfjDXpa3IHA8gT6NrvpOH1vQamlhCGhQk9CV+AHe0jXub
XDl0Kh2H7ypV/rtV9F8U9LBjQZcg8IsZrXfhjSwekKq0JOqfZFM427fzF3kK0AIXQQMOgFnf6yxw
AuJWIqPbrndTq++2lsVLbxOm+ZMkKpAGIJyw2PYbmWKk2Q57XpWLfF1wkGMB9sHzeD/aahvJFXnp
gdTBRHsXavr6r4d/Lq07pyjtlWDUE/+mNKPi7Z7f081463VzhIombibzDS+we+/i1f+KzqA5Zi73
OpP7qHAFaz4t4BszAejrBrRtCbWALFCsC6vpYgKYwnHBaIPnkNPPyU2N7fGcZI6awtrAZgz6K4dC
Ww3C2jQbKxluSc+EOCE4SAjTq6tinFz0wtxjz6i8F36IcQJtzTVSVcqFphml7atZ9Ydr554bvNW0
4Uy+ss43b1UiZASovmZ7vcdlFIIvsbU53sd3BPISo+UPI6hLeDqBMxFKE6JbhpzgB+Qlsz7V08Ws
ZXxRsPyyVBLpnQDxd7ElYSCbjy+s54ob9q/hk7rA+SDK+9aAKcvNEfRTytbMl9BW0mLbGTekr5bB
WBRulUkWaomh9VMQnS2c/ze7HS12Bm3oK3HIY5UH+Gly20SUVfw/5QUuicH8WRGDt7Bq5jwM+p2n
3Fm7JPReA4Z2OFRm+RvBBeV7VwY4O8GoQrHxo3kbK7OWWL7Tnjz97R6LXzs0YJVcMeLq1ZSLn1+Q
yLn+rG9oKpLDIj73sSDIEN6zN+uTfgENBFmb/MGVKxPM1JuTFfDtyIbeNAhR1YVBTFcUnCfnd92o
AO/JV2bsrLEMeIffkMC5u7DyGBNGBo+VT26hyDERzQQwEhMMPNCcuJIll1xw76zJ8dvPC63HW5nf
tH3QC2nBgXSsXxFSnF5DS3hfjaXmwudGYGTpQn4ZjYvHaSqvnxx8qwwdG9egCTS6oHGbW5ERhSiE
JXgnetZziAy8zhKYFgznlDJQzUbA5dj91s7YBujepwdSYea7ZKSpnX/2wFH7ujJ4bKGpyPxY10F9
kXpKhmYbJyIJR+VXNEekcWhfYa4ELRnkKW22PWe+NdIVQbRgwxOcj3DoaS+iNsJquHo9hGefNsO7
3tteneXJmMQLfZVkPOmcLfNYbyk4Ef3e+8UIWazg5L9OWTeCygFJY79Q0aE5KjpmQla3j6Eu2T6S
nV2FU90VZfRrmblkavx4CwkPEFjYiclsvIqd625AC/kYo2zdHld6AqB3D+Ds2T6OH46lV7l9i37P
D1W5SQRxLuMWEN8llTqtSj4GaDmjnybWpMNtVLKZtosgl6z31ZDFYq5aW1m7QZpWhc3JmTAUkE6B
jz4oMlg57+EYLFvvFo0PU5hzLCh4VsOK3wiGVHt+bGZOTWb3NsteNhivlzunK6wujoonPD4g/pyu
BeIhLYX2wYQrBBwSKsou0p+SvnqBYwjyeNSsAwKqQVlp1urFa9mB/wqPv64e7SzTelMjaAI3YAkF
HDYFqI71Vo5ZdV0GyaspvP2gi+MQRbIADKDs1/19brgCxHw7NpoR6aZVKt0a3akuwgPY7/6e2zON
0nKrukCnhgxzJPn/YiTPn1USE7nvAjg2GBM3MubEcQSsjfRymM+15ZewNX+lMcz4uu2m7YE9uO9T
HL3GsN4B1LblFIwwmO13gT1qiZD7NG842EXRzVXmXB40D6dtlyFP1AoGRY2NxBitFmNGt9v/Giv3
3c9vN9gmkhZTC7lyC/Rc6xqWgau53/wazNr0KB5BxeKuxG4n99PDABPWD5vifn/H2cGvc8dOLDK4
nsV2r2Ue9kf7aLaNNZ7v8vRa4VxSxe5/iZBe752aiBn/Eya3ne9BmloqSFmHzRKzKdVU/VKaSHvr
SNvBB/kPxf44N3HeRE1D6SWpdUnmbuw35QoGwhtOLzJyE830XN5uJABSjiaV7NwmPxDsYM+FH+Nt
9UAMcFUtT94k+upTse/w/QrOBSzrTJtGCYZ0mRY+AaMwT3oWRe4wFOimET+yaCNacTRBuVsml8Ur
s7ky9Gr/8Na9BsjZhuV+pUrM+wAzlxxRKOEY1o+ooIc/EPbjplLdbh/FK/TWNl0EvIhdkO8hufTm
mGzxIJ7zIfbQzp7+agP//YPA0jzrk/9Ydyjr4aZGTbUprgJOGeWNc71tQs9DHIiMzdFw+U16oMHM
jVCAZXPkPpiBFHO6meNyWSmUJ2J7dJ6uyLsJmApiy5mm0XpgxmqMrrwDT+sQEeFkNnS893fF4kOy
uBa/A5O7UDP/wzb/QbkC+UC9Ebivh6ZNtQ7CLfmVz5XmqtTjGy/AJ0qq+4cllnV7yX/tWwz0qqhC
/XVHhDfQ05uX17xW0ofynkpIYprgR+9Ig8MJ+qpQ08BQlzJSInQpnPyX/Tdu5eKDgnhM+c1yKey7
SpgdwzTePH1bUH5bMzR/CF7PVR8eWtgbeoPCZ9v755gYRporWDPU4FMNCXg53VUrDB1RVeQYNYn1
z3GLMg0+0AQSHZe2gba/P7yXDGXwK+jIkjvM+TUyXzfyYLxeC1r1mtBsoa8MtWCohZDnxxWi9Arc
clwftGTzW1XvlSC183MqTUpaZFnuTnrUNyQVa/dkKGyModkZh/+6KPJl0R4GKZru99NzjvwU97k4
Gigc9E4jeYQbJ+TEe6CkdB1tuFwC6X0yQYEAm0c0qg1NZtfwgFaM/4+sLMr6FzE++kaYDSfhipS5
Jh7+Os5D8ftx1nX64LNz/PVyXfTG9apuSxVb3KJbt87dcLByRIlyl1t1x/xSVWkp2pCI5gR8LcgZ
9/2ycTZGLe7QA5+g1sLtIGRpfa0H9KgzxUf9wYqu5gS70Yy6p4mkoUqmGCJR9lZ5xe2BICl1/Yo/
J6WJmNJOcvpLij4ZcR0uPLNAz4HBY3Uuj75ZAjxGR976UftwRsdYlMHf68XKXAm502XekMhtokHY
L8QhJlgmTh41hQSFDbj4iQA7qauVtUxKknVv/bhCx8pt+bHFfVYoA9aX2H83MxBm10LdpMs6BNBE
EWBGzLfpMM/iyEIpmINS0XWL2XIiIb2RoNPoQ9tSs3+HlMNz/ywCZwoVpCCjrQzoeSnj0Ixdyz2t
SMyBjrY8/oVSNNUOZ+m+HOaccWkRPHjexOYPitX3lRaFk6IKHrcLRW0WPhVhIeWXIIJn8rvCIqKx
K0WWnzJ71qGEk1x48cyCdwtec7ii/8tvG2RBagZXzx0RnIWZLku/fnmc6YbDPnGbT3su7UcozdyR
lfa7Dzcueg8yvyJYjw5kspUudE492VI3tveqlLj7D5Bst5XjGwpey7lqJec8Pc3aWr/+fcEq1MSL
H5Qx10Kp5qydbkIm1EFx+DwlphNNfnNg9s1Bmhz2AeysXSH/UI1Gfl/I8MWqKlyYfRWjPyUA8gG+
QetEFDJ4QeOY4HJfGEXVoZbwdASEqNQV+pKgPVis0oGGoihfHCCRGvhvwBS1D2RFbi/LCKYIvI3+
Mc5awy+Nul9IEUF0S1+Bxe45sYz0/kHd9geAGY/pHPggU0UiVYOvWABpOCCMMHWAB2dr0CNpMibt
EErDn+s5qvF4m/WT/cFGoABVhVWBsLp96W2vIVVGtWO26Xhk3yC7KQffkRRAJJa9JbfPpiSQ7p5l
QYdQze6t+EYudvnmL61IH7x/s29RjbATlN0Ug0yWSkOkG3vuD6bffrQR1/jHCFe85UxgtkwJvzAY
Z58LzuXvIUI/nq3Ki8GH2pnQcsXkc2NqVxSrAGVGRsB+tLGsRQzKTnMlQhQ/sfQhsRu2KhNIm4Zp
cKH2U9ekeAfiZc4k2zk0izk9cDObmRuWWT86lLF673aqzMJ0lja9TecxTNLOST6fAc+b7HpXPU00
pZGXrd0VXodBjhxYu0WLqe2E366DrqHMjnqYWIZ4cDKx0r3XkB7ybi7x5EU0B1+n9Vw4hs+Cdwri
KQVtNUN5568ZCVzhJqUiWq9LU1JRhKvPplY4YvKBdUqUqYn0YEfT5vFeNaf5//BE2ZVnzvn8UKP9
9EhgBvj4PChobxYuKefmF7ekvuusmIRaZ461RQ7caB00PkNudvXOkVX5TKec0lmcEZM9lkG4Qf3c
IIMn+WF6ffaqeOi9inzfjr4U6BeIAp6qi46Gf7tSyLOEuCptuqZdwkYI16o1Rm0pdExcoruFiIU/
1SRtFIqGzgufpqQHyaosrTYkBh+vfnv2QIiJSC1J2l2ImKmnjgWWylaTwACeCE1+HYmiqpFHIttb
d4yDFo2zv2M92tEq3ZvN+J665ahapBxigEq7/oeZxDf8lh/qQ+xMVWP8zDVsq/ihEVe9nAT1UgEt
14qhkzflE/CMcL8D2C/zPeQ1g2HaLFqnLf6x/KbfcXb7m8OcWh5HqRoBE3BSMIv87sZcc9ABsDNm
96vy5xaiFWR6q3dXjhQucZxjloknN7vTOuJdcBWWysTPSeEfhVOTrfY6W/FnVqzvGpfe1v8wqDzK
+h1CqyZhG0ymJi+UB9E7FGgdKy61NTLEvSAD9b2IQxJPPOFHdgOjv80OtW4jGULv0VxPIe1wC55r
vcghscgSFNW/TS7O4LzvfVbOdDLvdGaIKFTfv8j8pM9hGTs5LgFPKf5Bcm5hvdjFaR3QaoAFO7Qc
6K7t5AN1aM7uvmS4Kf4D0hpK9/jnB5NQ9GS/EAomJpHmCMElCwGBqG8fvxy7uFZIVPpcXXZVtMA7
Hq8HXQP/2XdpT3mhzjHB89dvyOHeNu0JHaIA8tAsL/G9rsjvdL7b6i/85WSpYKhxHUngwQ5L2SXU
ihFOznVD9AxcENnFs6IL7y1b+ftVhbFGgXpKNhXX9HDy6p0XpZ9LMpWWa6JlFkpntnR0pmzMvYwH
KzRBjBSGB5X9NFPDLfscUSDymTXFp96GWT3PXQbi9F1kS9jfExJcc4nb75UqtgJoJlFcW2f4tSAc
yid6pjB7/z2+l/EAVFPRtAjeWtMowuTIXON0L+OOJxnC9ObL5X62ziZKNG+O77nTwanVnwFKOLYh
hVmHet8q1lmZ3+jpjLOCv/xbn7hB7NwRl1lP75E1pvo9tRvEJkcaa2FDnwglj7X8VoZVykRvFwBz
GfGw7xXj0lgpoooZysBx5dIirT98nmz0MxbgTBrJd3ZE25yn5qce9o3FXacFnGhalBCsTU+WCr2q
KEyXS1IOpRixVImshTMM2+3QCImbNNalD95c1eF/9B19Kd7ZBeZE9OGWVhdozIOAqazGug+vasHx
QaY0A6J7Die/3uPntWDHlR8agBTVCSkGbhn9PbvsRcPqKR+40oW/eqQvlcC5wBO23tBm9UimkQz8
9RHLQuvj0P9OFMpBanAv1UU9alSWTl2BUf2iN3GUvVcyN992FnHV1B78R0xzEIx5VeFo/Wx3NN/I
1GtS9xs9z7qdcDV8nuhiWPGdu+kTFGtVNCbZmh//UMJusAF/ZKVg/JvUldHLtjDRFjWLjriGMGS9
dclirbBd4qhncrTkylaNIA+dJ0wFTNZrfIZHQtK/mROMWODvQpwJdFZboAc3qJbRg3nPOcWDYs6h
AYgqF25+gLJY7s6S0qbxqnKUmECfqeKyrsGe7nHkD5C1JtVoGntmB1NBOa76bwU2EBOc3CGWOW7K
QobVkfBuR0CuesNnTQ+R+naAOiydZM1I7kCQJMMTqelKI1i6rWNy7zQcalNxUxrgkfjagm/lns0Q
BqlGV+hqw4Wbdy8Gb9YkNTG8mzcmI4HQh7/X3JenJbYRz+owZCwiwwZb2hp78bjS6UFrZlE36k6C
Q6NLCyzW/3a5x28oBJm+PVuHB6GL7xbnSuOIaP+CpfbTbsneNiaV6nkvgWB2PUfBf8ZsfptuH6bY
Y+o6gCFUb6MuYRsNt3dNMllAxjAVrt2sUtoRKQVAAMtzeaxT3VHiDV1qAchlERvyV3b73mxGO2me
wQQT34L+KWdZ7KddSr8L3SmJ4oAVLWFYwCoxtybZIFWg32lT7gXGIvzAinG3IxP838yFbMhLJCk5
J37943nBxWPYpXCMHE7W8sU8BP4yVox7gsuhbrKD1nyomFj1lyUOrrwpAcCPY01JpUbMK8AGQehB
crr+jAsQ+h8Anvg0fAc1GrMzJU3SOK3qGveKT+M48LJhjA+OE/lhyVI1iKR4LMdQcbHHWE8BhvjS
kaaOVDQehz0Ps90FSjZzANtUGHZK7OTIvuYD44r56fr+DdLav9uHUsXUabglmN6jILJ3ohVNpS4P
GjB11sY5Ou6bFfk9nG8iNcuZ0tI0mhuByJpfVrE1uFUMwipw71IDpo/1JhH6zzo+yHpuKbDFIyHN
3f0RAsIQyi3w0clCsKRLZqE2gNKikVK37MkfE6OAlEAU2xy5i6C592O+QSOf4TPGOCeBsXvRbDir
DxySA37yVDBZYpS7RfY8jAXxqKAaWCiL3qwp8d1yduxsv7iur2vIvykH0kDu04DsyCZ8B8lPKwrf
xwZFSDmvPvIcxYbVkaI7DYVnVcMsOln6dJ2V+hxWpJkoMdmxOMl6tCD5h9Bi2+Aer4SQIofPKcjz
hVm5TXyUTSBc0tOZzfRb1pFZ4CbVQEtBUcHvyACLJz5Fge2c/CSjAsHe8RR/+L71aBQTujYKz7xD
z/mz9lwGtKTmaBg0jtsk7HD8cYEXHBGVlF1ptt7a22uJSHXTPUHBQ1CROIMIR3STjaiko3qvAYx7
Lc/Wqo/6f6bG/Y/3MKxC/FVcarQLbPBIo85i2MLrEDt2ZTLcBUdc2eVbxXV8E0kPoqJea3Ln24rI
6jgLzWM3f/GzwLnYQp3piOvSrgjEmlc5WET621j59B0ru1vZjSDpF1NC4ErdnV+IbQHSolVJu3VM
uHnavOsyLOCB/0Ly+0YB4a8PF7vN9INEvGchRbtcYRFCLsDJdxqcJ7iySwYScqrtZvvaJtkx7b+C
AblZ9wPusTQ3GC6PSi3vwb/+j/WznwGfvrLS7nAWl3QmhHs3bj1+DeYvaw2m0xMC6DGytCJJkdkU
kcRa/jhNgRBMJY39gLQL5swMS5W3uYUFQDJY388MIjku+rvZEFRZIWx4CilqZfddlzduch0ZeYOm
V98JnxE/a1Y/3irVqBX0dH1Py8n9jtC3Ri9D+OQle3kXBzqz1bnxoTO6JBXTZJfnXdo8pnOucVI4
S+zUMuG+mIqkqxW2x1crRz1WQf3aARhfwRIsaUUrOJACbIY9LlhvLWUqt4V3jifPOy9cGjQ5a6nb
6aXxvohZ4H+ZH+uLB3q3RHDelvb6pquHUzOXOPYAheheK3O5TGLuiV2aceOW4Ww2xHln03eP5ccq
hqrrATDPsMIMiTA5IslU6VqYp2aZ3hiuKZYB6B5eDYhZIG9mGE/scuMZXkPEayBVjZTkkmer8L8/
2F0P7mQCQCdJ5C3Al2CEJpYxm2IsmXj5vIeySghpvX6++Gk+LAAE0kcF7sLCxn9fsVdQiXTQjafV
9W7rHqEB0LV+H3DtcPXpyZLS2UN7AsET6fr4gcVN/D+wspUOMLm1pM5aNmsRfjhSe62DHbeiHPPl
r8iK6wxSC/LR5WfFFuaKDOqxn9gryfd5SlsVkxRjJqXr7qtmOO+3PX09oSzd0GL+Cs1ltBcohBuS
7biwJujVqGH1amMIxDHdA3W8OhjDgjDsTuzLgbWDaBBQvP3JiDP+ATSg8nNU/jrsK+A59ZgEHBr6
f1MefW2ZYSLmGGxx+iuSeqN+agphodeW+O8EA/iWTMvjlyhw8B5f7fnsBw2hUUl/yWKdRSnJDH4W
y9ZPfhbJVrleoYtQ9XoGuTfaC1Wzf18hhX3ok0L5DDFFGInMYtr+avPdfWXli58bDDSH4zy6KY/X
huA2F/av+6MPfSkA1QsdgMkEvNERoC9XPwVPpzjQi3zr3jn/LksRb+D9VccTtaac8pFNyxeabJcT
mgXioPrMBoWr5/kwQIo18F4VlZC13hlX1ihr7WRww05jZsGcDRBxKKqo05FIr++YXqJTMWFuLVfZ
+VMEsFtXqdT1ShM33SHL8fxy1ELcDCrxWJbg2dHcA8xZk8dV3i5FUv3cj/ZErK8zpm9LPzNEVhpg
5b18h3zdIF9d3KGnzXL/Jz0NsnP7Jk6C/wTAkRZcdXfWqGBe2mAAdFpQ/NDtzTFpJizrrYiLb54P
+uGFcm8JlCjdXcD9dNmK+HzK3SSj/1ckSajUlv9lv4AB/FOabyQisaj2jZqNZ+6SjVoOrTZZkFMT
Bt1SYMVhXVwKjTtlXB90PnVwDl1CRRtiztOoNB1X22LsTmau3SZL7CEjVBzw76z03iFjBZGQZ08d
M8PD9Z5WJ+O6KBQlWUXdYwEcs3nt16Fvk0l4/A1bYOQ473UwGWEplzWGWPsXqQkGcrL8DLDaDCRu
cEWFa7sm/pFepaMkrxMidrR4jHHAYoO841coZZTIRW/wKlCRrELI2kSP9Oqhu/KHI1r8RKwOy9tB
f0Rn7JQWn7/C/YFpM4UaXbX1++3orIyBdxBb9yZHhIB1ZaCKk+VDEosORyQ0cRSrN8js5uOgQTOS
WA1087m2FLQtPmY6l0Wii14+Geok3LFL3+nxZBKZKg10TNlalwcLxmKBmVlSgfW4Rs7Cs2Vk/OPa
kzTnQJcIEzbSs1ZzAf2321d151IMeHftyc86rQnho7iH4KNG7EEIi+Onzqw+MQdeWyPgxGd4d93T
tEMFrpK8I26r2kTSuzoIPZfPBDu4rzcot0mXp3CC8Rrs7aI8OQiDeGFT/FbAxocMFsRfHwYQbuxl
3yjcUdvHeL1JF3GPCc2/EzkunA5slK2SZgwA9FOQNGqGcO2IAqvSZK+B/JJgSM3oTM9YrwAge0oo
3f3iPRMmtP1GCrSM2dCWym+FCmj/DJktuTJoROac1HHxqwG19Czhl09wozw5X3tSkgEFbA4DDeEW
tNh7Ek/LDI9N55AnKTqVYzpKGXh+IFHr4LD4K9SoON5PjmC6Lt3Sj5cWNOyQK/vRjj41qj/3ZWv8
g5WyoOQRF17A+OUMiuqTVTIBsyQJiIn9TLqdQL+seKfuxrYH51LWnaSMkjuGlNmRQF8lgN4F/tY3
As45n/OT4dkGSdzcDLkuPdAhsiq3F7BQrdBlTCAinhvQd5z4iUUggOAeS/s9/m2GvrIa2QVDL+tQ
KilpXmCn5btmbY3gG838RsoFUqWSG79b+3eWnpi13CBWChX48AVVF34+7BKS4OX1BY/Ug7MhKDAW
b27wQLZtTSklz95nf72EcEQgElp0LgvQmcwr+Ry9AT5Iu5gYa2CyNUx4roUYDW9xv2MZbzhFOaxu
Mqpmb8hcBVHcRsoKiWQN4mgQGa4x2heCvEGptUpCDkye9G8SDIf0oOIJUnom+ugsCu+U8+VLHA+B
WKvk4laF6UmH0STyf6j2X2PoHQ27Z6HfM1OweAnP8NtJ7YaWgWcc4DxCyttH4bmZMI+DDIYuiSUN
HXnX0z34wyHCCZxTowKKcdGE/rBrdmMtAmfkHs5siB35j0HoozSsAa3XQE6fg2u9BGID2W5BtbqD
XWxxlDfNwmfW4FJDVnXw7LSdohKpYyre7GDjLT8MyQu7aqg9Ga0NyolEoXXs2m4yLAE7RcN1imVY
ihdW1FlPIqZDBjOVExXqJPKx9vkGSSc/DstIQ3M/EAZwBHv9tFl9XozqTRRby2RKQULf9lXfLDLl
LMjLuEtZ1UrKHiwZ7pc+tUj6WJwR0P8V6uVstNu6q7wopkVZVkQHucb0c2Sebc6tlkVXIpYXESO4
gNrUGpk2MGsVZb9dj8d6O0RWqBYwUpuyVvTNRwgq/2fQY8uZzGT0oJloQfFY0dHQtiqkQ9biuRQr
MCUUKEafUYVJiA14Tq4Yek+6FmhnCIweVlDi20vJrau86xLbTWepAoLDYJUg9g6Yu0MLuA2YNwfI
ROVREraHG3a6W7PRcH27C+FemiBJWqu/g3ebBwjmFU6TInx8u+K+q/xdyT+8TS7HSQHaPzrIt+FF
Gv2ePOeeMHMjcckk10B/T8AJNTwF/bdny9quOxzz/UYgp0Eso4qYHFLmf999IjRxFEHskzE4V56T
IQcp9WDwpklqB4RukPvqLNxrOFB5B4nnu2elktg4II780ghwieicPuz2NAUXFARdThEbUMxJfmu0
RMtXrqS/DP3WkybRQCsjQbHt4VTjDC0SAmZzQCAD+sqksX3NiOM//r7PnZwLiEmcyucLhzPn47La
KaDGGvdNrdDzNJBcPMDWUCRwR23WU7tyv5kg8qLvcHOySxkTvOl1skgTPc0zVmhgzkuhM5yMXO77
Qv0BuoHwX/X036qVKiosa63aau6c/JT6zX3OCMu0ER0s5YWgmoWW3Svj+uzWHN/urPO15UV/4CI1
drSxiTShQfu5BbWrmQC1DjXQHzljg0osa1cAsG3NThpc8dMpF22RgGHRCTesCc6FW23eEmkf1X9h
Ym7jinleRFGGycNWE6pO3OccwusSb5KAZtfHVds77i2585sJfFdoUOT6tuSgKf6Rmtmyhp9mS+vd
i0F3INQkZybPe8X6ind2qEbpObd5/Rh34pXLCjJqmscHU2Z1Vg6ck1v0c6A7301pqscjm6CPgM0q
SYukrMaD1ZqX+9BaYxR59Ktn8n98iCvX9KQb24pF4SuMNSc+WbfEWW75MVeviwF3NuI+GpzMy+Os
WkryloujIahJvYJN9caB7r1IQNBwc/UEykvG8cySB1fvTFqyPzIhf++Iz4Usu76ZFLLEb85Iu1sg
uMZhTLJBKOYnVkE8BqHTH+hPn+Ss/T2LQyjVY+mpLS7Ah7TTdR48kgf2AQVH1Jg6+0RSmCEhehnG
kJoiHZPXGQ+Y1aItmyq+FrvMlJu/CPZxWBaPMvZjTAOdn+BqC1xY0vw3mT5QpRtQKCeEd9xT//N+
lrzfSxF3KVVjbeTWC/wajKEY7rhIuj0ZJJ6r0IAKBOKXwmuRjl7TSt9FyB3XrALo6qDifjHUdDPe
z6KR7fVPjRWuX10KoDpMICoZAw2ybytXpcVcZpzQNCrOi92BC4FYFCBBg0hGBa9yLaaCmr4KDtMl
QTfa+/gyVzj1q+ZN6Is1hV1y7V8FdrD0r7R4Jt6hrt+FolmlfH9oIBFX+COm/ZmXs3Iw+irA58VH
VMt/rFc05NN+Lgx5llZxOICT+Azwdwr8JRIri8VGmns6E4XeEp8nFx4mbppfwWfwY7YOaQqIOsZb
oB2tAHQHfWl2Q/yGlUhCG9M5k70FxWDPsoY6YCgC7TnZ+KUVpaXO6LmEYD3FdRFZQPZCbIft9u1M
QWBcLIAFule79Jgf3Dyc40d7iuhx4E6e0z2aazTDwuU+OH30dP9mgOPQjBVgeKk9wefZg6D3dtc0
RxQ6AJy1uT9bIrTmEbV7ylJQ5msOwsdyP5T6/CSLBhU5lUHCabTG/BMdJRBQutatkJ87STZYyt1f
4E7kpO6ZfBeDUCi/rvH1Xu7qAHgxLkdsZFB0MIGDy3hoCzHObV2iABk/shE6xDejtN9EgPdrFOFy
7CLSt0s1a9I1mcNr6gDPboSJdxyT5fIDExINqA1gw2DCzKJrFtShyhFxpuTXshzfyyXOB0lD0h/f
WClkSa9AdhYmFQ+06NJ5ab+kei2aYNHpCSuyQ9IVq4Yo5koMuBVDl1ZhT3r0ZSYrsmqIOOP3JH4q
gASPaLtu19a4j9uwJ3/HyM+RF3L6JgZFZ0ozaNBb6CJc3/BNqjWOCFVtEZsh9Aoi7lmSzauNVFRz
HwIDHfOUWvMtbNhU8KMN11OZYNSkzYVJwk7cFLDpQFig7MrnkyGBlrjaTvRYQK5zP3SlV1N1Z7pU
FCkm4DcXSvgMGLcNPnENyc1NPFJhJW5nAMKctwaPxLzIwKwLutJuR2CY6xXTTRrY6DPtdxJaxqJm
FxlraB6T3R5pCsH9oXmpKVTbQ6wq6D/MMVYo5029B/SwWZy39xSrFhSRCqaUeUUyRiMKzqV/8+Dv
W5FOocGdZOF4HlnX87wyLOqfKq64wJLGL8Cl9sTPrsL2yvOwHbXXC0+qIwcMRTHvIAiGhB98sYpx
YOds0/EX1ImsLJxqfeuR0TP38aexSoRV5zimECYFkk5LPq6zN+GlzT+BYLEqy/aRFWQXLrIMfHkj
lcEy+nF5oRLfOmGaWTal7v+xC4ZCOyD7e6LuJkmksUjVtwI+0z5WGn/mjpfX2SPq44HmlTZ6MxS9
cNqkhPgploKTICOLKqloucP1caYf3MlDBWRxJwlB04LHrky5J3PgRBlq16g5viOQyxNVhRGr09tJ
4OjiN9CCH4zrWC+1mItiTJQWyLrUR3QzZ0Z/1HHNmq68EwxBh6Ax2V2u2MsLe/xiGgh1EydbWVZk
+X44ra6HofWaLmHGMiPsj1fUmbR5YmpB+IzyKA7Z3RRByKsuY/JKSMxGB7bXfQ7ZI8k25DFqOzMK
ePauczygELbLgT+kIh5EzGEpQpce4eFheH29e7SMF2AeNo/ZeNDgUiqxeqA/FM18AtyWJm0xZzAq
2ArECd2zncICgynycZNgEny4PYV5H/c48hPpQdzFSg5gnIy2DlT27Zb6EYPFkpl1h0/0J2SvgO5a
TxjJvSXhVFH6BtdigtdrKqac1fu6poCG2ElZAzceXxzoOOHPE5+TpucUdn2f2RyXhFuWKZiv2sEX
XtNW6NI1EPfxdrG9p4qpUMW5GGSeIeyb05nnikGn/q6MJbwMeU3BXSjNtbQvHKaiTKe8Ol+oUpfW
bgqslDJeKgahgUb4V2jTYREgH1F+zE2OvpgU8cUZSJStnDWAqVI+ABsUxbZg6rhv0ipzJn6m/C5v
qZMEntAkriW6Yce9yTsFjzTuYtwfkmzvGCRABfQIYYLFtS3DXW33ALvbOrM/iGopNlqMYrYPA8oQ
tY3rLuA/d/drGbKyzve0qf+4L6TYAXXGXDkxEKNeTxlCHwS52HKAyAH0zNNXHuCIg3Pu1/HVwVaJ
NLpvJpQUxGhjYmBKze4dglojo83IfmRBtr9OizXPUom++2u2B7qSDCk2z2+EvToOnZcr7jnxtU9H
XRXw91c/+ZPKUmX20lIHGHZo15lCM5aIOOMCa/sRBNeInsBwi0+nzRT2/Vmnh0Yl04PBr6ZCQ1O2
5efahJi+h1BSwSpu8dNYGdCzvvXoVfeqk37jP2nqeXc2F5W/ek23SdWPnQTFqgAtKO94uIzXmtMi
BTOHhZSo1AoDtWBNZZCwZ9+H5FGb/u2aD+bLlMdxPPxOE4GzvW7sLc7HvlfOG4b2OYz8u+T9kM26
HbDre8aC3n0UL66vBxN9Z5yY3xB5fx1Pe97Se430dzPjLkxx81IOEwf+u/kUWcM7/MiBJBeqGUIY
CCIm0g+W8NhjpkGhoLEHv8DDQJrVsv6txHbbSTSXKpAAYcFxJ9W133Ll1Wmb6vBl1MFw+xJVtFdF
sOICSG6VoAeOPCrQEbSl7Qa2Yg8YdJP1h6KSllo7Xfp9F+NMyVozPo5/kidh5/W8nv3FrZ9Vfw6j
tF1CJnGE+p7cn4id6UFHFhnB1ULOXfe6ol2rkM9/1Whxs71yLXaBT3aizJkLhtm1DcUz2G9OHB95
CJ7jwscY2wVazST4dn9paBTWUCkz6S066fbRG1JnZvjnYWJ/tj44eUyZ7tCJPqMC5FjIBDmTBvXJ
9mIN+DKTyQ467cP+U28DdvxhzUveo4U+9BNrw/E8ft7fiy2dz2sd5AIoK4KKjVgFxE1VjtzYrZ2U
3uMup6t9omoD4V2O9prsGDSvhJPhv9HsIwjGK7i369wVNFWB0qISGDv5WeJuvaLK6GHNezuGGtoM
lXeSje2hYpMahe+rXfbLIWEZgq7Nr7apGZDY/+jtQz9qeCGTXD2q3rARNqfLGjNHxdPyIGCUj49m
JdMUpoISGuHnzeLSAYeZwCgmKJNtYSr75IaKXbhFlSWaN34mLcNdhIoVFTUsprvA3bdBiY2dx7U5
GPEaUpNihKTTP44r+OAjuS2rJXw7EJObi2qRRl3BHOgEXHeeYMnRpwVLcibYoNpBqfhNH2Hi/eIt
0r7zP4vjKzqMqlKU1o+GiEvQZOTx/heeEw5BNLA2l+8BmOGcmvyIRW//iaYCZCKi4tFtOJC7C+sG
d0DP8eTSKZiglq/Z9T7twOLXHkxETfaBS63OJHqPp4///Jq2PfNY0KbdJkg+UuiZELIETc7h6mtM
0FnCLkl9XPuhHSqZBbSffxfQYVAy61PB8E/rdMc1GhyHV5PYqD5BmuqtkNK7Jg5Yp0vaA55v6n7v
SssMwkgMdKpP1EpnylsbRyF7Fgv3tO3A43TohKPoVmvLn+5mC2F+arbaLmuIYGV2mx1PB4/w7RNt
IblGMLiU/61Q8FmKP3DVF6KUr3vTCKT63mmO4iZzLT/doxw6cqY3tqQKWHES5USDbvOv6r39cS67
GVgkCR8v0PTR3k4B4T9REaE0iYxcFUOVXaML449x7mMPXbjPyXniqDNZSuOKlWliuPhsKBh5Qf+S
GTLDKm8dMqr3nU+Bm9CJH55OhGxLR2yuI3JwChve3v8/3ycDXf+ubBLPleY58dqpXBg4DfGAAtVq
8+0s3iXE0zCbQJk97h5FX+46XXYJit4eSVamibHdJv5NiyPDWgaH9luIqaebcItrtw1AYQgDtvcJ
kO1olxpUxyCISbjk7x/axiiw9HhWoBpNUo6yBqG+WpJL/1UffRLauqI0qesWk+8Hc40uDx5pPv+w
R6y2BUKUHASiet/+MFPO5QI98o/icK+WAXf2RHmA+NMoCnxEjXSTSNcXYxCuWUhpPrZlX2PelQ2c
2HoFitnB9aCFQmeiaL2TciIMX/0RrCiu3QvCj0MMszqi17xj75imJH7BNp8s0sFElxK+WLCgvzV5
rba+ozv42AXYaSzWk7pXw5ILqjkBiRtCT/JJB9Sk6DI7eK1zizPSEYO4B34NROZcmiOAv299LUak
jlwnWiLB1s2oIHX05GBEY9V28mpYUUAbEAXW+vDoi6dtOb5nB3kGPopTYC9xEKIdPmU26A2gAyYU
8bROWtR49hFc1z47hgWDA9VO0iAlqHe7TnGneZE4y7qQ0kSZiqNbmAk93m/Iumjih/6AQrKqvEyh
m6QsLSNLXmZixl6a1fRHN8jYMbCUCICdgqxMCXwZfFIVohISD/Z7VV1A8srSFjMDi0oaisAzNrMZ
J3QvoRuotangleUhmx8lhSvrZMciW0ZhwzGSaDPYLNqUzz/vl3qOA9hfpq2igxG+vsakzWVaEMZy
3Mat4LAXBhW0IsAp5WOXeN/8GPY1f3K8Qk2sF1ZmYvi2Ad1mcaZv5fSl2Ytfe8oCMFMzJxs9V80z
emmQbXQ4RzQJGu72pHc6DkIOWRCvhgnOczbzqxwPw/0L8SEo9JAgm8mUNBov3AYKZC6liOBdzFI0
hVvw7DRX23vTdP/lCg9X+H/LMPJz1OqYshJYGqfiDTk4ViLgftIU2naEczwu+ahPsAZrwpsQwTTa
kf3/F/osUa5em/t9V1FqfJGi4Dtxsfi0BwQiMYoIoHQfZlsiDzHMSisMHW6jo5N7UXDkhhjAV+a5
sSVMJR/4gyuSJslqDIqn2mgL1U8KMOPkSpbBeChOqJwY+PoybFLqRT+Tr842/U7CJs5czFyGSufQ
R3PXGIBQSxUL/sSKVgzxmIjIuDDqycE2rcepS784fffoe2wou337iTSaCqWfmlh5ByT+it7uaj0d
a8iysCiLVAlgr0E5xKeQKhqi+MfgDx3NELGY+43HJjaSTM7Z7clfD9YFY1EjHjb/9JjHd7UQWQt0
cINy+hCbf/s5qEBTl50MTA4oQ8ssmFxTQk8WPORg5wRpsRN7hslP7OaOcrQMWWDvLMiA4QfssYui
U80RD4Tj66uoKYEnuxZPd9utTM5rClA5Tb9KIlCK48ccoKCBBqfjg3p73CMdvfuFsokgFNFyESG4
yDUqSWCbpuxgVKF8YPDIc/HmOMdTuAZxBB77YjCAey6fPnJzcNTBby3JXKvfv671mTaJ1Xyogg2m
uOKCnE1hqe8OC1KCg2yuScPYD6OAweVMHhPTS+Z/muwYYSxV6cJbM0dli/qAmGYUoQtsF8xPwa1x
3ChXEPTmqQauyiSiDGfK8p7sC42Nyq7+4DtASdmKkQRyATfWPJqlt7PnzB0aawA6Y4oYq9zTIQA0
L8KxiX7d0hKgCPEyEv+rr0bv9qcwzs5faS+RwL1H4vQJcIVin8HaLQrtBQKwYiYkSJDpmm6zMxKC
tuIERbv68g6HWpN2Sv7iOpTWfKhUKeQdYy9A/O7gOqPUQk7hpuxWAymPL3CGhwelHaqSZRu4exVe
K/xgd4R54Vtp/t1uYEj2jXO6lWl/2/10KaoKqIDseT4cNwuOFoJ8VsZPUA5BBvDNZIoTAGn5gIXM
H+2EqXZY+Rf6i0CpZKi0ymWjAxFJBVzq47VoDFH/OObULo73ld708euMFNW2X/AKSL7Ht1T+FqoI
Lif21mjpKuzIGOzBaKrCqYJrZ+37G4xIQM8IWU+8MDxQMLqVqrMfxr/Q5KqJuBP9CxG70X5ni9If
irknel8ilk+3doJEq7PvrjqmoE91Td0dtVw6oTeaWig4t1RfPo7G1GiesriYw/ANXfBiKn79Vn6w
PMFyc6RE+f6Cd3MjZBQp7Z7jw1wog0fx7/QDgWIhZTOi8M8KtIEwl//P/EoGAeKV8xLcN+FQZbs/
BzyMY9WjvR7do7IW1mbHGtRkYIp8nCs+x3hqo3yzh9TORd3MWTbWzZ9zne30NTxBLKfuYPJ8d5/9
umGGH0xF1beUg7ij0nH3p4Cr346SqskhvWx2ij3M4hgsKcI4LlF6nRckkREuKG8kpaCljK+XMMcn
VZVlZS3x5BTdY3yl/ksjOFL+L1jl95dn70VIByKRx+dmkSaoqf5moEmBH64OuO+2FXskzLrISwrt
DK1xpIpzoGUios3yKjjWKpZnZah1te99T1rpuBF4pf1Mdh9gslu5MFC59WyEWy4/5o7as3IYFpcQ
0Dg2BA1eI41IKixQ8C2JFAsrKR73iatflMfUmdn8WHX0dBp+iKZneLdry5mUO9wk0Iv23Usww+/+
jybNhFWpaG3c5pTXNoyBk3/zMnrj+HvChA/y+ZEUazFgqyQjYXq7D+SZdpRQlZii88UZr/08BXFI
fCbC1UIrdxiICrEulu/0QAabdBC72RBpKqso9jJEavWhPURGYszhz2EU+OESP4/Rtmow4mSXjnMa
1xPf8/2oa5E9sGVQoggfHD9sPBJOFp54XB+pzc6DgFesqhxQqWFhko3U7O0hjDIH2w3Es/Q/tg3/
LVDBF6C69nth/LxqKiaxLVAPkJeEdcJqkXbeaqmRu7I2oEpxK9a3boAB2ngB3MZCL84Lzf3+jdWB
5fjjOztJ6O7JWq2VC1zG5xLA0lJKKcyePFll6PKHWNSZYkEZvyokr1L3t0jLEOJiA+mmRG73yww/
yGthy8LnwiLJv4hopV69umeOrhT8c1EauxtyKurmKStAjfiQmtpWAntg38G87dSQmtmz5VYRaeJv
wmhz5sqo2oVVjS9WxgnWjPnSiyjBMz96RMQdIcJj499G6E1+0n7NgAVCW4mDLETuktjRWZEjOUXB
1LJtq0Gh07VAuV/OOeod8B10q0mnk/mdQjLxFk9FC6hQ2/idwsFwmGEsf/LwM1BSIP2dvaXKxw1q
TOqQl1mwPvG0rkYrHbuqqd1gx9J2NjVFxbeqQwsVJ09VjJzGJiOm2qdFZm8biJjbDql5scMaO0k/
D2HP6TMSxpupcr10UYmfvYrTQb7n67znxjNtYgmodLuLq7Z88MCcFJgcMWXE8pv9ncVvQWtRL8np
Wo7YJBpUXpI5sqyyMavSw1oFjth2TrqASRAsOduStHFkk7RxhHUiHqTBvb325NGJrljitSCea2ub
vctM3kdkair/CgvmCrZI59YnbyBwCS6ma5BInkJWY/QJaHnyw/5zq2pEKJ0NY3rJjBOA0Ancm87m
/ec7Q/5huQrdVNBbJAbD089es9asVYK5C/pO6TXEFiWxtDAA3CTHfYzltGmaB3YO9DsoyoTY50ct
SxgccSuLYRD6FsQHPnyUO0xsswLM2DfesWlh9neC5jvLJDK+JLXfcLX4LSynq7yGa+38SNRFtqXX
rhA1BMR/6dMn9hMfX6w5513RNoReeBLCHkRFug7ztLDRnM2uy7AOtQpdQYYEiH1BUR7GDROGPAHR
XeWL7+WIuXlyLVO6Q2caPRNh189GyDdkSoOu+CqT/2bylsvbP0tb/rDwcd6/usA1vWxCLyaK6Ok7
YBJEuL/uCA5ctrBG9vvF5IVrEl5EjFbo4uGqeauLpUCEyMisQMqFH9MZ78xUtWFNi/lWEEYGYASo
LGC23nc4ee6NmRIMo2u/TfR5kanwXtGWD+pBqbcLvw/fpNV2aRWT8E06oQSOu41hKfTaoRut4SzJ
LJfpvSInP+c2pU3tm36I/8LC7ktHJw6nmZMVDtobTVMJM9vK2IyXhewnm8dZ3jSYlqKLeeBTr6W3
Wt0vue2i8kEN74K+LPbWnjoz4vEbW/yG4Jsa6MqJ30FWVQyPc0tx0H41NxK75tfUKmT7LtlDeNWg
FH+s4XXCBSsDh3Evq4FGTM4P9cF+aSddwvYWroWYqRsqBF0RWPLF/Q9X618RQc0mwmNGusDeMQIO
tm525WrLpyZSEfVlvlXXnPXIjSesjguS1HbaBCd7/Rz9FNHOZolhYuG+aGw0Oib0Y5m2s5lhXOup
kqIEQ3KB20fMl8CJ6uRRZavbAHi8eh/2FvKdFGXKwvAosbgtudgNFj1jA3r6lgmN8KbKyGAMyvZV
Z0WtJ1q/t1Ygzc4I+qOLCo72/+B3Vc8xYQDKywHOggqX1GTpk6e34wDH2WbQ18oC6KIkg6g3YJic
SJwM1Acw3lYF5rE6pC45A3llWP6LaPfvQUSqP/fiZ8igJ0BAb3j/7BsJASGGTY021ZuHNwUgfr6w
GZFdN7XcLEydfDYLc1J5+Mj8rMKvJwfgoPKdAs2QYjIm9wFnrf2ucGZJzo3aH8kmFRpTInaZbrF1
yVgTLpQS0E5qu122gQpwGDaIZcVBGngxS8NwRoVre5eSDaiIY/WcZoAYDE3nFp8giwdatzVD6Fhy
Hl53l/pOVbrG90Uo0SkdfiDokSbgWn2kmYbTEXvCm8r9AssdCZxy1QQQGMn20F0EB0fuMWu+Sprx
X65PDwBPw5nJQI/kSRzCSZ13H6bAz7nNERa/QtNgvUFD/CTcgR7k9cKfR1HDqvdx2TuHmeNT/c7t
ABvxyh1I1SlBHtmIVB/odp9FR70CNlWUX6FhrIiafyM0Qzd7Jmjonf5sVQ49ZrQ7wpp9jLI9266z
373LdlSLaWVy0y+jpM/XhOpPu64k8P01L4DOZ/C4X1bIv+BJhiRw1A/JROozJn7VToKLbruXyJZh
5xzWFPBHfErbVZ+MeKMKSmIUxHbyiGPUqWZfV0F3RE3BBEKYir2HOA4zxQrFT4V3bTfTNCMCkOEX
CSOg8mOvCtUXOzfkK4I59F+xRWBHpQGM0/6XLw5/Do/ca8DJ/l7ro7nWFP0INFvHLanRRxiwGJ/Q
BqDjhl0gbtmE7znarBzeYOcs7vNbSCODPqkWHAPNHwa8SWlMuVp335FJmIj+fG6CeKhgjRXhgVEu
aiHYgVz7W9DI+4layvcDyq3E0xi9BXsBmQuGiEqZoAhRSjvwL5+0zOiAEXi4OBOwgTpjZOdXT3Q+
wFwoEiLU2TNRY6Ze1w9DegCgMd42MBySIfHIt3amAMC5MPSecw4np0tO2GAiuCOGrQl6IXe1ji56
/3k4ijtTWE9brPj8a9gbgDELqcl4LBgDeUYkKjIFjPBJ0ZDG9ML4cFN/VE4hmyTapOD2J3mmAyhM
wOh9ZzNYgIsvb0xL60XKUhwh5hfLX0OuGCwDWvKthWi9Ym82r2r7jB3Qr9p4vqir6progMwmNztP
yVYLtWcLKK7cxHjpCsEYqKDayfIqWqQNom3Mhs+JfdSkBNBG6LszYLVWHtZ5ZYaKiWG5ROZfWIu0
HebiJBmWUD2qsTxvC6Bj2n7jY2UmvXGyiJdJNlObKF2+se3SGojQfE2KWFAiWUO2I75yIXI7mcDD
oWZ9ZIGabnyObuG5kBJd5p+FT95l/fmAnirNga/CowXkE2B/Wbq/WEbgH+fu7aLPV4pow2Nfob8q
99Ns8xrxUz37ErIJ4t0iOR9+pP0oWL3kjTmyxcnQTFZgDQJv4m9LQTzE0E7OR3UjN6cWQnh38yWs
/amFq0wZtifn9mMHIRheGb37s5QT8/cKPJFMd3ekPmlX+658j0DYyvYUnme1MiUR68zPFnRYpE85
5RPh+BzYAsLzcxWrNENL9VjTwAqb/7WuYFkxe2OuoGvrm0izZ3TB2vHDVwNRQ+gkfapZKjLX+PY3
GScjVB2DvsHsTYAbuXh9gxd5LJTJoQJll1PFuUfPHFcymQ3C92OjlpWGZMA62ktiXGytsenfa5PM
3rAZlRu/5jf15UP518EmpxLwnVrDi1xitRbJhlm9FligNy/d8llVUMzHwzVxgsIC8JXskN7LzbyO
Xcdlc6HmVRlmbbfJelr2itXm21yqmPh8G5dgfTncuSeUnbtBsJklN+Ml4UHHNWLQoPn1ie0UWrXS
jqAYdLgl5U3PqTa3seM/2XETyTPX26h4k5i/3XzEVdoUzF0Me6e3HIVk/ZOpoCrIQaPaieP4cIKF
pdFYRbGkSLi1/TmpMifPXVeSKa2QcV/LBDUIlMK0NMgRuU79BHq3ZJ7dUb2DA9A4E7J/oEbrjdfy
Zutnrx4hAJwDrYJV4Zi0uI5DGpCgW+f9HuhCn6MtK6veVEKb4uieActDMX29SPFvuM+T9Or41Z1g
46S22oGIL8q7xPpoSFwtuy1M4R6ezNiP5ZPHrlOM90MDRvXgsEacARHglkOhYycE7aJQPVvb7zTD
AxoHTLe9So753MFd8/FX5P28x8BCvNOlIS3nA/Zx5qlvquwXDxgaqg9bSf1ulq+pBWAYn4vHnr+7
kUJrPY4fUjQ4v6bx5Ke+My9tBJMUBptfmrP8trOw/kAyqSdcknYj1sfvQr0SFw3FiQshJZqF0wm9
8HhUa589rVki6NHBRJtdOS1Dq1st5O7mTDiWLiwXM8z7CuNzxcXqzoDb8dsfUbKhj7bv/QV5QYzw
U2Ys+D291SmMxPRZwUqUVANYeNRmgM25UHH6Kdce8sd5Bx9YxTMTChqOP/QPxWSukRtXQGf5NW7k
/p7cLRgsjgwYAFcc/kqx3K8PIEQ5T9sYYA0siwebXqnsrM6Bf3ci+xYZFZgFF/abYyTtXz0Daec+
qhd+H1dOxhtWe2Z1Soumms5lsPzhEQAjoXeqOm9CJzB5TcS+rH0YRcREE5Hm2FvLwQ7mw3fMUC6d
c8praMgX+iZzKGyCCy34lUEJA9gE+vy6FFADUZH6qV75N2opWkvmvlcMPUQJIVvMOWQYjNQfUhEE
SKQ1pBxVeDrx5/+tQAurJ5Tv/eh7aJGwt0AyN0Q+J9ZsPAXJkbcQwSeRfLPH4Jim55BrF9vVisUU
sQ+5i+mSaE4r//LBqrcNYmLqcE1TiQKlTzhZbDVO7TBATnHr7j7N/gT/gabyBmKoNlaEF9E8BpBW
Ne3xvRIQ0q+j+3PCUJeQmVwYoFhjZvkoGcfrurMegM1OiEmf2UWjddm6/A5k999KnEJ4K84WoWqw
/wVlYJKK3ktJrLyj+sOQ2W/24e5UjTQFLqvSUpX92wngNXxjxtJedi896/KABpDN9SXbAxm6DCwg
kN6/E6eApOKoQoBZ8Go1wXxk5wZiz10qzVmcjWSf1dd8uqnkR5GZ0FFQzvrry00gAZvuI0khZv/9
eC/zO03d+nJx60h0soDZd9CqKRAING7YYXnWUFmHyfzrvEVGGGYCMWHr4OBdttWcrid6dk7z9EOJ
SG4PO1HVr/Uhbs3W9VkfpY04ia/4hQtnp+qOCcyOK3RF6bSMYKuTckK8CoisOd19xYibbTspQURv
KyVHiKZ4p2VKUznS2MqEXm5BCxijL5ROUo2D7E8KwzBZY7J4yNyzCC3Z82+xDOz/IC5BrusaDMsN
tiIHGb7ez1h5EtK01IBPK2XWXI/uFeyZS8sH4wXEh+N5Q8h207O2ptucabfJip+RYvuxF/2vvBmF
wnOAXFe/Rrl2alpduGbp4athjk+5lBG21hwiDenjdMaDgDbHsj2Qr7VeIMD35e7ihKdzNyrBWowL
B8dXhcYvayYBunhbN0wKDSqYIx8Z4bzirgFCaWvsVHR0lxW9BoVi6FbgsN9MjpedE7We5QJ0f4Ld
YEHw0JPDTjNrflS73NVXhh3fh1fLyWTx3ebE42t0TK1uASq7E4ZNoJXuXMx5/MrbEA/dviWwJH7Q
cLCsUEht/1Q0P2LPnnjpxCyB3tlgNUbfhjjW2DbCAtyO3tHmaC5QHh1JYPRkhJ8tMjDb1/Tl5IR6
jDXqQ8QoldtB///uZ/i2PWTZ3N7oBrB2h9au3STfbGXwpVobTHImDT9+tqybC8/idkb1+3rzwf2V
QhNSBBf3JDrX0BlklcXzb8RCumsQ3y+rJBz4g6jDEBn/xwUHN6LnOF/74T/4ri2HhzJDPFJ7gsKk
nGbRKERQIciWwihbSkeZtKRIXKKLrtRfLQrSYCp0EYQu52LjLq+tSYqKoPHx+FhaVWIki/oqso94
BsmC8K56pdbUwYhdd/oG7St/Doh1MEIL1Dgup+9Hq/MthKcxkaxwNnJTZGTxr+4bPIiT7fwkTzjg
k8nq3pHrDlqX3wlI1SjapAxNaWqyVe+38G49XXVZIjrOPYUYtXnmQkzGHptrnm1BCUkpzquLKjQ5
aeX3mTNqt5U0Ldo5VdyhTk+oefUvkatHynBah8VBcCbLDkKs8XVOj4PKM+peKONpvGuEX6WDFLM2
fb9FDqxTbOgWkoxb7tTlT1lPU7M7xr/o7grygrUp+djPwkHtWKWzoO233xshL1RzfZMMjZJ+OpJg
veDXpQSOiGlvvZLthLUPI2KZ0rw8u8XSbAWIqYdoB5NI0axh4yJ0wwVw3J94FtUCR+pMszOsOt6Z
596zKI3xkcQPhECnFj+6v/lUt18I+iJHlKIy/t7StBxsXRW0hTGv9JrRY0SD2LJzEPNEf9mPR/3T
sABI+/sg7XnIaAUhSkv4AsQYi6kHrzy70YudeXiFrVSNP1oUh0MBwKL6AaxzY9YXDSmWs0Bsno/B
H449bn5p+xLHDRq02zgXz/himfReropoKCTHlKEHi5s5MwNzeOLh5//Z67I9sUMp0OPFqsbdxqpW
He+uX1OSzyFhtH3nlyKalG5ITIs6f3EgXf5VvbxIqQlzYYiURWMMVwG+Sz2X5oblCU+idpkQB/e2
ssnyR/4K5dR1meNbGwRhYhjfaZCJbZ8e1FaJZvGdjq09ONOAXZvFYDG2VEFwC7Cy4YZXBTdD6YW7
fR9ftSulgV6VsAUQuAzC2gFuDNTD9MZWXpqGM0AopKcXXkaYKA6Mw4mEedhFFAUQJHMtSqg3T2hD
GFFLYCjdZm3gfpHgxK07IYbP039bbkpdlUK+mr46UUfmrWeV9b5lHG/ZVWZ1jlo9a1jIlCC87Ajp
Wo+EO2y6OXSMJWhr4sN9EpQncw6nixHF8Rk0f4IT2kBy0eEFVEVy+AKbFv76ezB4u+KjxxEkcepL
pkBbS29SmzJsHdYsqMFJOzlWK2tgfkj/7FLLTGhn4EesQplkRUxYH2sXDVTDGPPVhs7ujbqZiVLb
+ZzjEU4DgWAqlFWtS0a7uQP/KEIJDtnWBtovZyl6t0LoXqkYCep1pmwsaUkReAW67cXmaa6Yn3O0
q9LRaTcq3cXDGqxspPrEXAhDGQveunM+MS9LYG8gYb6CLvSCCH50GE3oBug6jhnD0Yce+yFysak/
Qj5BrX4Tq9KtcrCQ493bjW3dPuhdxQ/V7sA4R1HmkW3PJwm3QnJs7nfixGX16aTqXv9sQB6FKVpo
lWpl3tVv+T+gW/rxQT3xeiYeiWpQKpSLu3Of80z9cXoPG7wh2BwqO1XxfrmWCPmUkE583hHhW4+P
KB/X+e/qevSrUctVI09tzNTwZBc4SN6bEsqXSH+38KfSZo+g/xxpftiJmwEy6yTr9kNfePxw5sV0
ZVfq9tWbESo0FRiajQ75ECoQlzn07EqXSYmxfZyQOijGrlpCTO8z5D7HRaop2JCOpmQgXrgJlCtn
g1AJk9CQzN+Tkh5Y8nKN293hZedm+VlkW8ck4nooT+Cg+Xi4x8xEqfiXvl254IpGthLaY7YxkplQ
d2KReQct5dzOgVbihEVBsvgiGuuYOeW2vhZ/10AO2xdSW9fybfq5Fm95LYisE6xies8jGOw0OFue
k880oSo5zqWzsCSEsWbW2b3tEAtY8/Qqb+Rl5fi8DJYD/kujdtmpAJ1DHa3kryaVRhcYaNYMYep5
n6ZfE8m9AKcGyrpujcvhEjaJnGxYw8lk9HER8VdHYfU8nlIYz7fvgcQKjPGnZ143eLdGXcZ+HQQR
7yLZyeBMXqxfzNkUcSWPkJ7meLk9+HIZ316BRLH3gyHMkyhw6HBAVRefTvI0JrwXc+8Zrl35YoB/
TzcYmA9LqFG9oO8h0aa9CV6v9IlEmbXcSA5F0xgN369ohZtK5pLi1/rgJktYg4DnQZN5ycu4JscW
SfUv9DKxkESL7TJ8sgmbLGrziOUMJMiyGG6c1aaWkFxEMlgNZn804LbJptC8D5wfj/iMBeJaewDX
Fwnzi2475H/yp9/gt9W4dBQflSolQTfwYJTTKfeRZ9jtOlrsVLOtXL7rJcL5BoNUjYG6E5tPwpTk
Lr2uVidscfJOrvGSKBNigNjeiy4ZzAGomJlQVCDH++dDobboOMgaY30APr9ABz0GvgFVgKCRyeWD
pvRmwBHC5D/6HVrG8vkPtH2o2H2z8lRGRTeBoejXuuTThegQZGf1Bri0Zz9akqUr6E9EbfUJyuv+
eBhndlwwCC9SHAsUJBJxaCtbs8cDw1hYCVGnwO+qsGajtUSrGT7JGAQAKduJNDUfDwO1BgExz47m
yhtTlFfEc1rMi3cvKPT5VLCdpAVBepkFDInLaoOG+yvBafwSq8qGMJ0qE2B0NmbTuBhRQaD1SxpW
T5fkXSlE9mH+jOuqLUWOEgJJcJaJr69J45IOdm+3tLgsGRhaJWyBfgJf5r5hiGnA7volPj+otXU0
ze4tQJWIaTNrPXQsn6Bjcjn/eXJR2FpVQWDjQiWQsSdPSfeSey18fgfTDIhctnIvnGUZm/6j/PiD
XT4SjB26GrJ2cIAXi8QwMxJIz80UkSlbNokxWzXdDFqSC0iZn95GngS8Oe5V5gNA5lui8KPaUcVw
Ab6Cc8e9nS11cfhr2XnRG9qTkuWaGYYJ4d0uhFrZvkCouGa367K+7Q8y+HZGqo++h5qvR72U76P5
uLxU2a6D2sEetkAgoKx55sMtBuAwPOJUBOYapyySV06yEfPTUt2G1ow7lg9wSeBEOEku66/3Xrun
VMshBW1DAaOMzUxeR4o/nWI4F2hKyw8uZZCdEsE3hv2PB05FT4YCL8Fj491aO54mjWbGOonZbX9w
tdZXgRzs5Oj/cBDJUVYE1EhkfjZFRFk6RtuLtJmnW88QKVQv70X72uHPJQmjoDd07CU8iv3vnUtH
9AVoWtY7ChVKXzAjgird9Fdqx7yT3FYVPcvq6S6evM26Sw4yef1eyzy7UuKh4siRo7Id/VTZ7/Nr
vRRxXotA1Cjm1B4o+scY5yqbJNqCxGnc5yAtLwxQgAph9E2PNSQFCBOqtT+qFAMDQH/aM9qZzbwO
wQ8y6SoRQkF7AU8rGlyIhsiPxwMEEAH0V0xLdPSLD6BewGzWZr2qNHYnsBqh65mlC1Oqp3XVsE/l
/y8TXqIm83Od7xlNHsKsrAAdTrVZcO1GVgirStS2s/ZN+KdsXBlwqPFlplyat9acVWkTeMxP5KqN
Wt6RvtKMJTLYL7Xpj+U0QyR5h6d3vt+Njy/UVGR4uULdg0AklhOXRZ8aFxm8LUDZaDE+taY/zZgN
ebdPKdoExiLO5EF5WRQbdmDTbbcNsUlRjJxGWvcPHlGsshbQGhrs6cr6d9FQoNTh8UlrODuLKmUt
UXKGHxV6JOu6PlEc0RwL7+1CKS1s2YDOGsTOJiGQc420dYby26XgQ3i2b8eRAmoE1UlxXExKbkJ5
vC60ON41NT5neHb+u62k1j3/ZkLTxw3qHTzmgnhP+akHIURUWUh+AM9ssL5F92yU2PUjBjrBR3ij
qDkFPuqepFYs6M3KFq7OyHs1Bbw5XiztcdQcJ+WIVjJYeBB4H1m2Nr7thK0rWVDfmCf6AZSmcg7M
dMzg+Cfm3rK9phNHMiwJ30HKuIfAojGg6lgUmfGquEo1feTT/rfun14z2ACQ9bGjpHOnnLRdcYtE
GSrQ+BiM/bOofPLSpcEJ5C8xlFUOrnTcfL/cIxEAoyfjFsM/aVfoGJJE2w8ehKg38zZxrBLyI/1F
xP6EIElUOPUpqqoLxQrHcM7J1ywDAww0PnwuXcMeNb2sRLltCh+9i8z37j38pheBh4PrQm7e9a6B
dHlJyv48ApVWokkCjgmgxO+LhIRF6WKS57fPbYXYvUAYDPJ+R+mFTnikH5EFHN8B/69/3jXcGm1x
Hszchd0nvIrFCq3Zzt4c8czVsWkz5BnSLMTQ5Z0BwGcGfYKvbWI6423ZILz7j4DRq2lqjNuKyVRU
FmeQHGh56Mrm46+/Z0oeB4Z5QAnIdURN3HiF2gAfpt/0WgCTB3umZ9EFqrq0GhcJX3xgO+SZRbmd
tNtnBHOitapAi3iEcYNkzZ0NSZTfb/WpKYidrNbiFJvstO7ZDEwH23ZuiJ+do4u/etihb/cLcudB
FyduwebPayhwtuVZGNX5GGXnoU6Gv4hBrGgA0quypg+XsrJBjOwEYr4diRNxgjd3GHhNu2Mv3ys5
6fDSBsj0W/q6Hph5TWhtIBO8DFvTeuQBqpjGyQFhQ1nPU0rGQIboE8xNKVMrnYDc75Qp8I5QJFq0
hIdl+VcMIiSZUcSEhtUmH31f3dYus9omiGlRKXvCEmIdZ3zfGPd4GhYHWonef0b/oT9a57NwhLWS
/MjnpBZbducCBujbTVv8rx4RBhORhURTFUI2vwQK/YYX6jUNHoqdgzgfVub1JyU7mupNT/P2wbAt
IrP9nNRSLJdr6vn5GddMnZrdkXuU9nQR2q9DcPrwyvuoiPXi5lhyPt5xqlENRatHAMLo7uy/vUP2
zt+3R1hM1J25SH4KtGkcWz+xY7KrugH8mmtxv6NzXL0L5u3xTgRyo8vxQZblBNcRH0XN3CbtnaXQ
7cK/iZruiW2BiMM3wBtDJuPu9m9hUjYMa7F6on8qRII/sQv8K/W6AEFaSZ5oSpTdZeeBaTgxnsL5
rcLgd/ti14f1Z2r8eR0SxCyuiOp3WlXX+GAsT/+DshC2KfMu7pd7yzoVlMyJFcZ5WN2klDYoihs9
E4Ya/hjQp3ZuBAtj2HJgYBqHharJT4J/bYwFcxBpPj99B7zqT7nJ24FF3Go0akd595nlZTgravOT
6vWEbTFWR9ePoN2+FWpPF9GiDMLuTwjCcxXJktetC5PwoOqPXYuwOlzj1L6idckJedEVQ4pwqQq3
Gft5Dxz47hVTrSun+j75P2yVis5cBKPlchOE1nMqFUZjrdZRY4Msa6yxxZtxTA9u/um5GGCBJMjc
YmDZ2lUm2QgJHzp9rc0JNTq8DrCk6EJGC9yrGVfxzDmpOzjtyzMMkb5tBrrxdLH8p3H96DySQLso
sj9+sDw20W32cypWV+zD5hfPUb7GdXOkRiNwXk+rx7dEqztyfRi2WYxdl3SyWSzBs7DE3sqBcA2c
r6yEeUyqzhJrvBl+MH1f9oyJjlE4xHX9hesq4FV71iO7BF255tFnN85cyvTiFqg1vTtpk8mIAN8M
u/OaH+xgp6M4FonqqZeYprUV8moEqsXBy1F6lFF1pGT1jkEmbJ7Q30cMDX7i1A/ax9+VxfeDTEWc
pmobINig2gv9Yu6CjmS37ljvUXdyGXVrpmLhu23oPVAR+gzbGxC52JRzjcJD8+62a0fcw29J2zwx
JQ4nviuVPd4LcBvnOfE+iZSD9s4N7vCcfWPRFV6xFmZOE5XCnG8+mfwKyk7sAzt0s34GNDcm0IhA
EUAprMf06vzxuMtK1OjZubHTY+2IJsVrIno+RLiAlwRrSSalhgFDxzDqvVkPJKwqxduLAqiADoj2
MYdinZxgnbV/hPTcm3UqXdQ/2c8R86F1hYeqhDhMwzcyUDdeNe56pkfOeCKLuJIM9XOyVqHSbrzj
9G2o7OGNwmrQMTRu/vGIXuyCypcmfrEOdWD42HDKiwk9iDqVVV7BemngZYdQ+CCm+WM5gAOVS8s9
N80w7rUAP6rrOVni37SgdFePGNFOtLqTJOrjiFtAuVCU47ThZaHL65j7Xb9JSMfFOAcS+85HcE3U
NErLqoukPPp78x7UccJqMfRm0yfAyJUIJQdvCx4yTWW1WRp8Ku92sP62s9oxu54Gfm4D2oMGt3C8
JqpuTwjMqdp4CJb8Un/D9uop+nbVj1RDQZDLsJj4+SPhUlHtclXysKFZ5SnnPPwzd5SWO65AF0sU
in5EWS+cozTK0z4P/zg+PM1xMuq1s4lLYsJ4sfjWKxhtPWKK7E/XIvr3/5NTtm3G/POAP6OmbMra
ar1eUREDavQsMhzicAbsUDcLQgnKlv3TWayvLuaLS3lkutsScvdntY5nMJIpRwsZHFrGROOuqiSr
qi5zn1KYhsKK/j9/E+yNRPnWBVvwgMg3BRIRbOoiXC+Yae+VKQYmRyp8VeHJZIYC1b+73yhXJ3V4
meGI1poAnEM6izECMv/xaEdU+w/vzQSq+Ckyd/qAbIVuhitED543i5BRe1SRP2WeBPw17BSEOHuX
bVljslaODcPKfCVBSCkQGqzK/D6clSYmlGgn9U+15Pexb3J60saTNeIsUkpDe/wNPp6n7w0CHh2U
y+0EQzJCuCtire9SAgeXkrK3I/VqvNzgpoQD5FdbsgItCeT2InHpeyjssRmfdwosl7I0S2SdCWOt
oSyhGyzjUGL+FeQ/q4qmJZ9HtKFxfdx6+IOs4YQzEJSntrZviZttj8gkGs0Wihnd4FW2JOuAamtX
BpdjIP/XnTJZJA8MTeLWl6wI00//d8exHUPb3ZyyMjLmm27/tQ4yH3GCO5n4a4i8t8QCIbZTgyYD
3O4c0Yis7iEmyR678UPjmTFHxrLHRxaqrjWMtqLAA1TSFFeUtG0nlVR386+DIniTe5dfTx1Gsarp
tYr50bXzyCAy1kupCMCa0soSOI/jZJAmiDzSneQbFnrHSo5/V+lrtZj0OSE3cCjoHTmkps8GOCXx
QxNkFfNKsPLHBYckHJgabe2WFi4F7+7hGi9lqvawR6ZwlnmH/JCoJYuGm23+bZ4bG0AzI7qDAy77
2qCl7Y9CiFQ+qGhETPnp8CQOdWqqZSmAnP8eaZF2/2fHJcVlCfxkvBv2BF2uzDjujYvbOMAfX0j5
X3I+uFKfvgIJPnLBX777Z5NAHTfx9kpmzOEyBz8gbvmqVT1cubYsOjGkLrQJENOgKDS8VGu3spZW
WSQyV0V9A6gw/fFB6lrRtdPDC/YxuEZa35AA0FONIz6xMuhEx1zPU52D1jbUi+5JXKPMzB7s33od
/y6AJlBSvcpEiHFimbgVZHLmxx0/r0Qw8kFny+504ogKNRXQkxh7MNym5ll0NCmq2UcL8tP17aRd
7WOcTU7IiFcy8gJ5ikulxuO6SkWU2fHgAKyG7UNbpaWZUaAxivb0uVRZd5wUF3C7oe7VH8mGLTAL
CS7v76yH/7x2+ROTU+mGoj4+ucuiclteNcZ/3jqlewSgSQdxQD8LCQ3bKnqnDRiP25ox31kKGbPf
E7F17MSAJMfRg90Zja1OC+IrFnR/0AX+LEnwAkq8ecsf+X9sjHyTmxmLF6OcbZ910gs0RrjzaFSz
z1MyzrhLKD80/Bw7LQGM7lB94PuNf4v3j8tZojaw9GeHX2tfhjPHNUnN2SWDM0sXqjMBBOjnmruh
ofcStx8BIN7LzkTzi/o3VnT926WSRIaovFJ08XWS3WBYO5XVuXLw3ECNhSRosESea2vlg03uDOCt
+GV+2mA+n/Lt2G9z2FNM5DXL4pcFaGvNLFCUypfHZsDjYQWS0iKEXhMlREUbWB3DeRqepSsNGqhB
hhJkd0XjGsEH3oI+s6bRHR/9xo6utJL5p73hysAgUckHyGFVd/ZpieI8/kh0fTKBGl8PyVZZCbVU
3ZfLM4oq6nJzUuoE6+uV3ZBURlg57+UEoGu96w31+Tq91zoIPf4g3UzxTeSOnVFUQOL9J1Qoo1p/
QmRdp3//tESJf9OV++vISSJl8sA71MFpIfjNj3YaCf92iJOkxcFyQ3lTDRD2Wg0v+sm8j4antsvy
JQuWMWeZ/q6bT3zheamZJ6kazw8ZppReFc4pjzTbRpsiu1NqO2TUFban5/xemN2TInD0chFFkDvG
Q1MNQrZR3QWD4AtlgsnAoqV065mNRjQZRsiAFZv7Tsm+nzeB9lfJfjyhbcA4Iol+XQdDFNbEQLym
c7gyjtnJ74tZ9NQWh3ZlujxzoY2EmXnd8Mey02iUKn2Nc4cl8xm+EUznaU60NGGvrix4c8hXyujG
L4M8EtTwaL2y9ES2KFxjjQOhCOkanCpe9m4iLkmrPRYr8IPQCQxErITy0CtDMGYE56JZGoXLLY7s
l3Mo6/QFWKd+GJZPOlnyW/YMPAyoJdBUNf08FSetr1C27A8BETi/YU4YIuR7ovQwQckRYwBBcoiq
eK6solqekx6zfGW8IKIRciNOFk3U9qEeG43LXL3XibTe4Wf+Z4aZ9uxs2uOP3zgig8Y4MAuLb5/s
mCFMYlZN5f9dr2NvfP840xC7HX2ubR4Zwc9nL8uaPc+UUVQTtk0nyD1zpPDA4i3Gcb2lqGdSLNMv
YEyrYx6xkvumYrYFzVuwZT6jr0B5YdZjjkSGOM/BHXjNPfUNXhoj5xj43bhMIS0muXWRXoTRSakz
O7vO0WMaYEmdqehqit1ewcpn1z44G157fj9y9nrTm0xT/wtWOKkb6M6tkgchDo+9b93ivzGcRN6/
rV1IFLXUXXl4DR0s6p2uKBHBdt99zoipzpdGaZ6P5IUWqxbUWj2uKTabXODVOdUyyUJgZ/EBUKbq
pZFDwPWY6+0lXyXZyEY1hA3HWvnqqJPGyzawy3CQnhNwuYWknqfW+3EHEKRaQsTyzI3VgJe0O8dF
GZPQNJc/eKE8MqYnrvjqxCObb5d+R1lzFJiSj8i0W7xJy/SXPFZdxcm8G/Zd1USm3OUwGY9XiqGK
uYbDYKrgbCdsjv2GYCoHqoZDpA/HiKFQ7p6PHzOMZY3Vbhme3aRCHw7YnUJn6T9fcn1t8nLfJI14
upeO8pCxqCpy9UJktX5bMKapE++CSsrbDbo9p+rjMHuIluuy9r4lvAcDE4EeF2CNV/gI4DJG8Dcs
ZB/PfZGk/XSV6RWRHUVRCxQELZtty775MDSShjlcPCSVIIccND+hALUVqtOzVJfpFROS7XC/ZaF2
4cqYzyP1eO4K92Up3JzwWLUCXAl+YMlvRRdGTjXYvO6ImK166s/mSITiooFMY45Y9q2vnfgDoX5Y
mqWK6zCvrs/IGzpjTY1QE50tQfDR5aGcNPy4KrOQpmlxYGdNN/g/t+DR0Uy0LcPlbyHjoak6Gv5t
Y187cjKo1pQBDh6EdFa8v5Zawk1IeajsB+cruuUIFDyj9F1/5mhTLxRJnYV/Z0j0BuYppQDj7c/Q
fvEVIkXIAE/prDdHrKLL8kElOK5AN/jtBwYWM1diGFtX24Bu3Naw2T6vSf1WQ6EZkcs0OafgyBWq
sjwTXTUR5r/kJ6ziCyqkN4K8+eWViRkK5isU33VL3JG3+az1/6faQmBvPo7pBBr7qPn4YG5OEg+Z
nd3BQmazorE31hbwb3oKdNeflfQg37wXy4IfzWwD1LFLKE0p6uLf9P1PVSXjKXuSQIhXoGmvlTrc
qLwS7AUoAfJ+0Cn4bqQX4AVhpmAAXvs043aQYtL1Fm6rbQgs243eI+PiLH/vYeJqxHfP213SnIO+
EONkS/vYBm4+ipimTOlyV3jfCstZIStnw37hgesfAVZH32geUgK+7UoLBWtPKDH1R8Q9PYYqoRxL
/u1te9T/gIMFK7rdM+rosIjjG/tdGGO2KImarqernuLs874yb1fx1pdJcMNXPXXPohYSH2oxty1w
NwkhsAaPuHbO/fVmyRp09L3RMtSvYmyg4WhveP/r1oeHsnxIoTcqjrPyap3WqQSfZaC9IaTye3UX
U1n8mlqp0RVETGwnEjMNupmkmrCMzrMs6S2Y85CoYqUOl3S37FMtjG6DShDtXQ9GBz5QW20nG4HV
GPYa3Lk0vEHpMOddAL35TitMBJsnCdZdAp6g8uUprboCWeXkeB/jpjA7D/g0AhSD4vlR21qpaoDk
zJwctsb3buP+wG3egQQ9dhHAlZQ2d+GN9vx/kZfHES0E9Q3fgyJ9T10rL2aI+qw4RG4ECPN/7MoA
qBECSBAI71ArD/H3k1AUm+tRhsa+n0x3CsAx6HJwwG0LLq4+3CeWv3Cv7e6lewGPA56+GcV6jF5H
nqxIoi+oIt+DbiBFwu4Wx8eaRSXYSVjTzSS+EqzRrZtbl77QVV/g8PtWNRHLU/xihnnZb9xyIUTN
qkCMWdFKlvk/+ks7EoOrJcf41nExgMfuREXsqrccC91jpAaoDuEc9BJ02WdUA+B5vre+SyYeX0sB
pJ84Wzje3Xgot0/lmG1H3Y4Xggw3kcKqOXfsX2WC9nhzvGxVEdDSSc8DuObQ1HiWTg/4uwkbwW0M
1M1zbstYBA88InBL+3v+jsPb2oWWZkHHgQ+ib/9uVXSn1dn4m3og3t4148JwgUUiCxf3A9HL8kuq
ycNcX26amFS/XvBYMQljQjsCapls2ZGd0g4FaGxdSqtrpMBRjwPYoMU4ACzdFO/OtlzGbO06cFaI
exAGecGsOVIbh5AJdFpRNQkU5Gmx1qV+IqF0JEGaXvgI/bJn+MpAFf3hfH277CMrLwkhkJf/6rXs
DLL0Ti28TXCBkWafnYHm6pe3q8zdY0g2Xv+I9fAJZnyyvIwatqDNuIU9Us6LV1t0Kqq25QP6gKWK
gr1GIGOYXWpJsHOPgoMg5sH9P8aKg2VK0EJ9wHkf/OPJvR4/V03WHNLINn2y4V419dUr94MFSCxy
ZqJaWjogcORSjjCK4FK0aO2GpF9kRTz4nI2g6+ADoYEI1HyEH7+de4/4JxXe8v3VOHbqmzRTsmuH
mBKSNAE/+tnc91If8ESC1SaOTh1zjnAwUwd2TN+tqB54Reo2ecigKqntTNn/QOSIPcvlfXuwInuO
iX+YjIbPK8cTfBq0A+3UwVGx4JFmZezA/7w7rnFgwiSBUfY95E6sDnlbMjL8WKP2HXdjKJInUKx5
+rN1rl43U8OQRAPJ+SbnyEm94PD7M9d4jJP3EwI67nHRgOUQEiKNRkQmeKWVSHxnUlb0zSdHmLvx
YMFBs5TpnwYUn8GL32NeHmbvo9pyhqZ2d63dc46ilJRCJ8jCOy2qORQs8H1P2/DN+8zYeNa1C1jS
NVh4hanQVqdU9bAXGYTD9dZgC0QZFZO/18/NUi7ac3DQ5Y71TF4+7qoEU0GW8rD8tVueqceEBYmb
Z17QrMaiVfxSevhc/K9o9hPKS9R4ylGMqUQE5e/pbtVsc9R4w7T0cqUiNFCvmYhTqkgy2D5LVQ92
RshxKID5iWI6p6QBd1+Mj02YmgLbXESq+GxBg1oLC5uaYifsHOuw7kG0zaCSuIcnJtudL7aYLyOd
E2JmPTTFwFY0BJo0xlJRysJUW4T8uKsl1hVlcbKk+RMVgkFg0PdLRG0IFcGHH7F7fS4lfvNsf3ED
al+CTvRGiB49JlE2DefegWLoFSr91HjATrPSR4ulQ1Z0Y6sX82ic/4q6PdAx9D6Nl/k3KW8OCk+D
CwMgRks6qcmceN67J/eGyC6y9Obn3b+GGtupKnHPqGFoPG5UIULjNei+J6MRmuldbnd7GGJnFmFv
aaOxryp7O+N/38IMxkAPnVkGicRRU3YCuVwdqeXoINls3lnMCatULyL6xGPwh6bipBm/BYn03Mho
LspPGHo2D3cCD0yAB8mvuyXdQpPGpXLELwnsLgEbqKwcNS/Q3Da+J1JnZrH+rS1J6V6rvXK/FUJ0
nd+MGdftlWeM3KWIsdYiWyyOb9q498cva29oKMrH+nMlApG1/7mxrjbmzc35DAfpO/HZNWNhPtHA
Aplew69DG9nOcwVwxdjWbjzcO2n5kLJG6r9S78H7dwdDKy0VUpByhQA0GZ4GMNxxBJxSt3ySYw5y
jGtKRa9nMaXwiG5zC4dml+9bw8QuUeJ6hSQ448FUaNQ5g+aeityYBvyCAYCX8katHKSV0AkCRnyC
eBCISUT2U11xYB+3DqrunXaFCvM/uExziOX567KtNHJG4XDD7NaMDMPwDLQX57xVKKhP/Zar7F1g
MXQ68v5Z9iCeH3jdOv/XfD6ZLVtyYO/56ek4wVPk2GDkgYJevHTEUm4h5xeEENIimKSI7IfzrNZ6
JhvE2p+22dZVS3bc0svFXkdSGcOTtZGiMSSnOplclV2y85izNWXiQtlJFMB/If/KP6GtmRgJ3guB
Qjf78mwTEYIT7ftlh8bkrzkm7li5lkjB5djBMIVlcOJa1bbmv6xz2FwmjVjwjnuQ/RS+6bWkEDj1
PLIlm4x+5aoAvd/2nJN7vMYLv2gatWVZB9j2B4K5p2Z6wJ+GBVBteO809ZV48Xb+/8SFHYhSvws6
JDqYWzr4eqe2t/g1PniAjT4+5Fb8rKNnw+G214HTKAH9S8HVSMFra46XaEb/hh2Ao+ptHhk2aHkb
QGUNFxvvaZoolgqk64nnkCQxIkW2IyjUhMejae+c0eUu9ZZo2keB3Rxe/lvQWOqczvQn8ux6zpC+
+jUIddLTAr46iesF+JI+imVI0Vo96K1KiFMY+2kXJGNmxbeW8HIsJz9kloO2Zk9PUyLxz2+7wFNg
8GVe9Q6EDJt+r9v7CpuEyxRGtpnFhxAhii4RnyU7xhq4b6XiPJCpTLuHKGcNYdOYRL1C6GH7vdZi
vDJfXdHlFTOiS9VlnAhx7Xrx6Ks3IPnUlne7mrqxTNekQ9/WEGo6zCz9AJsFiM5+B3qgFB4qSvRD
l6jdMdcZIIonqe+ekG/ZDWSQFojdmjVXanZYh1t2cLp4Eh974ThxuFJsylYrDruftsET1SR0l23f
OrOKT19PwUxvOtIA3xY+sre5B5rULWQmNJ6N/Q8hnNBWKd5ofKOltxz0V87B2L+3BhZbNSCxoCTA
kIU1Oo98Egi2bFJ8FVXSc18TIWRL1Eg3vR8MqfKbiivU1cc5uqJ+zNsySGTEzeIN0fAOgZoz3D46
yklRC7y+GmONpiEI2HYyUuyGweo0QNeVmod4aEYP3yNq2UbzOyF5PYWaK4DF1nITuTOsy5zBnLpi
TLEZ+suJ+NRJkGvAhD6xWBi7HzgTi20qPFLwf+wEWUGiy2nizB8Q4cQml4M5dvldMVfseo/nYTYk
Z85ajtIfFLVUXMpZ18WPOPRrJMt/DIaKljSpnkppIgxGox6TtXXapnqJvbbOyj77YUdPUBe/+9DF
IPHHxE4wuIPTtdSQV8P4vE2ajaTiAnABBoRDpM4+T6vLfmHSqSYBaBuUT9ndQrIeoW7N/jSkjj6i
D4qtq1L5EKCxYEoTIAyQE2jYh9T7m/YPM6ff+2ldgTHkMoMVqDnmPc89s2LMvnd21KiDBTxnIPO8
YWuavXGXlxAcvzR7iAqaRKgK+mng8daB1EcmBJS3bJF+ZHf3BQBggUJOcXoGvaogtDifHf1+lA4Y
KOUrS28yRrwL3w4jQ5LGYuknAS1OsN/CGORfjntZgScMW1k9VCMQk0buVGSKSFTuvQWpOCHTMiH/
bW4oVoCkYqQwatoYz76ITVqIqxMGI1J9kbn+ebAdFfLGlsnr1n4t6Z5pxFvUUTCB7bgqTq3n97D3
E91jMcuZNvxmRzZUEPaJd8sRyc4cJXrKtFnLlQKmjPLXZyLu7PmBQkE3ocsLJrlVujAjneUyI4qF
fBlUYNXN1h1vL+FHoZum0y4OsaowiEsU6QBb67E2emsTvLrSta+rbQ3JuLyq7IXDmYeh/1XUPM68
nCwmbYFI8kZBkC5RO75NkXJTQd3titvJUklvVJDC9clBzYjL9wb6cB175ovqGPhxCuHQUkE9CDqX
wvabhXx1w+Nl8CD9qSGBvRZaQ0ykygfsRLysH0+dVZ8G8F6QZEnsmLTb/Qk7tpV051W20VmSW1zz
gjZgA/WCuFZAaMRfRWeSKCPzCGk5edWAHkKKKlArQIGdztJpWCgqEK+ks2KTBnieyVKa8bc3kvu6
6IMtwIg9hmGC68ifiWnajj5dHUDXuGQhYzdLUnMw0j7NVdzBLfKPdqyYKmI02dtZ5C3ljdIgs2ZP
FiipNKlZPSAopoG22YrZorT/uzegbzz/E14vGlQ7yxexiFkWugTG+BBUrkQzE5DK4mkKCIU6vInF
Eq6smovmolj2QhsD5+29WalrLOXVIh4ZWRtODOPFO7Kmg0nU8r/DO8HZ13cSgtwI4z4R/RfHTd8D
TZ/3jQWhq1fnlY+LhWZ3IDhyNcO8fbjMNGc0517gWReskHwPrT8Av3vZs17Jm8Nhy1dyFf7ivBlL
D1QAVgs1xxoHEMhUeWIuy0SLtTDu/3kLTXG96evO5UyLEfRBxst5Q8JsX79Y07ZYX2UiTFcT6to1
CvzSPD+HTg20QPBOtOudiH0kODoicCDHD7SLz56aAUD/LjYQ+9tHDKKrlN0wx2ECfCua7dxyiESe
meDgrwonwPG5LFhPZNk655EQ8CUHyKZDcSJL9oKRVuceyJ6vMhY4tFOc6OkJ4ffSLKXVbPp1IKYt
uJB87rRKlIjRhYuHzvFWu44dcODtKFtXh8vXgarlJzJBpcTAesrPCXMdmdAOcvGY2AqoWwHxc6d9
v5udV7ONvDLwOjvoaWGVh1AlYD63LXy4R0Et8NUoYLxTMHvaOJuZeE4y0dAuhuwkWHZWxRBAIuh6
Caf/3DCH09/Y30ocvm18TUm2Y5TQWQbQ7E066Pw7wKj5XPqWLNcR+FCHuh2m4dfCFG6Lsn/ZZH0P
BiW+NZSFSjvZB+IcwJzicaj4YPqb1tBN4O/9yrUbaeYY7gK3OQa63wTmk5OPlSJVHF5DZJVcQWoY
tK+EZymAhCAruldXapyEsDtnLQBvPimt1GAUUV51T2yZ1gzewh30nMEmdZvPrczdfW+aZ1vKBG/h
+sDyZ7eAv+AeS9+msjpEZA27jJ/IgW9vuMWJS3gK+HEj1L2WNjSNcWtqfPmb1eD3pXWgw7B2b4OM
kwKvzol3aKgGpTSuCfQp3lKPB91A1xjYummmXNn7zrdCrE/lyT0jP8Ok7UqC2bScSYAc6hjBpjlq
BOTKA1a8Yrq3vahQ8q86Ck0kHglSN9jU3Res8vUgof2IweHG/0ncpjxPq8ikkTPiJfcTTrgMHXcx
m2BD4nyMnDmMpa/1YYf9pngOX0gsEsS+mc9knNuXo9Q+JWv+h2hhsruhijYUbn5dOz5nW4ttZT8a
gxBE7wpT8oSog5b5MAs4FZMrkUhp1FQSFddQn86e9aWaTrb5eXMs1G4PN/gH2MIwOwqCs2WTvOC8
1EXLa/B+k23lqtGGt9jd/LAvOesmpEksl7lQm9bj0bIDmTxwmJGtlGYP4+WWFhEqBeHb79HQQv+n
CkS23jJbeRWd24OEgEYEo5aYBBLFRePy4ToFqDrOriso/lTpye840a/UDlkZ93uQL5paFx3aPBmy
yqZbGRyJN3UQQ0aZDY8xa7wEznIkro3PN/ymL+hmJoE52lgHMgPDrqx0UOc0niDRik7nYZwYCa9Z
Din+abLQ/GVeeiqW1n0qbQoJjLgR4moLFgVpKvUgKRaX5zKpaP8isKCOzc+ETxTNKKM3ee5eZNAB
YIrof68p0elU6e7OQLsEDXEXL03N6eBIo1+4aFwF91jF5oZCR8yo0YJs/OyPL4LBAU3MC85A6/V+
vCdjADCV+9ppjzMTCXoEBgSuIppMYfh9hOIx3Idfrtsbv40W+i3QHBc9HqhrEw3pe77pjOeTtMgq
j58sg2eMfGN2SUZCE37mvr7sfZxQ3WYjmjIWDwvA0EwKx2TtQ5WL5Tjk90oIzD3joTGDFjlCb+FJ
JF7Fx9YoppcTLCtHZrGhHGpN6P9O0izdStRlinPvDXiVKNJr+dcqhI1ICiAIta8iv4L069sNJvXU
qfRuafTkS7GzQQUFSnWeyIlLKOEtCAI/OO5y9Cq8jt4LPemXcmsisgm/TXLh8VlFgddSPPizrbhf
FHhF6Rh+3XiWbT+ycrTNyIyH8XpcsKqqq6OlsmJXCu1/ZI6S4JFLGK571gA06oMIv/1Lg7EK3Imv
c9N2Bt6uQLFmheNVFw6XY1S6H8rdK88Xe5zpxI2WtNx2fSszugdTJvdXqCxEGg2s9LKpAgzhFQUC
StB4dXYmKlRSSQiwyti9FWBUZ6TSqqzfvaDoYKodeO81fVFXVoMXk//fs2B6mvDNzbTOM97LzKdh
pLOpdfIzCOEaX6nk0qyMaDsT6VzBOJr0bt4RbL/lCsPKQTURomf4VXDntnjawlSjV4FkwfdYkCpr
hMyMsg7HB2tdKoJtB4gPg5xnchxYnPOY6IBRQzbrGRy02gStTDcO2gWwB1UFhTRAYAAcN/M/6Sb5
J9OUJplAnQRfxy8pGGBUj+LUe7tsf+nPYAfYc1Af06jCMOmNZgchytfRKEwhLLvxw2T6+NdijYd0
HCyae8Xx8Y+fkbADr9ryazWaasmFj3so0zGKt1dogeFgsI/xP2WllFUg2tTOM0AKt16TzmQf/+6V
Wvuin1xrWJGj9swRsPBa9uJDqK83HFGoJCII+zy72zGeDke29D4ZvAu9ogHqCBkRqEzWXNURxTJb
cQwoJdwCkrP4ZEPaigFSNQnJt0j8eH+MrySreF0bn/y9Jg4y9j4EziBM24/DoIvLDyskqXIfxY4S
LUCSC1xpa2eVdnbV++5T3PCif28mKMQ5h4nGJjyTArcrCXjvQrkoQ4vM43IKOX9Xzlfsbd05d8KY
Tc0hPT2C3PI/Nyvj0+eLJGXWJLrh0vPUPI1cUlB54Nl3w3q8AzVBST6KDopXfQ4q2GhwN2cw0Fbv
4bpquqoK6HarIUFYCmGt2Y/YOZYhHniAUr2wx4D/amWyy1tT6jhqt7hFvrh0ohr9/35oU8k3Z+ZN
oCBNfkJaaacMrdUIlEM24ff8wCRcUevHHvmn9Gnyc9Cn31xSf9TpGxKuBMtF5OqCB0Q+1RDs1yQ1
1/aOierEtUqAVJRgXJC8WAGwpmHn1zcuSxLpYuu+neobDW2CXax7yf4kvusolKwJUE/3ZC9gNoE5
5hH5VEWbzWZASqBzDp7bKo2mrE9Cy7rXzGKHPHhwtKWVt8G3o2vi7FNTiDgtjsqhGiANkYILdQzC
Vrx2W8w04GqRSvKLjFLKrX9GDvlMPM9Ji91vyX0Egwd8hYfq4t7/LwWWo2p/932NoNYFzr+i//jI
wqQTCocHxy7GSMLLd1zqyCgusowLQlQE/kn8UfnNHwLyLaa2efzVTrN+sp+Dd10KkEMI/Z9jHJfV
BuEVGAz1p9s8wyjJOPLWMlLMYE5WAoxJsMfHiLzY8vTbE7xzOMJe3na0OHxwtbAjgMom+OowKQmW
1aESUc64ljTr3uAcoQVVX+a4ugx/tPK2I3y/UYT5tZwTyHQtMbMoIqCUdXcBX7sl1RWAdhXyIYhI
uFBXrs8m7SXJyYwkWroG3bWWCJM+Q2qHR7VRgJigbRxnIJeiUo0kD1gMKa+XXX9Nj0I6GzP/3Y6i
2o8KdGYqKSnPKk1RPmDUSbCJFipfjVrVlE/LR7b6IYSwxZmPeVhnu9KLAREd96+wsXS5xYWXJ6/I
IG/BOgKGuIhk+0d3cHN5qGB5SEbinHNnwfEmJ+PZmtlwb3E/g/YUj0uhrUUh4sGVCDHIyVO5SPyx
g3tbvtbaRm2GX4PpJqxIMNxvBre+GbNfrODYDItlfzd081bymS6MsRhfH2wId34poKQQlKXy9VQ0
KEieFm8FzNgPGkBHgUOIBvIIa3znXJieNEopUFo0K0WEvfHduH28pass0iYlpqmaIHl6QzYldWEa
A2odYYgXZMbjyBsLzcPDePcdYhALl+I9aG+44dFeG+E094lQVl2M5mDrOxLgbr/KbW3bOjNgdViw
8IgspDaRUB42nMHEJ+0jFnh0sLv1CuPfwsuea7WSdoRtf4UwsjqC6VK/ltOj143mhNzJFgS+n3a5
xR8TAain9AkNeG5Duv3PQ5THrKZOeBnPbv4ypu80W/QwHR0jUrtf5xFXgZNu6MOe6ubPVB0VTaF4
WBSHmBD36KGRfUQ9yn5cJi9MEpwfMvfzCbgizcWJRbJ1TKYyC6CvzHa8I4vaY8xQunGagnIvgxXY
LW9RdoFGf6XPbKP7uTdqXpwaCjQ4lUOOiWRhJlsRDYWttOGoTtdG9y1SwRB5ObjE2zOuX9jPhCMz
1wM1ivHazfzQ7hwnMagZeXQOkRl9SONYfaVlYdR4lZrVQ6Iif6noHMZ02HvkqRsz6PucWAdnJmDb
OMCMAnQVBgLM1LSfqFwfBmgoLkYM1V407TDon8NvYk835g1TDU9nOUa/d4HNzkWYbvVvkjs2FN2D
5N0RaYb41dek800IdFGlYTZpGZb/z1yHsX+Otpab3BQq5yt0Jd3YYORTQD3/h4y02kMItQ7pmuxx
upB6nzouHwky5qTxI8H5m7gDuibG0Ce6Flaq2GAYoKvZKNtiYvODx6Z5y5xwRHf5ZSWGrr3BiPj/
qNsdYzXeIydyeDVH4qlDQMC/vH9h3ZDp1GcfZM7LP8XC7/iDQxpSSV7Z+/kvyIJ7NJypDh82WqCN
8Eo59DG1pRH8g2ZtohZlf42JxJqcZrsugepQYiv9Y7Svsl6Fbq1S4qkyfY2gX9wwAlAxDUH4Em05
/wqYQtLJjl2g859nQwCEuyUM5CXHf6neM+YStT+lcHWuFrIpgAPczgpaynADihA9jXKLsKMHK9Gf
tbZTgnsatKWEj0m9pxDRmTdg6eVzi0AzH04n6rgjTPWYvLKwThGWTlgvKrb6U2EFVxMH9NWmtHgw
zsmIqg3lBywz1EPeDHhmqrWRtvLgyGo48eBErx2in3oJsDCwQ+xgSg+S6kuo6E5VKVft132Pkylm
Ne4QU2yuCh8BdsM+jcgG9jc7vxlXjWbgfCYK9at+WwVIp1jscUqReZDDcBmbSLeO7tF5pdTPFtVm
bP4pWf3zmqIaGkgopq7ngTxpsw9TGUSIqRGFSM3PZl2Wk0NL+QQp/xCnqaOo24v5CalAPPR81rBj
HmHx4ESf/cHfJjIuEqQHWy0mCGHWkLC+XKj+skuT0A9xrpjC6O8nAwG2FiW7VWpsblQaSOxAMG/f
5iswtYSRR/CksiNIMMritVJLY9pLwBJU2ebdwQK95NQMxgEkiQRgh4MM/JAzusgMQ5x0EBb9hTYi
q284XRrT9JP6VvUq5QjjFZ6SKHWozzTUe9wk0zKH+/dkf36EtDbj2K+4FzjhWGl71yKehsQn4jLA
6DvSnBl0hXMmdU+Pxmw/1iazAD4sqZjO3w+A5Q/G3QBJ4fw7HCMw1lavQ86zFimzaCgE2KXg/5u+
F3a+zL7IjRloWiqfM9r40+Enke3acKH4l8E05lHw/NoHCbIb26Z1bHBqOAJ6sN/zJOn0BMC+p3kN
DQFVAigLi8zL67WBPsF3Vzp02s45SPK56jGTN7XkmgRM80YLtxYCr/S67VriaES4UJSnFrzNt2wW
TRKb5tCQl8BAgr3Xjkc9U/zXcF+kEKrjz7rZrfYEPeNxQYYrOZj0+bFix2jD535WJwuHJhx79vtj
LDknmPioUyzw8IjRIwstjm12PRXXxs0etqvAi1pfLzHkCPQQTpc2eEIROKgakiPu5uCaukbXOj5H
4aA75yvWjR1eW51s8FNFrw9BRyfYLeAP5kpsxnXjKmvw+j7SZgfmP23/Sa47SIOc9d8nH2sDZwdd
xbY07XQ9skxBY0/FCTFvbJU3dJnLCJgoV/MsA9fHL7miF3H9Z6/GWf+v0st2q1qXVO/21bgXjqbm
TZXv2fZojNaFRR/y+l2OPFT9SoWJccUERYFervrgw67HeKrQCR9sFiDGBB1dp7RBcHf69sAc/QZt
b+Hgg3ThdRv4O9yhbmBDFlGW7emlqPKh9MK4h7UGWvPmZ8jf97BlFy3Oby5wL9zz4lnNvLyDLZ4M
aXRRWiYPR3Ok7+Nvp3jRpghMub5cIt8cqegK5tDJZpSKw1T9TLt7DP7MmDkMeWajRl/smsCn35E7
sn6QXx4UtILb7HVKcz1r7H0oM71qfa62MPxeYdiy3fRPhURUESppx3/oRBLo0GnwsxodAaMtvRTB
SP7jqoSXB/VcOh9iDlTlXUBg4M83pi7COooY1OPQqdDleeikqdMVcU+YR+JfiBsyQO26xGzBJs12
DBiSr6EF9cK2Jt5/CxcMbjBLLQNMtHbwRQ4srz1hOMQciaZN9NMYuo6EG13DZQ0vAgp0r/6wQDbQ
spzZShh0BeCeep3dxgPfveOvII6t61c5+ShX17lpofF6Y2wvvDURYW+rmdBkHP2Oh46HUuqIfHl0
ioGaDI5mC/hOsEMc7larzulMNXhKBz8AEOek8emzxCsWze1cuEXD8HAf3uwvWGMP5bFboVk2So5p
xVbm8p1QI8W1MXWjthLElq272u751pTaAS7bFN2rEs1PljkbSYoQ9SPpC5L7c62QVQkFQ/DT+sFi
7RsrOvOlghel1ICBhSZ7Mrn7trXRqztsWTdt4mHPeItrhaoe3Xa4qpwLhw8SsXr/z/go4bQlYi0S
Il6dXuV0Ae6JgrrfYagi31mqwQ9maiTmPt8R0vZWppe/uokro+CsQJC/RpzIhKZ8O7uI3IS7oqXu
aJ9PCOQ3qLf2g9/wJg2edoVc67FQolFAH1NROyIHb+pk1Wu159bvnBZK6PAErqRBlcCvUBNFWNag
Ah781if3uaPJ1ignmO1UcWyEecOowgask1I3ARIhqi2iAsUaZQtn4qXeKL6IFkm6DUYef6PGPrjR
9PqreRalyjfu9KoDZ404Pm4jAnldjyPUGVxU5/AmqSHBy3JyUdvH9vUvZqXUPp+3Ra7QMGjzlmeu
DlnPFCDD6pJcgmfa7E6NxxI7NnqPXgfs98OGGfM9b4Jy0qqIH4zQ/sXJYFvFLGCtXKFoGahfQu9Z
MstzE3K2/YkIBvcjZt9TYx2IrQC0kLI3MaWICVYFZHwu8lCNv3Vt4bmnHcfrWDpIGOsgiuPbI6mH
HT/qeHaPdTslTHXyhIE2VngrXrnh+8/C/lYgG7OfLAd5HE6CeVjNY9Ck5TpFW38sL8RReZ2H5ko/
Ki4SzfAtP1a5BDUUcYYwagWfHni9hdOm4/GvBGPgFB/k5t7JtkU14JfyhTXv1s9zvW/z8Iib6Dl4
0zQyatW0POlDEUvknZb1WV4BxNlfSUgWRgC1CUCIAax5gESUudKIAoF38QS3KAThEsrOtMMEKL+8
itZzi0Sm6UEvL+07nWb4NuQqaSoF7Jphz5yO5vUwPBtZMNJ6pThtRRebkOAZLx7me7/H5k5QXHfR
WcnVFoUKP13IJneiXUA+DSw1ZtCPTNtXQsP7IsIZu/GWQyZ5EQ8nrAlPMEG9ugiUz2GZVq4rLK5+
SuKyEq1VQopZNzKpHkKu4gWTNDuvTTrv7bhq5Abp6QWSYj760SsP3H2/tI0wfq+d3CB4T8Oyosmr
qWZ7VkYXTTsjkE4sqkHRlLKGVRlRXVVJTwcX7Rsbm91TDrmUI3RPs3s+poWsyb8yN0YHJQ5d/zS3
Dn3bi8pxlMcunyV+A83RKx9sHCocSTX6b/Dp3aLcjDF4mLYmUscNc2tQU/B9YBZqoUmJHGNfHyHt
qbfWuy8eWBTMJ1kDkMo7gCZmMhd0+obIO4qTwpBnZ8Id81YeGyG74BT5GhTzvrM9lXKqWBjckbWK
EgiMGQlQaEBN30AqbCSOSPYEHl5+BitIJscYcdRp0NDfhZY0NVQiDC+4ICiHzSrixmqXIUVZidci
V153WTLWFIYvA5AE07BeIDVFoorSnM1Nih0toqVRWmHFZOeCMkbQZrfDa9GxESgU/I1Cglzkn4vJ
a4cQNcgWeLJ8dIcwxEzV4dNEJiBEXpBz0GthPrCgI6dGxRIz92R6eEH4U6zsU08HvuhuRDY5Ay+S
OQMH657P0FlG0wYW72dQozPiL9+GnCfY+yqMIlS5Wi93QlOqo8htLKPeFzue3DNCwjZX44FKlqbU
t9DZzrng0kx43VVEDN6Hwl576BYlJX5Abui0ce2bP1ZktoSth4mlRR83DYU551Dg3jt+HQuUROl4
gC6a/VvZdF8i8hq9l5WfDuABy7t3imS6gyf+AAa6ip1hoW2bzQGtceMVJIy0SFmfZweHPcPj+mKf
hFu6NC8jypmV16wbOq1/kzvoKbXtnPgxhYqSIWceDGNV8N0hr/bdJq1OuxCYUiMIbY7v5GTB6/MS
F66iuntL54kSNC+MTj5lhS/k/YgbfVdqY6C7md37cDqlebs9lQkBxWLsMKYrjoSIuDuFz1ZIjb2w
KwIRCkoiyGKsBndpb1KBc9E+s7a3owe5KCBdmpZ9blqfPawqJ4D9BOfWAtOBWIt5pnn8Z6Gssb13
8KMeuoFMiDB/gR9fE1RPHHKibAtPxkc9XJKpCMlKdlcJqeN/mz7fwYJJu7A9b/6v2WHxKYg4fMUl
rJSVyypi+Xx6gyBai77xpT0VSqc37/AABacMm7GPTZCDaFs2V6SHuC9McQ4y91hwhy/dmzcue1GH
tEUeBD4WdXUkWcvQaoU2001fVaNJ4KEKxHJYiB7e1rDTkTX/vZPaNM8vGpaoPX5xd5iW1wegLgVx
IUWfybLjyaM4bWKpAXurk+otb+LwZGseIM0xDiOzPN08l08zMGRimfgwQqCaTxJIbYcTAz5OBS4H
0DBn5NW+pygnfjzyTxgP1OSXMbv2XjC2ew9i5/hy1UN2R4XWIGaHlvWJETP9OmjZR6yVl0etED7K
TbkAYK4ieaOmqwl52taFK4wsH1NbnWkmK5njWBlF25khiRYiRvqplirjk9sgWev3QO3rL9ROc5JD
CsOUi6o4pyGhMSThXGCR/DJOiI2C4QDbOTYZrYxOMlaq6rX+uq3/Gacnhs43j7ogpnQhkG5FSLRw
Z4wokunX6vetpL78BxOo6lNlkeaqpzI67jtKMHFmX6Uo7cLy4OxxZPOM5efmdldJBZo4JTb2HWGh
uK2X/BzoUayjEdAXAVuhrNktADCKkZ20WlRoXeFFc9A55G8XEdW8yXjXtC5l8BfTcLi/fmM3MKmd
1CHKU436WjIZzuAUvXjiolD3RYLcnY8TVoMuWfqmrEzq4Rl2smQNzZaPqAAGagveyRPjGmf3FzYG
Lc57EF/VQRK60F7yQr+psFCwELz1UmVszq3ImpCt/srghkRh1pOYYv7JYhpIFzbkvebo3e4uRXtC
CcH9tkkNEKVQRlen41sXAtNmQQD4/Oj2IO3YpdGQXR5XA2b2cEAIyQusAo/PahpvlKHrPRjQPymA
8QqmnOCcdrks0TUGayJzvLAA0vEOJYR5LM5ENmEB03qFWkZft7Xy4JNM95D6sjBEte/NmBgP1arL
xR95RM+YG7bdvCcDs3wYfzcY8qMorW2WYEQo76xAk2w/yPmPc8s0evATJsIPEsEd1/EqWmZgYjBd
bDgMrbt4RcUGodeIPRwJNSYhFwfEqehp/o2UhPHhVI+zY/2L71n5KZecaKLaedTUg+a4/8H7nmg2
LWU3bY2zDuQCFntnTpjXjVL3DWBQM1/VjhQ83yXC2IoLNKp8SaCA0Dwtl3LmNGOv6pwTjonLNSTX
PXLJe/HFCkzjVdhP8sHqjqZGUYdwhgRsDtJNIdNs+oJES1eiBwdfGL4taelKmPi7LP0u5yqz4br6
aotCrcKxDz9c1TeCuO/RPKJ0+WZ+cSk3++MZFSfb4Ywem5zY3O7KSYdKwwvyY1RplR4feWvkn1YK
6uAxxRgbQsE87IEvbQYbpE+ZmQK90W0LWlqARdpPnAjIINJKwfs0BSS3eq7A6ICqW8SEmiqY1a08
QnRqG6p5AsjbDc0IDfVhWEEqcIxihGnAaw5savS+I7g3gw/Y8R74GDDqoiPAui6iXTN71dV05a6o
vf83smYiS3M4BkXHDQhYWZjfQQvtfH8AENnmqwPus4Iz5YxBQBCnJ8yXjCpCvPQ/ZkpgM/vJTq/T
roDPPv6F/Ki6HEdu1JdyqUwTZkPEw876Z6XEVg+deAB7Y626FZxO3Zn8J4HOCJctM4Ezh53F8axM
QQllD3UJ3Dzb5rHxwqsFJbJ+EfvPstNln4mZhWfz4TRHIshpMvvw7bz7igY/BPnvB2xqmmnAtZHs
RJs/Bj5rhTRM4MNeSHwiPgb49rYtpyb6HrdGVJsNUKvL7Gsru+A5XzyKksgdAU9Hb44nY8aipX11
8a8v8m1kpR9gI5mvQHxWuBG9StMlDtIl67ikATDxHygiIRSgPUFpOjj4R2QPl4rveZE1wmRQzX7M
jXFUkCkw2RC3UJllHarIcADAwZlfdVOQKmuzLbvTjeF0ag3r514/BW/1DGtVT5lAqBi9RebPrrMb
BdOarjEZK4Rq7NiWwlirbVZR076d7EB7YD0i1NlhYId3Qhb497SUOQw37riVhOfdmE2KoMqSRc1x
TqlnQ7Hube9gqJ2S+VXgpVphxfB4UyB372betK0Ccbjlbf8u/K6WxtvDHWTqH6EXp22VuzmuZYAJ
sU/+TcCEwKFcmCRuy5ph+Ze2bGdJq1+BBRIZtrT9v9RFy3uF9RkYe0T/w7QKy4ouOgmHCyH43gTA
JMrAKVOjDKawoAMKs+mrXzczEH/WAfcsTbbpJQBEFNdwQV+L7GPxw0FlGoQkJCdx8ztsVl5pL0Ie
Ybmzgmdk7QMADLc9+r/Ky8o2kTbf/JTd/PiOBQu53pc17CA3MKK7Z4z5CDWWjizvnRyWz1v2UKCQ
elLwIHD87n6nPwkVe7T6NSgXpD4bXbAONFc4cYtI6J4RGFy+HGzss3z9JEwMyI520hlVk3rCNF4o
3VxiKUMbdyWKQIoS1phfLNS3Ct1e99c32+LCGYIuyr6kHbak/vVIk8ZxpnbDFQhI2Qen5gzeyjsg
fx6UZv1X84lKb1Ja6EdrCGQEtaxwwEBuAhkdhaf+rIiNEf4LtXeZwaQq5WGzgWvHpenM+QSgxINt
87STkhCXVG99C6KnK3UYniNsAc9cN8vw/+OFgarFWYIi8mNBciQGtZCLmmk5jrat981zQk2klsXf
tKGJAlgvcTv2LOwC1rVrmUJLvrP01AcAYnmiBXb5WCm3BAJ5ov54DiuAn2zBj/Ag9vEyN27u3VBf
Rd8yHi4PbFDG3l7fRnxxlRFjjthOhV6LgTaW2bqcPRmGrNJNhLSj96WVCbLmXeu9eP4C7y+0b2cQ
0PbouDj2cSSBnU8z0fXQ+qSvhOP5TxfsEvKGaOn0yrL9B7elR2LFTWdtkorwMeBVpd3RUNEtqc0p
iibD0McocOrPpBLgeACQgvrXclKiqutwEgYKjOg+dnUkWwvaq1Iy4xiWiVPwAMBUfact0aaP2mmJ
/mNbso+WLZX3H6olLtfvWVitxSSQEWt7N2K5t67bTf9OWDBHd+bWShMRezBxc+ILhL1oCSf3sD9U
eISTxopXAHX7UM/kn5BKxTky9LrGeSQar/n2jKmH0NlOUinQozLCneJhAea/U01/L3rA8dpK4zvZ
m5lpsBuxMb8+KRWXEe+Jm962HjH2JVYuiEw6+cfv3LtQci6AR8VnKYmMG1FgxFGqGlVDd6lmo9uj
tPrcs+MQ0umDu65s7nGqefMHloszXloXqZ/aB3lQ8tQRdywl8ftE3QJ68cqI/BKecn3VTfJdFLpj
hQ7FjZOXdca/yFnx2FNhBqsl5gPzbUHDtDfEQWbRvgfYBa0WX0x5ig1pz5YhNaL5Z+jP74jGBkWd
CBhxNJECnrW+qK4kDpKj63eZywkRHinbESgvsG7ClXoZe+9fEIszjkh+Ith7uSrzeGD5a/zeXrz8
aXy5oJsJHd+gTv8rU7M5bdxkOmiOvUAuwzldS+oCNRRVmzyN8UiQUqkydTRW0Au/MUkzIWt49xVx
lCUWxqYY8OQDpew8cFVrq8oBuqHtyRYaOvbnMUrNCcB1aprfyoHZbYBCOZP3LGnmRIPQdLLZFZhz
y4/hup1KjJTWLkH2hJZ5/L7QZWWGdeTQjmTmjq6Yyb82UaA3YC7tReHqvr010IhmkeCRMKlj2fbD
toDuSuQIznxsrDGPhBtWg8iHteWbTsE3dCNKOgUuV2x9jGvaevCj3qQO5aLztSzossv3PjBq2ffJ
QBlUlVIp8OLz9+f5V33zV3YujNrq54zSLsQ4Yvc7VWYHfVYXNOV7nSTqHa+lRAs0G3QfB3m2Uzja
nbhvLDg5QxRS2AyNMBsBSmqRhERhpXd77NdFvXg+PecMZSGfNy3mdshPu59b98rKpmUam/SAmfrr
uzxvH6gku7bNKhOsZBlxP6dERuvjgVkQhvXx7WDPHJOwIu6QA3lDoGUMggf7PKhfYaYKQIiXaWqT
tsUscB7WeBiz2ys+qZpdzBOiVxW150cH2DBH/TqkDMLXPkA1aO4WbKRM44AosSdrKm2gqerrBOhe
uBwDKQZd6YsCDx60KlKFFyxMqpPgqEC3xWPOZ2ykyLQNsmeCppV+NKn6GGCGL7T7dl9VviWU/xf8
rSSn1yyvM03oYmC/cUGkU2U3JIfwhc9e1wFQdNwjfNa5m+haMZrD3x2rd6KDLQw2ZZLIfCit9SBN
B1HMVCXxy6lpYy+k6ZL8Ko9ygVVMld4Ijjes8HsmEvIm0VSMTy0ans7kW6CXpZztOjna7cHPZOCD
+Ckln+FIo1rMAmDXPyLtOi54RqAzRoi7FyZqU/U4pFidldfrlgobs4dtkPQVoDP76ZhOWzYF9il0
p232vy3PN4ajnX3tq6XlBBBSRrTQjgdWPvgAVN+mCTT/S74rW0XxaZdeav8X7NLMFzd+S3BG+nPh
UQCKuVkzxwvaKa1e7dWU4F3TLr2dQVXgv0SNldb34tIAmaa9zu0YjXL/voqzkxMYx7+D2jcwCwHC
gs6lqYRhF27mrmSfJDn8Ka2UCcNkExSOBqgvubYNUWXwDKnJq+jV4grqzzAjEaBGfhKW0HoDrY7J
PaIrNQO+VcqsdMhDC7deiAVADtn3TpAMKrm/+KysKjVjUkUcsTGIetRighvijv+3GAYEPvuKO3He
IDJW0RWxOhgBShcyxXGjP7iDbKyc2q7oPC5qX8D3QvOU40e38p6gDHRf9F0tnyfKsSBw8sF2+rVX
QiznYycCgEbRVByXZkPyWPVVeTGoGfxW04dBO4mPirGq56kgCnkR2WOS7WSxVkVLv4MwF+Lv7yyW
Mw/n82e3MAEGa5csoGmSBh+2Kn8Exm/1nH4buU+NwxW19fLyDZmQS+PeNUAN3+Fl0WYS9rDoE1b0
NexED/jZQfVgWlUgW3UFWmUbVg55QPi6UBxLuNgjbBki2aHSmutkJ3NIkxtPysW0DwJWM0ZKjHlf
ezS9TlJOS+Kc0wR3XUUPVWP5PWDy/+dkS8j4Jbt0Mx5P5a60aRr8ewV+l50un7qRuN7Y+rSBHOI5
UEc/c1k725Bw3KF2COUJE7Cyhg3oToL3BVukr+AGsvkzzPap/tNd29EVY7UE8EIPoG/atbHkXNQy
mjqjtANgb1FiJBevfFU7c8wpZI3s9V7uOUIqf9+wv9gaoe+WPorR8F72DL81h2PMjXbloELgj4YV
lox9407itRFQj2f+4BEOkOBxAJ1JjFJVkifPkPqthTwxt4k6/Si92p6x05bTNHDLhQN5TwVLeIPL
8l9GrQ5FD9bQJbdfK3a5OpuXOOuDns/qM0fbIw6ZtvEZ3FOcGKR8DvvLgJqI+nzO8kqHjEY1bNeM
0Gqz2+lAhsI84HHBI5k7m9CbE4GScTLiEHFNj4REJS2JNuxCuwRr1n40vIUgvyqpU8q5L6rcdyex
E+j30jCkaoc4mkFpeXVP+MHe8RJOrkFmZW3rCekaJQ3f1GmyuYlQ3R4K1EyirID5Su2ov+6soLA7
vOGNHhDO2ADm17MITM0fvFTAAI2yiyp6UVNxR1V3BWGp7dhfTgXi9l7jZcMk5VltZUrgkY4c4BBa
3J97OZ6aubYmv3RI07Hnkbc/CzVkpzs0i2pJJjj67aqlbMeSyIkJYacrhQKiIlp07olPZABF4kKx
WHYr58DKjgTY3FdtGFnWfr6OKu4rU6C//buwquCbgx9jIM//yujWr180R22+dXsAY0iiDEy9KSMA
sxq/Tvp+v3q8F4Wi7Fj+tL3b1+2ievob98wgatI9xy/yH9+NEA7q/nXjTenwseo5VRh12SLUTFqn
EgBF72nFgmW3AobmKPR3XAg9H06nHgXjKExoBO2J0TmrnYfTRw2bhXjI/U/uk2cldbtx+tVirOR7
M3d9HSHZPs4rZst2Nsjq2Cb0dhB2FyMfLbpQ+dmrc73FEtPwAEDLCT4hV3DCiAymtU96Hnbr/QmC
4m+PLtYTvyX1Yw+Wrw+qmamv8JF5kdGLmN/TIAA2Zek2xBzqakDNIYrooVnRU+zHgOHcTlqNTSNx
JJbsVgzz4hjPXEdhFxuPB77VJeAhTbfBPiG5TqlLXLD7armzY0vfV0P1URAeMwB6ETzXLi2LmgWO
Qsz/+ZsYHz9B4jUAYKKd7Bq6YN7Pg0v5SmVqGDppC4bZ/orfyyJ8l/Ip60JpgArZonLHvvaqxno6
hKUKqI53+uFsyhUUV+s4E0t3Wqms1je4drrTn9UO56d/EzNLiurTY42QZcnh+fjnX6T0B3slVg/i
EY61rCqwD3UHB4+eKqQgDSLk7NSq045ed09Wspi53AYBCQ07uusrqw7WepFAHEriHA68NWx4zRjS
kzn/he27iMvn/3fbVpwPUZJj3AAIQRjBac6IdwWTfdR9qVYbLjh2MZPZdBFDxwmYaL1UK6Nmmdu3
brv6GWjd/KqCzB5/MblbHkf7p1kOFzMKSQzPr7wqc+5m52U8+imqnidf+LwARgC4bNEwalhMEX0c
cdOIehlmESdTugX8xXVF2bepA8NK//r/bja0+cI27+6RSRXLTigJ5sbvUF+eBlQsrFa0C02dMFRD
ymNypU2cqREBoNbolPq539wF6mUF6f14sn3EcCZ6r7RsG4b72TnEFYOaBNMl9YMP7RK30ba00En4
U2s8J0j4ESSze82k6oFFQijQeoHcdIAKwCO2HY/0x37lT3k1z0ciA246L4PHds2lrELC5XS/nDd/
fwdlBx2rD+edkmoqkSkIk01iZ3c67Eb2iX/l8RVVvIQ/jtjrA9Y9DsSfUGH18o15iL5DQrj7ycWl
YPAiMTNWwgFHIMWoaYc6890ecpZByFQc3O61REkfSAkfrIpRu5K5yCM1VzHBihGwxiPuFwO/Q/5v
rNzDr9SE2gvzrf8V1F7y2fHEkX2jV0kmFMGSp8fM2EGPYBm+oHpMQL+/vCfwE7keMG62+CullL7U
h1QDwlaNNM5+C0hWsCIndTU9VhebbSwFe2T7GU5cP2p3sUN6rU4A3ZM/xEvXHT0rS7PZP+BkGuS9
7SNPcWMq5T+BlIcp5nWETu92A6U8zhN3G+mLSlx5tCa4NtixBLDopTq6DBMqM9N6w2wlTkhyV9nE
pu+o1+eJMxiF5XHoKxrgdsesxQSDgenDRNmzRIWjbTBeo6gghz+53Vfhu7xOvU0Ft35brdjvGe2a
J+0JbNIvTGEETNGu/QnQmLcpuVJ70fAyF0FoRomlxYp9Kf/xzqmsC5/5a89Gu13uJ+5fEtOev7rB
bwKtpY+wWmrgeoQSpQs/KKePDHeWMhNfMH4chYH4ociVEd1zojAdN/AJ3WAnG8jgDs+esgDXo0QC
HOuMw8fiM4yPvlBb6wqMOLZOao8YU/hIFjI7Cg7hB1qg/lT/Mm/7CuEetjN2P8RSV9boqRJDBAUb
aTUTOGRm8x9YSDf9qu1PT9HBTdD6fAyHtoFIGoNfDhgQ7cXibL9tD+XjoMXbtoEvB2r70VGTztSw
FrIGxT4/2yRvUPJQA11Lffz7Ac07INYYUrAWs3mJw4g8gZKEAipaLRbBh9CzuFR/4VjhI33dGzOc
ZMz1rH0HaFGn5QJ9gGFWSQceJBD/jYTohOI1r9bFyITxFjHyUkcfdlilT9YsamsZYLtugbGjb5+m
87CFxvTBg+wPNJLV32+6ijOBF+N00ucJ/orsvg4hC3xfoHCIWTjildkrfMzVd5xMWUwxAHGiGpmO
b4+NgWQd+VKzy28I/Kl0pNVpyMe2PIRnP5OqRnoOF46W6RK7Ytbr4ILixE3C1cTRVkECKGSDPwWM
8Lj5OH6l99f9nOrSMA4wIjIyyB+t0Ix7aiaEcDR5aIGZWw0zovq8cDFmuVmSjS2hPQeE3brleHkt
gSSl2JxO1pToQ/axjQXnamtut2t3EqI/tcnZdOtmnx2Wxl4oUJd173wOzxDrv4lyaEgKseJRJQ26
NyPUnVj+L3zCkdBnIB61ZvQ+5PJ8Kx+w7CvgGFhf9kq/iOvh2800Vxb4IQPgmVF46cfrk+djumd/
gy3KZa36DDe8cmuBcKoaPa9c3vXzxSmwUZYNFQTkWm5Ey45z44mmrz59nqX6E4utSXZ1GO/sym3z
H2SziOYph+4O9sz8Irl7S4UGZVGQfkY3u7vYZqDt84DGmAAPEfZJTwQ8UDqmRGboAZcGMehITVMo
iX+5LnLg6lIFXeczl/HDaAFCa95n0pnLjbA8fVR6757yKOeZWnQEFBdbstYX1+8wchi1HSltqzFg
jw2PB/9+zzook4fB3ZjPo4dyl4OyDNeU0dwfKwKm9BzUIpWNPJK2qF6/Q+ugZvRAIZQ1sSAKA5Vh
b39ylF06CgFTD+ud/fFgdx7yrCJc65lyvNfqjc5rwCrMh2kGL8bYcL1cQAYeiGmbHvcd3qyNEpWC
hc+24e5JpqLf8eqgwHjRd4+NgwzILFM7d4ic00dJpTe3yFhAXK9QIW8vr1aYU1YqIkOaAUbU3GZl
/fdUDhe/tKOOsAw0x1fpCpVcq6iX0R4JLvmuapoR9OSCdtniaAw4N8885v2quk7MjLOStCuVYE+0
2qvvpQ70D2WmyDBtXwGbgSHCOHM+PxngDGczc7OVhx6v1bEVIBGu7fdSirZkPw0QMhGS9rDMjgGW
61+ewEi/V36xKx6bvAjuz6Ms6QJsMYJ+6Y5P/QsqNMUXnPRMnaiwaZoao7nLUFKIXwANn30ZniGl
sK/M+QpCPaaeQEuMRsXZhD015p81aEnM+eDEDapYVZdWhWL2/0uuuJf+INmYLa+BavXhIEK5tiiW
R2JdUXepTBKwGzF1cYmTRoiba76vV+y+4mLQfn+66BFmilP7juXrcd5ievdBKqod0YFEdFdsAwFR
nGciVUfcuD4smcOhHBTEvZep6q2+Bfw5VJ01aghjE4qOeJsPrrnUNSDrjgOkqTdHsuodKyOrcR52
dCp5rSAHw1Fzxe1CdzI0kZWee3ZPyS2wq5LK6hboxvx754IpVSOZ302OXcMPyo21wiEzc4WCsW+z
+DPe2AK2j1KE31WGr1/E3+vPJbReagWMvOPchTXTrURcdnlRiH9E/ejuqmgwHLM6bgbWMnmfegfN
+jZpKyvYvLglRL59bgjSb01u2bqV9dQM/ujELFEKWYSgjWSWo6J/j/7NDNnd76AWwp0J9qvwXu2Q
5Q578chouEplv4zT/lJ9L75h66xc+vX8UCA0H1Bf+jacf3G/237JcvCC032JeceChE1h8CGA1cSH
C7Rz2mjIg2pcZ2SU8zSqnmjm9OUrp6Rv60Nprl1kq7fDussG3xKf3AbSYbJc0XwG3usOcvvwQe2I
KzlraNgWR9mK7eEQzb1dtZJIwsy9Do66/RqA4cRAG/D+QpyYMDYg206CJ+HYkN4fDTPpdgZBlZ54
sPzHlnkL4j9QMfLgFbHkAKg3iH9JncV6tq6FtPGr118l5dgANpdrS+m4oEF1idmmHAsSXxIEbbuD
Gbp9+r09FczlScpEikZm3zBWIWtrZmO1o8Zh1cfVNL25xIYy0HXuWvOoCgOGU/4aVqvyX5e8+jS2
eHTTFwikwP6bAn12z7eJEQmVG2ylHZT1rLLxPTPLlkdt8WeHnortWPfbB88PyySfIByIPuV/uRHh
U9EumoaMsSkwdrhqz/temhMVj2K3jSlDCQj1+eMtAmNq4QyU4K3pGLNX8pz9J3AndlQRJngSpMqV
LeXW6/3dsHcBXDAlpG1UPQF8cvWTPUad7iHOqd63AlddTX9WL9T1rqLE4cIkM7FsgqpVuD9z0lwt
xiKRL8lrHDseS+BU/63DxNHUUBxooIYV8NH9DyVz36mbV0r2Yr8XhRa29egKGlc3C6h0VGU72M6L
iVukd8lY+EBwy6pnIMw1RsPm0zrEeteKEIeWFQCAv8EaONuWUEna9LhDAkvR3bfFZEMwCQmBJLkJ
9wr0DIwO5KiU/heJHWQuutq9YzJqlKG/vfFNOiPuqC6MPWxWZEnfR/71cHzjZEhif6hCzzK4eL5k
qvTku2lNNRLhK8X1mL70Hg7ixvZ1ZsMbUsgA8mkCcI95oYRC/J2artORWm/sNUNyVel7RAu4yKcF
eNwFk6CEBjCW6AeE8NBKmv1fK/TF+c7R3854C5wGO0PYYoMOHIWTdTZ20Dxzpr3p8hmZy6MiDawQ
cRNIWDoSAOlbGMHv8CQvtjdtMZwE9jbQO00Frq68dIHm8OCH8rbkdnSGCSQq2sa797eJv8l0D+KC
+CIjg0XnTUsWgd28KB/X+XZ0IFCxuqXLGXpAArMsAxPJA4aONkUwS9kqFYE+G8L0O2d3rkd4FB9m
T3XL+y/XOo3VqUoNpgcYcV6JH7x83Wkaxa4DOCuWuyKnLL7OFNoFUIQP296WHfWlo3ju4Jg9qHvd
LALesRB6afXzKOT8chPANGpB309ic0w4TuYFKAFRt6z92qQ5UxFfyu60RU6jfBQb3cuRolir9K3g
mUQtL6VrRfEFypD+L0/3wWdyOD+GToMbC8I2V40zWQeK6ZEqbr1cjeQbD5jq83t8qNPqQZVUbZ4v
IRbnj9CfxQ1o6t8sJjtQwTpYL/rCRtfJjyCqefEEW+FUeHYM5XBJmry7x3pZEg9WMIsLHEF2j98D
JF+j7N4UE2jQdwn1U0uqBQFtuUoI3QliMkBu/NoXjfQNBFlWC7kkGCgrqSrcF6dnZJUtb7aduymc
8HSRDc4N15b6AWs8yg3suMQ7aaVLpEA3qRbEuRQgttOX9bIneMmqmEChmBWYQWq2H3kKGvivBEz7
oKq3aTCvPj0VfkvxOqLR5CUeayPUlpMreQfkEKQ7GsrIm74009veTYYrKEdckdFDnAjJcvdkoSyR
o0QoClB/rO3YGguU6zUm2fBA3klbIy2bYkBOryZr11koaVRng2z0i/780X3jYS7i8/5fURhmmk9n
SwrP0opEzjhvBN8B9LyrlhLx3qCK5UBnLPgAuSpstSqrjJ2eIZTpt0qAklDRyglAbiniO7SXwJ9p
3hqm+4upx+5U9h0zQ1Rk1i8CdFuAi5d9QGRHBEyfkNgue3J8WEmUw6067wj1sMUNNLRYjc0gQuBc
xEz37F0LclCagL5xKxm2/+bYebfSE8P8iZTvvPAy63cFRMdiLURqAui2RiNnwoJAdZf0kjvi3HSv
v6ZuXQBk+m/Txaz1496Ir5v7M31G1DIaA1qXE02UlkQ/zptRCuR6/G9TgN5FAsgVmCTsXFOk7r5r
PS2c3sEioZaQb4Kq4iiyF7yUpICHMeThyOCVLhajdKLh+7kXkIqAVu64rR0dLRb+Gcg1r/sB6pTP
lv0nY+1nDXDsFBYw6ibmrZ2SaC9vJm4rAIIrQgHIhyx3RKRoeNRCRA97HLoSLHjGY3WMPf30rE5a
607MJPrBrY8LS0pBGJ/tNEkCPJiGJfwavWIHnGi2koRRjdnyWrh/WmTWuTV/No5lKwUUo6WOZP3a
88HyPqLvYoi1kSWh20l5A/+y41xCtrLYWKiN4fAdipnvtBOJT7sP+ZnoiDprPPmNiHX6Ub/paMmm
SpYpFfAjWZ0AkLsyCYJUzPDL6GqzW/sjKOZvRbjsv4jy868JpdxBV+IwYOvuWjuY4RDl0q1pcgU6
jCZ+kMiEJLfDdHAneKCgesQop6pg7hb+smjrWjYVVFmowUfq+QRGkIyqkRc/rvYAMIdnWYlKg7PI
4ow6ZF7/i72AMDDHan6rsPIcvnWPJMUIqFZ4kZfjID7OJF36lqTYldj0PzXCYs/rDGHyvMiJXtqv
z9DGkkf/Fo44khwHwW4/sQS+Zif5qup5HSGsRLKtlQaRYwW3VtawrhagS7AFXJrdkrw2Ori5vJVY
7o+xrl2fv4GSx6rNvX+OsNucr1lVA2gYol/zbVrFf74PiDSQxEskZ1xoS8IROo7MOF9+kJksEf84
WT0kjHjTjIRsWSF+88ZvbOL3HPgpnBb3nSRI/FD4S3dqwQn5jgbJFGL8iVt2/LQTqY5hVgZvcLNz
YmzJSCiqBOt2PZapU7t3kQ3/ksfezbyMHqVJSrK2Sssk1CpuTuAbnQMBEEmgsqHU3hlOKAwU9dLZ
VnNxOc7otVfOhSFifNOiaWlyqDuaFmi67pZfH+uKqKmUrxAGz8LcH6nbfsS1ecIYHHRlQZqgPyFN
khKNTCaA9dXxq672ZWSF3U36NJfjp7Sddilx2y4496KxRpKQRFZYnangDzsiL//3G3MkW4y8ocau
qflg8sc9gE5vPzdAYNtb4F0bG1h21wlNBdm11Lokg/iSk910A55Fcz2q9iDhAXYrVxRquz5sCAKf
WJHuaTxU67S7dTAo0RJfbAyzivzrsfF5dthoeXRSIk3eOBiTcrEdp+izY60hsCeYrEJur/22nh4l
5sm0Ando/BlnX7aUemSb981KeS5BbsIh4udE68UnQ8aVCvRlpFRidmtPewCJtOzcHHXu1CooM/Mx
8dTLrtyBttRj6BkMPxvjOwmFq7yfXVUxZWixRmdlj0t/kcupkQK9v26xFxF2YedtstEKA+93WaAt
PCoaBb3jsimxzCXKSC65mOh6mYB6LH884eac0NbuFA4PXqAzWl6VjidRmjsS0d2tEk43Dewl1zaY
nt8rJhx9QPexJn8oiiC7Z4buMY+wurNT223o3wVTNwVTA5YryqZ3whkyiv3r6T3kRKT+xgNUwf7X
3qd/yQF6JpuKx13mmD1NIuLLgTSH7dbRn2stOiiCX84qibqCIiR6wIj8jNN3auUJepjMZO418BU5
4ErtrUqv4PyAOysbSb98mckcXHUM2IwcBQmKtAAmCDQ1iIDa06BhN2VE1IxcNd+gMfHch9WBMnpL
bLEm8PEbMYX635CUOpRey4xUzhvqj6ZMnwM89Z5xI/aUkKYIJh1AFp+QEjxcIe4iz6XfdYAIeU70
NBOHCpvD0iZ/gkyRo6LRHFr9YfgYe+Y0kXEuAMOR9enZU6DFUSDJVWEgRRk4py7C8JiaMzcw2Lpb
oMIcBdiraDQyju5q7QYr8c5UY6HcK7CSNLprE5Kgo48QVgC3Uz+MI6ytu1Lq4/KrZ7v14w7GGwl+
/ZGm0TcZFcM/dVLeSXar0UV96crDXiDFwLvWShBDaC5Qg36WKHdshVXQw9mqQOkY36jJ6SRH8Uu8
ztjxc/whButXcamNCyPQq74GdlN1Ms7Xu5YgkwcW3sV/87nXl3FDcMeB/jHhytG1ipnlNU4eEhJB
1VNLZSDJDNLZdCXS5E77UTa+4qQVCGUUOhvbO0edJdiL7qjCDTKnBMl+FvKwRCWcVJN6OJy4Jj4Z
adC479cvhlkShaLago8j6MfRAHf1jLgXn3MOse2wxI+kGIa1hz7Ttt/X3KCrqQ2awNhl6FhFbpb+
YivWFo1Vhyx1uBUL5sQ9Q5ZLl7zbW4jsl+lTB85Yx0w1xKSDl8XTAlFx/a0Qgs/oGem6+RyXZOGV
lX1Yd6ujNFypPtNgGCOQEX+D5J1k/TWmZqNf7awMzxCdqIiRbLQ5LmvWccTGlg6v/BGov0zW2ild
BtmRRY3mzNz10jDXGKo94+rzujVILZX730NXzaBXDmhRcTwYslubgyCuDMVfmv4TcyysuImO6cEk
nIcIf8SFxabK49ammTzze8TqWZRMyuTvGgJMMFR7WhoxwL+G8F839nA1utVN8M1N0YomnB6nmtbc
PwS2P07NpATamIcJ2nbXuJQkCh13o8YbuheiWB2SKyxeOeDy5sPHQU6LaFwGz8Uxr0uA0hvKMI/k
KoZXd/CWNuwze4ZtIhu8VxyX3oDT+X1yPo+GsQgCAJn5k+xn+BTQxzR4U+WAvnC2SfHFjhNdwjqU
P0GTj7i0VY5u8hbuHmIql6ihHBzB9MIQU/JMwPh3Jse0AsH0wQKwvEg6l0HnrwnRKtHUarLdTkeR
4Uhu5qRk1baZn6UDb3QiDUTQag4lc+P2aGm7zDwmcfrFd8H1oA/Y1uGc7bpQ3oHlMWo4IoYfHirh
f2IklfY/3cDKVnnuw0VFKlxMsn8NBBlo1RJNphgaB4dyvCNcdKSua3C11K1IwWgNsTBgh40Qi5nO
2ds7XLd4rjWJv9jx3tL2iSWZscK1TbY8W+ccANreQdQFvaLeAw65VJNjFIHEvI8AvbqmpjsX+w2d
yHq+yfSAsGigAyXho7Yf+1wO3ueT85TkHWRTGZ/WHg7fiYWDYcOhx4osp0M6i7v765BziwvgGr5M
AJSRnzCKZPlwtVPTCRK7KgdHFWwjYdDy6c6+k2zjWKLVZIUxWtcEnwsbRJ8Ui8x2pOsg8TXvIj6Z
aUlMcajqlCLJI5UwWO9BLoBxkGVbaU6TC9S2csrdVoW4o2uKEFXl9LgSFR2RDrNpTo0WJABWIxOB
xmHDfcxk+L9h4Z7NVj/mXpkbDP8R9y+W3comzladzRLX+gzxzM0Tk25vcmy/L/9O81byNOdg5ZK9
QfRHr2Aov5vsAqwb2sRoIPj5kdJ6r0FGqu4ZeHnibriQPeMIi43Jfa86W0b7qG0kHbJScZ3O7eYT
CbON4zSF/yvBp1o4Xk3sTuD28YKwwpV8rOKJG5uKFac9GnWCxuO4Kl5LYPem9v/w2eNJqXHecVkv
OaPyLkUJVUyAiKvMp3Pv16aZyEc/ArYJ0yCQbpLuk7l8zqbHKC6v2Fxe5Od5mZ5OSd/bCXBRpVJv
e22b3QpEdYIieoESpHRNs032WkEvxQ0BQewE5FIEEUuzI04SjD6uelGevM5uj0jemOtKwjJQd/sm
kIdgrQjNs3whhy0kKS2bujVkH9wvB/K15WnXgGdXOiIg05+ienL0giOU/jyUv0xEpZVqP6Xx8j+h
/B69Wb7972ESz6MiAnzo7pTNK8S9TZhWIGyBtn/pYJya4BmyJg96CeDb77rZord0PHuYV4bwCB9K
D7XVPdAFsaBtew/2noARECBGY2bxBEICsgQX7lSyfqcE4CTFnwKt0tTOcJFwczMvOvg5wiNMy6Il
1Jwy0hBGrL0JvHQZBXDK6vdygVzh5BI3A459OTKRyRuVj+3crXcGZb3MORTuXN0hREMF03SaMKcV
q0hbfKqrPZIEFMmFa6nmDdp9FjMAbGq0JoKdtCseaiWOrNP8IkN2H1g3Mb2kPG6qn+0EY+E/aHK+
JBJXBcUn3xbuTlb6NLhHPJ8Fm8t/gtjpmfz7TZQobBv15qi1tBeT1+9plE47+JvPbX2i8adre6cU
u8YWdvec2HnCS/N1uiGt2bMd84Y4y9wt8GIhV0KrcMh1Zz8a19NFQUzEBhPQgJrN4IdTJMtUr5Iq
0iyD5WEUjHtGsQizifjvljtsseohrwlvmuSFl7yeT/V4M1D1Zn+Xh3UC8tm4RExxuePybsmMST5B
NiAvgEso6xXoAj5iXUMJAqopVhNNXk1s4Wjji/bxhmM4urOU9TKmMhPLNhY7aUqpf1MdrUWmfVTj
qVztUQEMUh23MYSeC5gMbNLOptjBJ1K2hoGG+FSOx+Z+ctuzZ0m6mjKAVTqSuQswqdXvbanRfYjB
SZveVtjontaF2bo5pnHePUCcAkv6KK+NZRjDxa5hQ2Sucqb/3HY2WUGwlbrsRVxDeA8R8BMnvqm5
sGyQH/Db7bHDKtcfeQTyu/vj/+h0wTxL6UuVpZKqcva0CtX7IQY80K9gFZY+UFoEan299Nz6EqrL
lj4eVFUonDNON9J0E/N1snBF1zu6Qrcx8bRuZNAGPEcmrHatHedeGV57wXdpAVrqGwLdJ2wMn4QH
Xni9ecfrkBVamQWu1G46BFp/Q7k1OsFW0tD9K1CyQefjMgD2t4acJ84xUGUVDSjrX0TZ8za0fvay
jhCnpKiINxSqho8Twj2rMIIm9Qf09rWecbqImEwIYfvm1ZzuqOYDd6KOEyIxZvMgo3rSqcE3ZTCV
VFdt5FTEc5jEwoINRB/P0FmOz30SWNc/Ps0DD9Jt2b0dpUEnIRAHDwEbP2geV0spxYJ+l24smzpT
32HfH3fp111sXIknXz7/AV4XJZdWRJBoWETQlUM2nQp6B0/HdGTdBW/Lr4RoQSEPfeP8Rq80df/d
Y9lw3TssunuGHbiCHY8aRQIGS9yDqjXD1liYv/g6Wp8cqlcnjROXSJ51Si0XFEnWZSxW9DLxTGe7
Pi63YfcPZRRtWj0QFIGcOvfeKycrbsFkpqEYfmmzGc9sSYnQ+VM/+QC5+ttw9XxQn4ZZR7yoC+nx
JI4umhXWerXLLXG2hkWCXskRtJ8CQhpRZGe5SbNQX0lpjP6pmCFUyQuRhTJOidcj+bwn7RE/4JPh
P1QRhw5+yTbHxg1QV6XmHF/Icg3Hlj9BsvuLaw9vpaT6jAeq5MDXlkWk0uUiSKTaKNTYODBw6iUr
cnp7Gk2pcry8Vz7z08Rm57aXLDCmcJ+yUu57/jCX2v6cH4R30km2uhfIUeBq8K34BmWDvNflMDMo
GHT5ryMrQ7TM3RIzuKEYEUDZrdQyPRH8rDsGu9TNha/OKHjgF20RZ1T+JEm/DlpFXuuXuRfAb06E
GfM1Ke6Ee0Wl10CQzCmA4xczJ3ZJTGpHI7aTM2SzQ08w0k7G5EHJ1SwOkjF93U0K0a/9l+GkLg02
bJf7Ooj6o1i0YTK8KaIwnbE/Qs9TrOgTA4w9fm+i6Q/iIf3LHpjdXUa5wON43Rt7uN7i8bakm7Qk
oFz6PXCy1PtSofIpkoPAaVCd5853s9CVkCRiBuRa19ilvviwdXHDw5m4sD5WHB2o1rIvnMVwGQXH
/aZ3Iuq//vHtQ4Dke/XBEJfex/vY+qZN8EFDpg7msNCko+7Salt+3vEVMkUr5W7+6GeJoZIc4eaD
PeXjVAfTFS32lV5hWKtEHDXgC4Pgl78/hYOrbJGQJoQKe0qDMJnw4C6DEu6+uDeyXlUQ3oX/tVvl
bZuLfL1vMRSa21+UZqSiBS6R4wWfmaXiuPE+KEcMmJabUJNgqny6hytFbfARVp7oYqdhShL9WeTb
3mOPEeVjGKExGVBMCfEomKTXLYmQDQu1VA+RWd9mUXCfNzm253bYE4THZMKhzm9bmk72atM7shkU
6ECF3s1ujVgePnmPkys/SPqiwwjEBLaT8HQ/FTHm9djSuWvoOV8pIQPaLdmQYColR1gFpTFEAX5w
YsZaAsKJ5nM37RLmB3QK1i/rdllHptJRBQvn3OfqLrPfL/0Ax+V6utnof5OF4HSKOVAKqV0wXmnq
xFtPrqt5NqBPP8cZIPWxUB3O3RiXnUj6nk3gNOkadfwcxTeyNQnA38UaMXlLhb+v66d0dajfe49u
uN/UrZJw322QJHqBIhbiLHWT3c0MUtUPI+3+QM+dDXEOMt/ACUZqguHIXa+xmXz/iWjze6dMmHZJ
sTvEXIh+vVlhRbMvs9aOCoTSZ+jSR1NK/EG1u4SSNWkA9UD+02UPdWnrNnSEfZ9/udN/7Aj3k5Gt
LKPBbBUNWl4n2Irsfz9piO5OaX9stA9URhCZlEB8vqXGTFjntbCBZ4xjdrfDzoOwVEtPkxuItlJ3
0yvbRYAbPhAEXd9B+JfTYomOxzFwAwWGx/5vLNb0sOchHXL3cwPJecz7WMIURZCVDH4Q6FGzf7Ll
PaS1kqCJUO8bS/F7ahosZXN0JCjH552NGW7JHdng/KxnyfiZ82hChTQ+8jJX+GUbaeKG6RO0bqLi
T/H0W+EqK8emmLQgcp+XlzDCtPmYN0xR0Hk4G1l0dmr7oAdvgAYduZiQGZDWcG/p2eaJ7xnLeGji
3y3NFSmHb3ojjlsz/YYFDm0W0G2yoeWj8+4bIgsyX6PvtMuPheMqBKluOf1yRiEXLCGTEKBvxvBW
qXMAhNZIEgaztN06KuIU1QP5M2m/R98v/dbkmC74xNE7nFvKssRRmKzt9ejrsjywva5FV+cXGpIs
ywwOJnbhxGhEzAxq52sZ7qwfUjCp3i2R7UiwYzExGhmW3uwYCQYtse0PXeXn9oo5SHDKW4Cxmuwk
CWoG159unkvUCdcS0YpYkNExntXzeLsCS3M7QVHkyA8N3BhiKEN1oQ8OzOEOddCAzGRfafSKpSJ5
tHxMJ+doTHkBcJSwNHPv3UnxveuSuxGP+IefB8uBMOmb2jABgAHGhyDZhaq1XcmRC+EjEyIjWvS4
XzAjOTpOJidQCmBdQrU5HHWBR/JUqwA1LflD4K4w8LmuxUpsm9LRoVihj5/IQ2OqrFaH8UZTiTVB
LfV2Hbz+2L8hT/+G6ZDfaO0dFloIMBWJVadiukjOLjZVWat7zl+K3hWMTgu55qK9isUyBgK11nlK
l+sZ/dqaxssKRoXUQXCmDdp4vAc+7r9s82J7qDsWCkmF/VdGv7/E6mN/T3en7vqYH6+gIBwge83t
f30mN0HLX4V9xH5KwVS9CniJe2SFeTSxOBNgyXrGqH6n4x++N4BiD/UA2Xik43DKxvMtschtrswB
6ibe6DuJ1h+u5H6UM25rm4Lj4BItyqFDtXbRPjENElu8W1WLy2WikFfDsD1rbRUlxSZqg1NfQFp8
3ot/hYZfHj8QF+j4XBIyYWKDEL/wfL04cKClz8NAaYZBsFTXtGdbyYJ96WO1gaNFqn3olhqeNYrm
pPkPCMmZ2dAOQ6aSqDoxBZdvn5uE3tsDZRS/3P3RhDZpoT/2EuD/i45Ex4Bf++lxPN6IbGA0Qjwu
FWw3XcwcIHGUffhqLab5r8P2FS2zcyRMRa9Dg98PeW9LF+fDAEKd8dR8vp1pKxpLo2FZUua104vu
ZybTzwxb/i9iuP9Bn0hepJXXbz6TobsUj8QC4iu11tNpxnEqiompODagzxnWW2CXazokAv+ipYZ6
M1RGayP5zK68f265BvdMCeiz3gaIjVFMKDJgj2m5bnv4/dgN8X7RfjfmEpDVZ0kVAxJ6Xg4ocoAm
1wVYqJQVgVTFskKajaFb+4dnn6ff9d8wWaY1aUQq4Mx/Ei5mjcxzEVnSdGdemUCMwlUBQCUKqEJB
XfqC3YOSVe54n0jNzaSCjKnHVeOLeEMNoD9RPTTTHgfKMVzi2tzC6nibQ2uekxFg18RZAZ572rsI
pDzQgdqoOBJX8zxhFDqRXcKarWVJ6RpDGLcRGBstu5FcALF5ppeS3qftBJCy7jmDUCW7tp8GaRCH
T7dHScNa4anqOZUNTDB5l7Ffi3Jtnp64/gAjF8QOIvnR9PbuGzc6P1ENKuYsJQr714O7jXqBmv/w
S/xONVhm/iyOCSqv7mMKmnLg91Rr1JLxa+/SzHOskEy26mdQyRN+Go6tzz8/+eiJ2XbAZv72zb4m
nxinS+y/DxGFw91jFPzOD0po5l0B+qyrl86HfXJ0prqRSYw+hY9JzB/iekGOhhrhA3l6UMwHj5gy
DH9m++WOLR+V5EDDK0XYdvBeKBYY5XWjt0hT6CPDIl2cEWzXBQWW5yFsNB5Cho7AiMWiBkPWbHZa
vlhzSAcbfrZHWmvL+LJ2/rwYtrDZMxOKsI1k+TEv3VxegNBMXpt3cLyedILAJsxxt595tTVbjKua
r1dNV6A95NcEaNJL0zFj2n703ticbnne7WzfXuA0iyQCy33oPQY4YEOvhvwwBOOcJwG8kI7zGHf7
8MzIt8mDGPYe8j7vcQevCTiC1QQ2w7F+5BTjuD3EctOzwY/uxt00vNBGoSqT7cDsdvywADL7/5re
CAUJXVzdBWmfAfEhOPcf+cvfkqbGOuATMqc2MUDWLDQgEP0FbwnnZlPivfhTXy7eISwGdw/wltma
kxjTjjRryK3YpapmwRBZdj8laj9nDFC2Gl6KmbJU5qth8RoAAA4YOrEAuyuRm3BvPJrxmDG71Qro
V2LciK9blB5rmwJI7TuDpWi7iAP99+FwYc6v/VN4vsAEx1YDBJI9qzfNdNtZTKgFeFR6nNRKdf/c
HhGL6SfuRJ8s8UPj2gz5Fks1k8Zecoihc0qiJS03xdF315c0lP61KZEdQuOAXpKEXe85MKrAmXPY
n7w+NfzI2LhHGHGPFBP2nzbUYzkkwATYhCL4NVkDUwSqVxNVkA5S1Bdd72FlU2X5TtamR5wu5eWy
q9ehs5ox/C+hIvRjIEM15Qd6S3v9taYtPDrqdPMARryid4LS9b7kVkRNaOIbE8gbjYsmWrjIa9Zs
D0dXT47T8lBnCNSmAxVc9uYSyEFz509317WW7lMWrLt9VrewGBtgct+j3brv2H0X/e2BR7tG4iCS
yBN009n322N5149zCc/qE/xz7FxUE6QL6SwTHRLQ+SORSjTVdOhjQ1FVk8nZMaV1spX0rX1hSMCx
rGN3FUhCMbynmMiW18zEGu2EEwoZyuj+mbYn4J4iDg5wXqtBzbRw6rN92KIqBf+E9Ln8toAxiY4K
fcIRaLomUBJGtayqEyE7es77beIwAKNhz7YgVQnEff445TyFOvvdA8ugs7BvQlM6D5wGnYDOmChk
O7sTqJ96hJhTAqqNCIhZItSbRbqNp792d+3x7KTNFp+UAyPSPuGwDA+RabHrwWdRbqpRB5pm/2GE
EnlcisZqa1KTXOb7LdjTBsPsxjJTpcPWauAQnqJXECxNl0o+o3UZPCk28xJ8gKjaZi+2jhChfjQK
SdVSSoGpLyUBUMrghi2xnZv6THYr3Ldi/u6qFNhnXLt0TrIwZFpL/ubMp3D6PNOlXzGwEm5j27bv
zVBftPvx/EK7OnYHQ6Qaq335oFaJGfrtijbkAm5/5cWt1IZeHYoLUP2to7sNaHQgctq3yf2XdTY2
NHXOZmBGmay/4QUcjUTT3a5NOvbwNFXhOsgCKcf9uewhpDdicnTV91cW3qu4Hd8US34L/V7PRIMf
6UCxqs+TWUjOUqBYjGpH0wUEOPNHSawjX7H9PY5IvohhdQk7WGMkFbYfNm4O1alePZjN04766dlU
03tXFys795f/BNlXEkO76PTapnF3cRlavc0gkV20vjYYYQNIUenEofQSSZoHzeKbdIY8OX16MKeh
rgMRRvZV4T74zSLgvDuxlW7hcDyzz4DFeKw6uDWwELDC/TVJOXNlwD+Zgptz0Lszf4eI6EsYVXbV
OFsyKqxkR4mLTBVCx2N16wIMBpEnqytyKEEKDcd6LayNTd/kRYGE90boBBZFE5divcALOA+eHmM/
z/aYDU9+87071sy5gL0f1MPnmiTvtrhPG9zFBkGxxJAjwMi9nnfBoTt+UGd8Fx9TXNDSLgBhWUJ5
38I/mq+shT1YafGjkN0L/FcMn+kCelyTbN9Eu+2cAAPeIYlgJLrYQeO5389iuKSTqnGhvBq/WjuF
0EWxaPdpsuXCffqkgjHWvMNE5M8OjyenUxwrvfkTMUtME9x3c8sUASZNZTKP5SKqhVGFm+ekyBlT
Ia7YsCfSDpVb7cF7aMcUxGj9xKLf9EHylsoKfvxZAxNxG90ObvZXr6RV45IQwEyC6+X79gNiZ800
4WhSPG69A3elGj3sWXKalKWdf7Gk2PuIRCdUYZjJFpQIWgu2gCQ9SyRLaRXu4qQ/iNCQ5KV5+Zhm
CeCHhxA4LccDEHEsbEnLYlprWaHpP53XAXtmGojWgxc2eHyZ6l9tXyvaZs5Q8j9GSDRFTVa1fLCr
6LNmbXd9L80VEwZnk1Joq5+a1K0k7BO4dwmBrgEV+I8Z3Jl0205DxuAlsbfifVn/ONJurODXr+Ym
MuTerrauQPo0e91iCQaNsorVAIg3OTo9rUxSRBB5N0LXVu33gxiE2RtJHHMFVKVUEeQMpGd9bzo3
92Hbf3ZHGN8iqE6P5f2NeGWFqjiX8ZZsgbFcwKXsO5VwVSJOW6Nnf9b4L+bnGstfJ3haq7IPjNPP
9Qs3dYSSf7cpuXJlhdgU7aBGQOhFt8o5tY/J5AUo2McHdyiMEQQWMx9YR+zz/MS44N8uAJ9ZRYdb
DTD5mnwOmkBUaQsh9mTtxWOUsQX2NjV9Ia4cKVLyet6XWCx4+gfVP2zVn43eysmAJjvZ9v9ZZ4zu
C9qzrYxFDlgyCTxaVXC50z1pxtpaZanO68fyE+1sYsGtbgTCcS4thakMvbzxDlDf5TDdzQRZKNdj
1Qp/Y3AewYS+rtUoQxHRbpBr1mMbwKa1+58iIKiNrNPyufQztF8Wfn8LDp+dRL9hPVCJtuCGLi34
hukz5lGccRFvjQ8BJ97nD/GXEqaAbOC1djWKeI4gDlIuSwbT75rZmD2BW8KdPAaZgbxPbQzhLzPC
xZae+EU8zUWLgChXMrJ5L74LHQyEBIqcu7R2RVHnm0I/qkMec3EUBQRMGDuu6S0KXGUWqnf2QhPy
KEzAzkub+hrpzheLInLSA3k6eOu3vRunpgfj3DCp79y+mbMv/E2s/fa8ELO/E1m5eBURAatIh32d
yjIhYcKds+OimDOIA5MOvRZlZL0Ty89DfmqAR+7OHIfm6ZS4CAtOQQXlzOkquDB7u10Pd9mTrEi4
uFACx1pB5Cox8e4MNOuBWLmvWUoXLTPBud+W2IXWqPEYV5JguqjwY90e56AruX8LxvY2DZckGXrR
rpvmPz+OawfCPs5/5YkYE/Grmg0sqtlzNIHuCT6ZU7peUute3tDqoHt5+fHlAUIZ2GKuPAShpyc7
+5TZbtc4mlZ86LrAUcNZPlnu8q2UEfw4d5GzVphuCuFVDpm15PtNWKFxDKlXiDUqWNPMuLFrED0u
Fpjdz7DUlpdzM0HuD+7Md+14E7yl3va/Zr280qMJorxFvLg0/EprMn0sesqqbdwc7MxXdyFlgKAV
2+mZsNP7M3uWm22ruS4dT2KfjXRUt1fWcbQMAHSYycBTYBz97i+cvSOgfn9T9jMajdnV4+2ZSo8W
E4gO8QYkvJwRggT0jNj8JVsBhJ+VbbFyDQyGqu+a8d0EH9pDDn6N1nSGeabumPvJMGFIQzw5i/sR
KgDxspF/We9dcIZEaruoczGIfDzZ19JBAjsCSwpVAA6fxZK9Vigds1FLcPF5GzZhag2P3PL2hgLW
lWlF1mUswWjJiGW3i6JJMZ2P4YFk+02f+apZ0a/zK8DQIyZWYKIBNCnp76PMA08Veofhxxbml0xR
iVXAyWQyz3McLQK7gxk2YS94+/j0KyI3NtHWIVQ+fg69lYG6ifwnQJEcI290+wumSTzvTqN9gTCS
dntaTUqjHTuVyNk/kyWCVulakWBJaacJuHEPkTRUBSNjwFIlzlylqicXg9icS8anAYpIlACdVY4v
ZvlxX+5Si+hGpjJMjGJN/yMh5ICHqAS/wkbnUKeNT/Ywb1cd7veMvk8RH0IozirIynTb+twD+XZS
7h0uh/Wyw0Fp1XCf1RRNxX2gk7wZpOqa83/tbsnHvMaffUfp+L5UimDjEfld7OwYfSIC+U3K8SNC
Pdr1aPXm7F5stYtbqRj2Rk6IkjPLi0S+LYhaZMzuWxsJQkPGteks4GQHCX6a6vRaGAMxlD4Tbw7v
8M7r5yXoINwpInE8zfjkTZwBW/9vK3Jk823nCBH9Tv5l6FE5aOvYRt4DZSS1/cteLJAvoV2AmnGJ
4PA55b1tF3EUb9EuYwFsxP4Ls29lpEGP+zcGPqBnI/0wZCA3+vUjqbRGLEyBfwcamOMxtod2TlRN
nHiiTuyvrYnQRdr2woBgI3xTm01Gl3gOoAR68TgOpILQ83hFG+UU59mp6fPv4ZjQ8vnWCQENRr3H
UHkJa6wjivjl7TOdJZPFKTF4o+QW3NWnIBXlbR+KsqE+UNNv28iWicMD+khhLqwTldp0ytkTO8Xe
O08FipBkTRNBEeXFtsbvr1QXzxTcMlmoik3C3Ooxw/NvCQmMtWKRyvFXdLkfz0bqPqoR3IM6Gg+l
4E0m3YAvkZ/NY8sY7w/JSl3XKJ81Kr5GbtzCF8UIkK7II0dODyAi71A4MDF4kvtj4Up1C4iVMDC8
9O0m+cSwcGCj33yr2XvuNfNx9TqhAvIuifXONtdYPbEgRzXnYdXSGO5Vg6Ycl86lMpq3HOCq6SRJ
b0yEDjQlzPJi7EIsx3hBlVaO+dyVWVD4F2EptE+Ljdc9YZEgbPH/if5Nwm+CeHnVL/bPthrPyCIA
mtvQv82qRQvzthax1RpUI8EW+Nk5ZCjbatbKVjy6AukFX5ctL8xzn9hTVyj7NGbdJE8voHXBp41M
D1Nqh0DlWSTe8PPyMNmiobPL8S3pB43U6w6QHFm8aBSiAUnX+7i4mXwSaa5U5zv5RuFExw75PdO7
qofQJ74hGynYkG0xnooCR1Hr2GJHcDz8S1vb/bqQ1uXmrOpExoET2k2tfQubkMkCAnnxGSidU1iR
4I4vssYucCUqAdJwpgYv/g/EvgcDFZe/icyJBpEkawC2yh75UdavEsWinM1BX//Z1hMHo5m/nMUq
9SQiGVJbIP2z4EK2X8rzdx/uBGk2TEQFxhEIDY+hrIaU/OfCgGgBmsUAmNCLWG7P1kxeCYnlp7WA
9zVyJ9atPmfMJuZMxLQn9dua1aM1x23fbk8j6nQ4ePPmTxCQ9J08nznKW2rd0i5Wp2GfSCcPR4MD
+oT9KYDcxCffFsY9gqcuZBjAGj0f9RGpPih65kJvM81Hf5XwrRd1c2SJKDK2OiGLshUFRoa4NbQp
rYNXxufJVHkR/WjBJuSEZSlKYtkIhvvbpt1fenSAWi/xQ7fOXzB0UeRgIbWgiOQq8venkCyVx3io
jsUGSLc/Y+lfoCjT0K4rLBuSbuM6x70cjKh65f0hQtTbHodiAK/OMTPpaxQJYpQQDgj4f8H37tXk
Vptqjfm8f8j6ulFNzTFcuWXZ/Ec5bnj2xvqCq32hi9U8M8eTeOaMnv3DBCuc9gMgbfVslKSP3yyI
6Pwp9o8WTcItQqTORDIDu1Kngr3eOhE0+UsK/LSg84pQ3X9nJeKbnPEfxGs8onBsDa3U5ktetgLV
nqKmN2IZBWnb3Xkk1r7J3UuWKmrKkOT+VvhPqdNAebRPPJr1kfdLZi+EnMAzfLPB/OqzbtJMn7hm
5h9l2G8Cb7PGGyqIKZO31KETKyow3q2QZ3w/BgKH2/pGyx3F3YtyUCYda55lp/ejITeEyW7ilVW9
NZA+rTnBEXVbWqaWy40kGD5U7F0Gimq2DVxfJlRwZxzgSt9m8U5z22lnevCEb8VLI9jnY/FbbFiz
hGhlb7iHgpKO1TPq9XHp2ibKEzBfL2BErrzs/nOwzDSFAL3X/QmK5TtacjRJoPYm6WSSIhqOOgmA
ixd3XGkEVoAkkDLcgiqEmBeyg06lMR0V83ILw6CJMybuR5OuAsjx4xnOeLdvwwqaJM7ey5g4aDSf
qRZvVYiqUJYeizSjikaMTv47802Izxf9D41yww5BWjyzdMYUcX4gtjJ2KqkcxmdB8wLmVoUtVo2J
8/Opb3JMhzthL0fym2SGbyv8n+lz6gtnjld7giJEgES/ZbIKtkwNNrSincyMjsdqfqVosNpa1oqv
p3lImkrm6ecQ5mFFYluTOj1Y/WXvmUIHbp8leTjBhaLMKHvrDS6J1TosWWMPAzM4xI9lZuUgNZ1T
jTbIGDT+POsrl8lhRd+i+YNiPJ1q3f5P2rb8aNEbG4PdDFOKVOQ09/2c+smCsV4X5ud/H9J6FAjj
lULIiFZDqjYEpaWeKf00oRn/fEh6cKYfzFnljuewjAk+DbtrdHcd+hhce2Wwdx97Lws4dklQNyxm
3/u1A5JHJhQeIz4sQg5efX557osOdwIYzyNAWNJAUrm8o1/nn7TNlyV/2byyHELojdcnFzVQyqOL
zw/afy8jCgIj7fM+sCVs7KMYZk6zhllpZmZuQzLfSCMjkeBA2xCHPQrg+fpNZuzUTe9NIbBirCpr
dysNhzwkai2MAni4hrjd6+YV3DzoCuZktTxV6o4liCT6o1YgGCcoSEfz1xJSOAiGoalpwoSe+gSc
MkfhKaWecU3mJS7f1Zo7dIh+dEWvXnxk/mkEdYFMHVpZqx1GHjxkiOlLtTgIgVdR761oflrxOSR9
vDbXcUaq7eBnQOuGPeB0VCl7uMuZ2qea7CploWlXgLhejRTh3AlsQZW11x5QRbQ5slo+hnQ/xs4e
ECKJtS3lIvOOLS6DngSEzRFbvNtCa5jAQoV7Wxl4mPLAR44mdBs9XMt1Jdu6cSJ8ufOaGgnhi+hU
DLtig2nKbaVNDIFilJZ/tXylqykJ2BjChcQEdB35SIU42NDy50kiW+XyifaLzPHxF6rXIhUCWkS+
mF4pKqHbIr2yGX5WixWtyLI1yOeTtTLSugTKBTXNfDwVXPztCJeGrhh2OQuMpS0jBEa/xDdBOfRV
tlq7ysDP+OrCWCRsqj1Fo7vMQqifD92zU7lfFAq+bDbN38BIQoLTYbMaZw9C2UsI40G1uT4slfGj
VnhwsXwF6YEvl3S9tmnfU/u03CFWjMVkX6GbZhLW9HkXcKdeclOs/WRMzNndH48+CV3Bmoryym+4
CkzziL42F6amdkSd9kcr+dfab0F0eUj51Xfd3x1pFAZx/SlAfiMGjC4GoMFahLFCqqIvmrZqYw6u
6Rc7C+v41EWBFY995iQXUzUiqoVsjSAsmTbFeatqhkpUxAWYU3dXDZ9lF/XrGuq14n1CxBlqktu6
CFX2uZhnPcDvjG5h6jpQ28kElpXhd+xzbOSTUdfjibVuXC6P+o8znwyDuzArXDQTNNBxYU+7KIV6
1STGt/MceGNTg2sjthqR5HxpI2CXEQaanPwPBUCPAausj256JRa90C8p5/sGahMGSIwjgRyJ2v2X
ygUqZvJ3Drj7bQIMz5zmCGzGZARUh+4jO6hmj34lS3LjpzkKiE7iRRrJP1TKa8CPpo1HUHj7TMfq
6WbYIEaSEDd/KX07N5kHy9OOLbw3Hys3zZT9mV70O8Uzb95rstielolLDKQ7SSxwPQeveaBDx/ON
MJG7YQVyL16nRpXZdRivx/qhllvFUCL8hZe4ZouC2V1kK48YWWzljL1R2zMKmnIhtJmx8xn1zHeB
FwOxshmQzHQax6cgujdmIv4wlzjnYsfi9vFY0ejOPeKfJD7SLZqoH2NCKQ2Us1S4ctMhvGFQlFC7
IhUwSH118FHJoG6GWOAcvNo8bmtoMOr074YoDRBz91C9jgOJ1wR/1aCdkXXbAbPkoqduOVOBfmPZ
Vi/GNJ7+nYTYgB8qGr3ovzdGyupuSDICzBkHEeCxo1bst8769Hmf7CwKVMILBNhFdDH/c4vfBuQi
/AnVnp5zMb5wLR8mXImOvfDWtcZ4J6aLrx8z4F4JFxEnH3cwx6Uvs0uw5B8Il0acrIlSgk1W8aNr
ruwGUPxaJM3pflaoF/NjLMuTwhD1Fo3ZpqKlHOK51fyi3P7fQsrSoh/7XnFNbt8gY4RYEES+qOrT
wC9Ir06ojlIcFPmub2pMJSn2gZyoHgLZrwXXVXm6Unh91MMeTfDpEVZsiyCJr4CsN9XvXoMQcNrv
GCLK8N2x2nlxFfRGuJZLS/smHP9GvKtVJZ/7sFNMMWnYAKrLW+9pdtfxV36LWOhiImP6KDEggxAa
aO54QiGknBCgiLW4Bp7EmcZK7Dtg/+EnLpFj+TLc8cM/BDNpMIMY3OqOm39OgkCsgjvepDOj2GbE
eoZjlty8GH92aH+gwjSVOGEkN891UpRz07fJ9ixT7bysFm/3U48WtetOhMpQDhXrkjLHt1UGDLmh
9CJP5mk47fds3D+fX+EpyGBSxXkYl3XFlsFvGWmsSDLQ2Wi++cTMB4K9gGSaa7R04ZAkoNONyoD/
xGejhVKAdWeZAzVfWp/EZJv+g6eguCoLZ8if1K1Qx8LKfMAAhX8TJreV6c1MdUqF4+by6mPmsUI0
PQ473cuYIRtTtfKEe129uHZwEst6oLHpGf3fLykNVivF9ge5+LPSWi++2pZNzvGfjmHXtgohYfFk
en5pV4NjVYRHmbrI1bnsAoUk0O1LtDC5rONuc7g+XS1+LduQbiUm5nmjFVv9MzSXKuUekQ1TjDgy
np3wIW4VcZhZ6rsTntQR9BLDki6UzNs3jQ2urpbH64u6IA+RTiwlk/dsGvBfP6qfUzzYtHWr9IIq
Ni6kEOIBmQ8fwvvQLkw06cPx+NHMUTjoykzsCpiyHce08/1hbyw4QgNuNpwDCAGR14Arv3ilb4z0
XcC0AR9Z3K7c28OxXvQqXpfNi6MgAcNE2d6EOVBBBpUMxOvpQ9gjkSUrncvJPRc7ZiD+M03jJXP+
muOuX+dO9tGBGKsgSAhq4SahZJChhxxRx767xa5gNLCzDNODlMBu8ISFIc19CVUxQSseZ4xz2ieS
rvt4hEW3X3Yz6duunyU9c5GekmUKKZ9UeFD/0AeWxtA9GjDGnwSEsd8XwDq33wcC7p1vTC/mWzoL
iG+wkPdm+VpQfAPW8F6ZpQU++25B7vthmwJ2ePv01WRXqGsNJr4d/IvDpFQ5BLWlGy7kdRRwLFXu
+Fcchb5SeMEDpjaSw8tQ9JyAVaDMVCmnGmIm1dzEK56bEx/AIYF2+ZyIMhfVpRrVg3oOLePUzlJL
bJq24pF5AnzmqvK/xDx9MougxIXSpqTwCk6ds9GjeWpjmbupkPos2566jw/RoED+vcaPVeRhDu4b
kJPPKH/OwTTHN7olgkZmPjheY5B7EoZAMu8YJrNVYtuExh71KCAL+V5HTv63hBpe7/3gKWnEcejb
OfZQwi/7DUixjqqnwPbV3/a7QHUxAh93XZ5/N2OEEVptv3Qk65vKMNQW0jHvT9i2A08MLZRvCjgG
CMB+VvlxWKy4JOEwoJbLKcASlnPtjpWecsmQsGr5hxbH5pBIudnVLgV+7tw6AyEgh1Ef5+wFhqYA
tkMOWhtVDyZfQCkKsE+Rc/XsAjTP6w5/wf+UCWo6e5iQaSXXASYs7q/P5uKeO5d4OEh+xTZPFPnp
XcHMvAq07Rtl1ARoLWLvVyTKKrsgGt1E5JyOiUPSTVqM/SvoPsQjNV+ifSTy+SgQyWLipRJ5TwA9
YjWw4hL9A9Ass5d09e6DwFC9pZh/2AK1A+1Ynp1Q2vFOimUlZMfPmCgRcLOfae5c/2VayMk0SHaS
7h2Ud5zE++MpFJVrbYU71uMewjh7P+2I6/x34ZGP+QQmVZ8VySW8ZEznBhLJi1TMxiz9oBfCXFtj
xEMbJvet9aWMdjupeml9mytX4NQjWSN0GYWSgzBoVKn/qHcZJ4Xmd/3JqjkOJCPHgqRWr06mLPN8
74fINbdQsJHbAa/1I0SRn/QNm0YrC7EmjUfd9JSoV5R9jwVq6B9dOLChxQSdtUlkk7BFxYO9XPuh
uMu/b0rxdOs4Lo1RG81DyJwHiDOcjDISq0LRT+VqaOIAWC2cEWFAd5O2ZkoeScX/Z1c3TqKw/XmU
Er8k9BS086cUjh74Kxs7sjKNnvnRU1wccud3to2IZu0k8FVkqXKO4A6MJidKVCKcH5LgUewEJpJw
NzmUkYQq41nMeXdher0v0quo35bo1GUpPnivWfoKN0RsqtJBsUN/5i+zOp0YMWYCMxoKaFL1Xqq+
YUVtFBM9AIwrLlYjC1hzrVpXC3APrGpJAA+X6CSycGOS4l/KJ7lRmZo/TqVB7ilh54PgvBAlWMJ4
nXWAGJKkyKyRG/uURdYCyVyrfQcBe/uw7+k8KosRhT1ocfw6rjquYVGs1T1w5VWIsFi3SKB45Gnm
IHy7TF1xbXrdcQSVaARcYrpXQjMgSCcjmMe0mKuNwm9mq3T4GlNolfvq9GLiw8fHKq0FdIxL9GXD
OjRWNOz/1e8pj2J3WZlXLWoOatp77t2V5hpMkao+2EqEJ2QqAXHjNqLI1CgxjJ0NBrAY5Yr9DqY9
GBOQxkPbi5m91UBC/d2AXJkd3irXhdrsG/fuEkQaF1UDEQMwc5VDKNUIW8zvJ++X/3Z0qjjvcgqo
vMPOdlqRNv0+v2VUKG4jcz+WhqduhyvCyOnTE0pM00biXe4DjC0lhHFxg5+2MT45ctE7sjXzscaB
nXSjAgGj3XO6bFjXB0G+iuzOZ/RMTpAtmx8rK6Z6qT50dnGUOg9bcVPvoKEniMiU2Equa+eOrOqC
FwF1KPI4d71M63D2te/orB81cDXzmgHjkpI6G3AlWM7wSHJ2EI0buPv8VGJQbdBQihl2kaWOR6Cj
Sut3dz48mF+CaG7UEWl1VkgkkZbMmPEdihOJ6431w7S7WpTbtV+UL6LwBObEMi7484mF4FwGEZzi
T7BrLb5r09p+EZJGBMh08fhqhE6EppBLKOSU5c9n9JxVrkxlhUUOCvOZv03dI6c3iDgS5Scyo+qg
VRg2f2vVAPcdGZzyXi7exnI/DyksqbiJMcxOs6gDz/Zjwps8QQXFJt94Esh7QPyWe8Ds1AaGmJ4R
siKyrS1ebzNcPTziqG/yRR5U04DsF8be9d7tefJJ8xcqjlWjK0mUbAsg/mqlERHXD8Uix+YrJG+4
PvsKK/1TgONE9S3qTbDfknPdSCDnf4qEP9YXtNBJTu89qAlP8TLbI6rtFjR3fzuvlJ/bpK/1qN0X
M9RgNtmn65Fe0Y0L5J5+vz3A0AP9Kpr2mi5a3oKdfLlpOeEVKmTQkvAjv1jG4Pu4NMVRPJnCluM1
Csv80P/hk9MrXYF6p7nmfIUuT7GiB3y49bZ0L6+btP5DBWtxGj43SuV4Bfk70BBDYOlYNp0NFf1V
AHUGQ5czHTR7hxVw8Ai2j6Wts4pyYk+lhGpMJzBuva3/2cLoHcr1dV8FS1BECxaXivziebaw+BlR
odQqJHkw+qnE687N9EtI0fU2Yn0r5MNy0P4qMo0UZM4qPj4hzycLGENyzvHL9RIBuy4OihYCKb6y
alFk3TT5+d1VLoBZnktCgQ1W5RY6nKhepXovFwYBdufonoseVJW+BSwsDqEk+WOvwHez6iGQlhjJ
IjV3gCPP6P6iz7t0Mx+nk39y7nZf323cZf3+sw8HRnX2qPrj7jLUbjtvpbJD2Cl8Yyxww8dpqdx/
M6Ylzcgll1yLFxCCYY1zv3/H5mTRJLsRU0X2nu4g1Kuf0q/NDzjluQIWJ8REWK/tgmd/m0EY9ev1
OpGhjS9xL3HyiwAa5oy7e+OZRCgrfI9TWzEhY5BJgKRkqFidFbPWPyHW0Ay+Pl9L40BmDXPrkdoW
WE14tLi6vBGbS6/5INSyWehG44RIA7t8F9HJU/ZBYxidiUjWi2yrUISwhE6u4aXxP/aMvog29wSk
twuHl0Zfjc5Rh3iYO122ny7/jIIKhff8VlpmlWOTM8+MlNyvbLO/a3lGjcpyHLpHy/G0jJIjWPrN
XtE8WEEGs7R2Avf6KzqXAfQzc/RTHShZNtu2QqpBF3Xk7EhVvGZxRtqc6tkL8L8LFmyD3LmRQ3zU
QJQTtJnhOSi4AQwgsgyTYdvJVKlqdixYsFIbruzHgfHNw7L2Dm3Vyjw3XE/CMcd2cuktdVY5Yb2z
tV63UsGzxi5IUyJNLt3dPvPVMtFlCEdT49D65EHSJxg0D1zVclSja8haaQ8e3cgTNO+Ag9p/8/TB
T2QZaH/pLTU/r50PEkRmh1mhc7QxfZRPbj41dv7zHDJGlVH5PRTh8qyjmWMGbz9TNTQUmeacO830
9sE4gyND2LC5ICUwsASzTpWdkpEE9Z5MovbBs8Hhc2HO0w8Kp+l72QZGx2gL/gev5u2dqU62d0l8
gdI9JXH1yV+6Oug96BdN/+vE6UfI/fKTCrqwZ6UcRjlxnz4Ziyzzl+HRVwK1Tq17/1BuXphVVr9m
yGcQxa2eYYP6pdngmNBIq08TkP13vf7v2sh9cvFOpLGXu054j55BADeIzQ1LH4C2UMKdWLuNnUIy
Tjk+co78ZOea21F2IZfPXjm1zQ2YHH9FEH5S+tvuOHFmfAnM/cyuLzWZq/YRbkIjJkaXjs6MZO/j
RtI/uMp2SNDk5fCcq+h3NPwQdcQs7ZFIBjSSasJP35MbtxAxZfNM6NalCjk4KFGQuCB/ngAqdtlg
+EpacAvBIoGF3EADKCs66nryVHmN9LvnuMNLyZXMdQoBShCga5S34naBgfgCwG4Jwie0UVoRrq61
Xc3v9W80VfXVQ164sHwZRbEgqy0cZQpqPeW9FoeETjMKyJzM/8VbFCsCAFB0H3rp+iJdvcfYEp58
PniEJA0OiO1FyMsqlgjfZF3P5mNrd2GQoBuQqFXie66SoToXejVETGJMnqb6L0gQbnmvuxL9h+Pd
zFYanrqHkfORVkKRQgeGJamNXcovY33mk/wK7I4tKAx80Jm+PvI9T4qf6+orq47h9eEU5GU2H+ft
bn+rlEWm36XehSgOPxzR4WqDI1XfMHjvp9lKX7Dkht5oxngVTsTwxjZW1iQcF4a9IVzAD+sMM2jX
AcRyEjDozNjuCohXwcvYauVhvAhnmGb82HBWvh3e+NaLa0fOCc8fAVu2rphf++HErZIp/bB++fBU
8+UIDuRlmqAjLEseeity1PVSh1ce3lwm9Aov0QPjiDIMSd19CEb4zSIrGRuo6sMkkweqPMJhaL2Y
SH3R0QB5iANbsEHpb6i4OSyKotQ6dAqWiX4UsuFTFb8vEFGcHMiZsKv6pVd5TBoEIppErMhfSGIh
TFQjlhTwbVsZ9vnuWGR6xB/UWLJMdMMvi4Liw2GVbJA8XH8A0pm5xmdqIfizby5OOXEh6CF3m1dM
/CpoV490XQfPGhfDYK2++acowNzlosKLihNQokscBjwJWa4o0HhEvwuljgWO2jnzXWBdULrRKdi8
aNnWATS6cdqaoRvFMsHEEpAeyADvLCS1EQ9nLFnKbQvbxlJvktrxTaKKAspMIaLV3eRhxWF4tbcP
xQkNAPOYekXEKZChLs+JhNJ+/RJf1df+DYJwnp5VkQ+T9fJD9PZFsQDMk1DnxXoGQCshKW+A3X3w
3PSXxHw9/GcKf7DAZQ3Aox3ImGKe/9GwsfNWGn55fHstTS8Ngqfvc4pM18x65BjoveTLhMvOHiTc
0S3bpP3w4Vvyl9nRaJy4HyOZ0XCYX3Qpqia0fhizufzOO9s71Kn4qO338LX8M068c7Bi7Vy6pMdS
f1L6L6TgwNsOJNTVKczNqPzlGFcoAhc50zhlUnFSaUKDS+FnFKmCw1vY73wfxZoOj0z2ZDx4dbJX
AJJnxmH+89LC0kZuYVvyVRV6f3oFJa2lD7UpG2uodcwlDWMn+3C3ooDbzV/orroQ1bns0Srjm5Ap
u8w5VT92m0zbKOXkK0KkJRLm6hGGjvvg/VxkCMao2UjHNBqZ1HOdPwdtL+z7QSM1DHDgs9KzJ0AA
VuUdhVSwj7cken8kN1/975XAi/mIFkF4+U8etGUKbEK2Xm6cxB5NFDXUJpfzbctmqQsIeN5NmzBl
AjN5MdbjOjf3dbRs1gzOf1LVixMWz1TSO1rIFRBf9UxXybrpzAwAuA/NoAOsEC0tfKE5+akyxARt
foWYVRChzXPeuN8UAau46EO7ACNZyeLxzqyLHL5bEV4fOemIC16fb9LoeIHVsBypc9k7M3Z/fAm/
R+lQ7Yag6gPf83Q4r/tYuj+N/KB0NTAlPpZnnHBeDNSyO7KR/6d/HJAw58vMjvisxdDwme5iKB5K
FGBaO7oPoTx4kYCIXDkhYeqkCKjkbMQGDzAr3Ikj/ms0sWprFiJZBV8yt5OvtJqFdXP8m444N5cw
kZiLNbctsikJ5gqGEUqZ94bgGqUCWrfyceVwIX0qfmDx0Tiin+z7FspEj7peHyty4ms//hj8qrfl
HmDPTIdDNrDj5plzENzwMOz4c33Vf+HXNEsMPYC4W5WXRhZNoygMziOdvXWARl559zJWDSbIwGy5
JqKX9Ozx/ft+4FDtQmpWPR0g341xcy7hyoYI7HQGcKSiJx3qwVWhg9MDZzmwwF/oV2Xxj7ueXkmz
RxVJwcQJwi7lbrDPZxFvOxxs6p46cQOrYxHK+g9iOKpGIV+evDUATlLor/SRJiBx+BA/K9uWGbvG
VM75vIjlhmtXCV81jFm95B5xeYTQbITWlVm3MY3pdR/uiObaXehqjsDc6tnB7Ay+j3p8OxWoJAZc
qBoMUTvmlmjgGadwLkDzQSJb7ETuShLdyRbbuUb+DLUaMBM9Gjy/+G8O/StmFt3ouQII3UJ4uvjL
t/ScmzKthYH0+J3Wwd1pDw4bekW9ExEIxHwuGsa2H5Fak3ZGhmi75JtPEeb0RIzW+yRpYQHImvD5
XmE2bWA0NjvBzaBNAwcYEV/guaNSF9HNMSZ97ebbjwTFHApfk4D7fq0f2hjsipmHMmZS5OOTdRiD
saNw7B0S0uvEOx0ITT5AceJJyw+21UrYp4vBnYReafV7MLTcn2I0hbddT31zSoe2Xzt2hcp/VqGA
mXe7j+CzrG1rqwf3p7bG0dfkqr5ESWEyuqp/GCbKInFNSn1FRY2b40Zj7XxMa5WEgEDRxrDRQYCy
3WGV4Vlwyc/Pj0F9wIKSYETBVpbp5C3nVFN+fIhbfXlYSWvJlvqm8Ybr1fUet6cmNxTBTRY/lFfF
3Ae8wACEx41WNpSSKKrgrVQSOfxhAHv9xM0q/9uDTpvkqFiEqZ27ZT1OSDd53EJVeRrnjWP1m08/
CQK2bczGbQpPX0Im7GcfZ/MpQ6k7duZ58oD0EcZMsUdOhzPt1RUgpXATMIACmtMDMLZ/pU9zaK88
5F6mbd45yBmO/QeDtnCJ1nOK18b932UmBT/ZkQf537f+nf0jZ51GBdEfkfkZ+ZQ1MYZFymdhFrCx
bk9CF7iYVePyXKG2psdrOy6Sc3Ib2JshNjBawWSO/w1h5uIs6uwE3JwUYu5KoMM7tVrqpkH7Fu+T
TwPvDopaodJV7fuWtvvCI/NCSXNx0QdRF/cTOpwW3CBFE4JVP4p1oWiTfdvc68zj+LW/cI1JEEXG
gblE2iNcNxrBnfFyFUjlEdJM9mTs3asadpP9EIeLYRsh0Z52gs9erHQX2HLk3RNR5owJ46Qvduc7
yorCkiPuyvjO8pU+W+5EJX2dGudggS6hWEWcHxV9DuJl8OB4IbbiW/wf9oAVHQRIx1bZ3GDoCfYt
1myp/VC4nX5dVZVfq6MYZa075/n8/CRu/GAn08H4lXkIKakrhp7y5P4G8oVkNRvclwRD+wSMNbgg
CE/zWYwU7jPDfn9c2Q006BxFODNzhzm/y3jiOv41DyCn0PAO+tINTMLPPy0NY3FfpJ3I5lkQMJ/m
j0aBYjzccKmaIZ2YVm9pJ+mv2YLGMZNoUmMNhN3hx3SXqm/rL7tXXJo4cIQqyMI8iBa0upUT36PZ
vBzjE6y2mFpZ/fF2tCr3r1yGjZRvfTrIxTraESDXF6EoHPU9HVaCVM3zFWrCzX+bX7+RQHh7DNIe
ERT0VAS4g8aJy8ZUJl2Yc7AVemRjLdKaZlF0S2skbf5DejslvbOAANVn8oJgEjv5fnFLk2ZKO924
kv4+6o27LoyQwgMTY3KwA/NVOEXkIQAkYPv4BoFA0SV0ei7b039LjEbD1c2MXf4HGcI1Pi7IWxLZ
sRVSKTDoXEU//+Ryt64eTxiUKj7e3EJNXg32FEs2pM+qLlyca0XvI/IzeY1xFeVshxW0i2sBaMPE
6pYyEJCxI3vXLJ5N//lNzGWow9jOxD71mBZU0z651GmaY7iBJrIfIY2Zka/Oy46KGkOt5p7bUUfA
a6l25lFLwIwVXcJy5FBfzFnk/EyzuzP4AGvnn87bUGrG3YcmCcNaXfjlBnAY2/AN+WY0oNUfeF9N
UMz57R/NjnYfnfLGBYW4PXOEjiCjVcOV1MggwC9Ylv/2VCk7E89yVf4qy5pn6WY8AQIzRTPe+3Ci
XzPnuc27Vq52Vrr13znBUEUZWrPKgKB7sumA8nZ3XypOaBAzdK9Xk93XqjLlHwlL7r/Sf0N2ZZ5E
/RsOyJDnF+Hehd/uVTnScRZKBAAdR21PxPg9jL7wQ+OPyUs7i5PCRqJcNDNgv+tbXOGNxYVgTjzP
FZwgktTKGI9U4yVfbmDn7K4/veugKgZbBGrd62pc+P+vagcG027cyIPn+dzer6wk6HXzOkV0s2Xd
ANtnaPmV+tflo+Xf0MpExjEs5n1RE2ouZgAYBiKQUGSEANWh1zt/9X+0JPKVVHPJg5ri2+R2RLJt
LZG3wKz7tqvmalFe3qrMxkrwE2ddt4++WujVS3rppOtIOUfVg59sML6SJByUUj+eDMbbDo3i6VWC
Kq/7L15WKgt7cgjuN3rPfQUrUcX1bBr0EG1PtUJkx+ttCbDVa7fSrQ37ZyWRMZCet81RwL1Ddm8T
rBMVOYJcSpo1abYmaJcvUga9Ib5A7nnZQmHlOcGxIcZYe5EY5RMlG2LcJujiQBtXXTtEl/SHrhmW
TyRXYepFmZognkLmbyVY2lPqLX2moSnYqdFpx0KdqT6Prqb1fUZVWYSZm9pKC6qyJ00/eMGV7Q+g
/XwQ9thUzxhM5qMyqJ7t9ZscAnrfVTLRfsBQ/AKXJ+V+wMxJRk61nQEYSRnxU/tOwY5kC3FrXnRN
lOhW+W/2rna/D9tjIhOVVuNS685nC9H30Hxxdln50FArWTOhl7kIkB/7RHLP4NecR0g+V30SWQsc
BoSbnjA8QQs9MbWMG97AzFkHFPW6+skO1O37fEEheqXHoFAQuSB+WXH2+NuKFF3j9JEJHc6olLJe
wEtzzM3G7NCSXd9n1rHr0lPJvFiEBYrzqfGSZoyEFhnZK9VzfrgmrfygK6qEZfPKvPvtPr7tTrok
RX5wUnZsI0ftXZW1GLLdb+fJdvv+LmqdKB64CWbrOIhHEy8Fj0qw5hUzi8W7i7u+uI6CUBq/KCh+
koU92bMsnTaKsujahR2Kp9j2f0tRPqTFKFccvky3pjyFFFFwi/51P2GJy3OqbWyVxULnVQHxEBH5
wMAtiS6ZoNVfp+AvyQsaY21Ig9wvKwQLCvQHGzp+977vhEpLJYLG3yHIUN/VMOMLewEepRGvCaHU
jCk/kZyhoHBbpKJiw9Iuq+q22eD00alzDqGgMiARBySWXHuMZ0PA44UcPthnba2029IDCS+UDtqI
LkgoQek/WkvHwC4ZjlWPLrofG0/ZNInW/BdrgQYhBoTClEk5Dgia4Nuh46nl5PDmcAtaUzZo/bzw
/zyRmoaSMXg57/ct4ugcQTSrhBpPykTwzp/wRzMsH9/6TCtSEZjfKFct8prPTHL9pXdHMn8f0JjW
g1ZCnmgRfEHrVZpO8HRJU+n7u6N4XCw6BvPN2+W03ahIsAzY5g1fP8DUZtBtc3d6jigd0+335xMT
vUgFQeq2Dua/40R0myIFdbYux7/4zLMvA+2kerHFeYFCiIx+uulQvzlyfpx5g0BxuP4R7ZbZnuU3
RbdIOoQNt4a2iWb4qMSLJQcRiffejJ27scbHu+B9FA6mZTOlHRDqWcCuaZiK69V8EmrDmaffcYui
9s0L7PWyy3BVA1DzLaTIqg/z88j6C7UeAGcuQXN/f5uk4gLHRtwB6YIMki3ZGeMyqwVOfGyeDmT5
bKH/7rTmP4KOGWBhTvPbkesGVfvEJKIeY0MYQt6s1mGbk/o8DzzYZ/Y/ZJHNusKbZVHxE4JooYy0
uwISmKaNYji//Y80GEFju713IZep3e0FCQ8j0jbzXhJvDb6oLV2HgtzNX5KXPCpsO9O9Yhp2mvke
qFCMrccO1Ng2G4gb74iuKEDeseAREtd9LG+oVKNx5AejsbcSdZfvUZ2QCsbLjDcUMXDByCu7KRxJ
v50X6Ee/RAPOeKGbMMuuQGz5L2qV6lphz0b+TcPoDWiOfiMVUzpX5DHA0Xh2/chL8BMpGmW3wz7E
j1IVQ7ffd/1mfdLtTZ+cIoSWroQgdZlD5mCvliW3ZG03xjduPwrMr8bgCJxSsKRb5JVxVtpp1U+1
Hm7OZgETHjUm94lN13n28xPisI8UR3sf0KgnoCrOayde1CfPWfdskUk28KWWkdHfm2bXaP0baYyM
5JoIrTzMOzOQM2oSIt42cz8sUDL7pV9KZX5B9wQv1erfKrroD18iFo8/lPZ15U7foTt1BrTGihid
BfABzhhx9BydXYbe/i6D3oXVt4zIaxrryW1NYV7AZBCNgCuwQWrf+5VJmxgNwimppsq4Uj5/kQxN
LCafElmvbD8Gup+Dfkc5pywxnqhMF/62GzSLAcOVV7cICcRZl4FysATOaVKgdi4VT39PCHDKnb8I
fXWyqLIkV6ZF7ctRahP0AmtPOcyr1f6nWkof3UYrmLCZbmDex05iK90QwjTtBAkhKiRUONztxm7g
Cx3d7zT6NJWU3DZtg2zWJHIZOCjQQlb2NOMweYEG4APYHHep6qey5pc/bqYCso4FJAQNW5saotXA
o1JPinr3J/bwSY/mKCRO1S8POS+WawTJGMUxqzFl0AKm7GzUN4av+TSLW4YBniZ32zD9ujMFuHx1
HaW6YdnA6sO0OGr93g+jjFby3DGw1Hwil5oD2xpmg85a4zbHP3fd0h9xdAmxNGsoCNRXHwO9kF/x
8Zav1ggmnw4u1KPfp9e/yE93eL8WLBSrBGtokFbd6oubDo9cU/iuCt4hfTWNVmy3gxQZpsgeGMZG
OXwIBOv6OyMbmkHhQAXsykuRIgrQuYEqslgBJbxoe218009qywRD9R3hITAAvqyW8otdEgCF/1gC
PubKo9LnXoMMxfT1WnfA9hyIn/OgkL5bt+tpabZdr/+fY7G/egTY+nCQUbMmt7HXSPvgoTafz/+X
9gCEXwFfsQkoshHQ+ooRnD49fA07KPnSpPHXOm1De7f3/J0ak/T/qgKj+km48FvjJSAnA/dFeaCc
Z1iWvHgSaaBimMPE9oeJGPFehvtmN3dEkJtq+cM3dD4gLMMtr2BBFYAeYHn28eywoJEeFs3r3pqB
te3JLZY81K9SpJMvuxiocTkb7NdEqnKAOFJUy+QJSdc2qRFlS159tHXAEdRM2Ax87b660cL5lEy9
vnXNkkdOY3FZUTG9n24iCcfq7rtleAfGBnzkxQKjLBdxIOeBqRo69mzTzxRwKNUsXjm1ICKFoSpQ
V5RO0GsqZEbyPHdnqOJM6aT02vrWz3TsDhzGxtn04oxyxenJ4eM3i8P5xzXshN/MA7lFB9ojsmAk
x5PSTGEWVbSWndlRYluyTAH2va5nXyBT027Bdvs7sYiIEhcHUfAef2D3nNLGWyM46PwkwvvEYI3p
788Lpxwg7f/HugPJ0XbKaonqwwaWMBnaYiJGc2cM/WdekkgYMBIbSLc5l50v2BDUc0c/cCkjbq0X
n9LOLvFj6OFVjAkrjlAOr77f7P8z47DoQe1xfGQ/jTJusQVoMlxvK0zWVToDGV7SaUqmlFmGqCIG
1Efp/ZsAHpHgEK8fAoWjxKv+BpFK6LMsz3YqVsRxCazv8uArYjymdybtmWJ6G87o+Tj4c9snJqJZ
fv0ia+NHa6ei7rayAfMVIvc6swBlb2LkZfybKK3R/94O8NUtOb6tieeletHeYIdd/DLpyWkGdXSI
PNN3vDC3QFQxBynFcNClaxkqPQlWQ6mlN4Egm0Y/0fW59TLQEAa9oaQ2BUMNYS+z8dJtueDsDfEH
Sx5l3Ov1Be/oV+Gs2ZnQpxy0kOZiRf8zdkER0w/cjnxIr8sJzUpvojaK31w/DMialKKWCHRJSjDc
B3VW2iwPuz4QoiKoklAuZC0vLK+/wVveh83ISiBB+IRp8KMtpPwdG4hxmNS4uQ3rs7synSeIrCEM
y9YOzgOvz1ckGwBcuKOg3zC5ikgZvf0YgNHVPQURxYU8O+dPW8G+pj7x2Ib5WZHw5MULJe+4KwyO
xxvA9JHh5u/fiW8RKVLLsmI/fIet8WBeBfNiTkGEYPZWd308RwplHLoyZECW8OXDeUmLl2KSUnvQ
vC/g400KKPny6c+/DDpDZ9iPFxv5vHILKDuU5wpXfgMmbPVWLCvLnHneRgta7TLYDAAj+IByPdK9
uOfDgYtZvJs6PO4Y/4kEBNjHstf3lrdYfWP9v5npinveGB9MVlbDp8kizGUhwp+OMSTQBL1lqCk4
0L64JvU/rdraoAAT4c9fAE+l/q9zhT7qPX7iXuu/u5uhjDYKMkiuX02uG6Tm+x7RA1TY1Z3MnOBk
Ls1FZzIr2BOc4BLkqQkvpAVDktzaOhRk7pDMrTf6lEdwinzuTtjvpwMxRwvkII2KdAfx2lTQnuwY
DwqD9FvPcL/kjWLd0ZWgzMm9DW9BOCzi7JXXbmw+VqKIpXTCpiMS1Xm+vmWLQNuRtT9k6h+6UiFk
v41YWzO+qRRabYkJqDtY63uoaVGxKcagE+A4XanCda5JDRbjE4YnAl+v6VSgLOOhGASiNZXu3d5+
SE80jiJZ4iSmzo5HNdizmXkERn7uZ+V7t272mhizXkaKCQU/QMEFAj8XfZQTXmc60326fH0vJBf0
xwavZTwnQRj0DbbUMJqt+qc9LpSoA1pHqmQZ8muQfDv7SWi/kDWpjLZM79V8U66kZC2mAXhlAn7q
1p8MW713eQWyIz+x8krM07Fk+v7IznjcBKmCJm9WiXnEwAb+SpZnRRSLfLq6Y6tSPAQTN58XDMZo
61VQy5EHqV5ExzooZrlt8jVbgMEIwLPqurR3W0yEmuIsvQsc7einU2gttJtNCeVLBd51ohPVw1/M
vrYazs5GyXZWmeyYZyKKP7C3zFBjSG77vsL9PhjljoVtFNHzA23HVDnLC/hC5W6SvNCuT4dWVx53
ufZzBh1o30sSvQF+DIchX5pQzUSDLMaa4v9i0rEG5Pgo4SwZM8+nW2cDJB/wORu/IYTL6+6Jljmn
0dtcxYdnO9cPK6E0ZGe0WEiYYDWxXUFwcVSDPJhcSUL/pOVFhDKM48wMRBfCiTc1CkV9p9NgPdYW
Yqq0CXGpXvRLASPenjyInuvln7zkh65B1/iHe2ygY6502PTTdO9//sZTcZkXVwEhiwWUTAV+IGtj
+gAHhDzcAyltwegKP5yoRw16EgXi973A88fmePuMhYCWoGNo7FO1t2uQWuXI2kz0Ij6yu/CzNtlG
78HOHmCdhyviifwwUPeIvYxGxtHCjKzElxWrfW314jmlrkycv5LUl5G/h4PRBusaAKdJ2stpxiJs
/yX3CeIJgjrVOgRiQD1Yn+guGxCwmjpBTiSzORkqpJhGTTTlEYK1M9BbLbcWapFFo8aa8YyxFQkt
0RgZcVgQyahNWvcfoNzwwtZshPrcWcwkTRt0uSv2QW+buMnmh6fehslF8W72WHgC3RUGnLEd3IPK
UEVMd8qA4xizBJEWKuzUvTyD+SdHvxZMAOil4NBCNFwV8PiGW9Dnj8kkLhMS8PNl0VHk4s7UdFE6
zEiWwuSaxLeppah2LieIK/HL1AKwFhuwfFK82D0LvjUKgvnF8KDjC29jU058HyZjDqWx796wwlBO
GlA8S4gNjYARsWVKmzTQiUI0pQdSD4AHoDhstfxNBh0UowkS+ofBz4K7OCueZC/AccTyhHffpcZk
+ybz9xm32U+oQGvsYtggjMP9VPGD02CkYC8lSkZ3JaN4SmRGk2IAqIDMCIJKOGHVkxI0C+BWMXz0
nOdmvZZ6VM+OH3CxKrogsUiTZJi3CQGceqnUKCQhtfAokwMp3oT5q012uRxsIu2KJIxarln/2OAC
BQ1IT387Tbqtl5YnKGczS2iW8zvBOvClxRBJ6xb+jdmym++gQBBON7TV225L+S+Jun6Thsu9nZpA
4lllUGnTWv4SyTEVFdAyPSSCLAtIpIZfJ8eQt8nDykdAZNPqRrLhQOrPHnySUZmm4OrBTFMRUTyw
gGef409rvAqVuKt8MJnWJXoVrwdfS6ww+o3+6C1KUTvuOh4vUF+qWfoIrdEOUriDrNi0/PXoJ0ym
+08970sl9ZBGmSNsV+RdhCUSIQj84xdwNoHipW472HxmV6AhAJzpDK8NyZAyfuZsH+ZWkYEtYIe1
em/eBysZeV2i3Dom4pIT8wYAjKE6cC5eBnaqHrs+8Mxm+6fNcVPXHPKsq/cq2jBNXMSb3uXzkIi6
4Oe/3QbE1TPFlZsayLU+yxVc31YYSZlvMIgqYWvlLXGnOueYGbFaZxChn+DlNHtquxuV7S4Y1a6E
yUN8M7zc9VBNCumMzwqsAYhW31dfBE8tR6NllHRYnZ7Y947IlCYav9LBjhet9uB5L14OZhwiuYXj
LPf+Wu2J4ZpRlUm3W+PP/82H8M7XoxRvxvCbjsyWhBm9GOJVO2hknt+VchUkoQOY7T8hIqTwIp/j
NAhRN9HeKvK2KvkCyU7vKmWmT0OdozyM4Z8OLakA5BswclQUTetgm8eQgUk8Dj0n5JxaoRU1tc36
guFBmrwD7KwwR9TrnZKJ9+0lgPMHpZtekAeugSbB7A4Xo/cX25lEpnoygU94rQT4Q/4pzb1sR0XD
aVkDvS9kZEw0qBhgs0T0v+t195d7/RszSDS307ERbjZyIvyD4Eq9C/CUtrZ378qgFTatI5wKb15i
wZydbkMTibQiJhSLczr3U6eLp69cau0eb22RazEjhrYCiBxEFuK3SIA5RpI8kG1LJ7JHMDFtrv+n
vgVnUOjcuVCy7CuJBN0L34SAEfukytqArdmaouAYUS1K50ENl3UJAtkIMMC0MXEUxUYZ6xkUHsvz
qAt9jyq4j6ErpP0aqQ5u4jEKM38eqHRXMn1Us4BL8y1hJ8mGcZBvYqp4JLAoGTTt+J/Xj263MxCf
OWFHo9dMQwZyMreyMQr61nPOoLjDq3qwnCWoedDYEWtofb/76m6eL9rAtjDKFhNhtU4RU8Pf7BEv
0pDUwz+in8ON1KwJxS+3QTsPr/SJJM2JxYbyJUfi1Xc5/zSK/axiywmso1JSSIF0m/5pxF2BwrSs
bnRZ5HfYQv+d1AESqFybX5Kc2sE2DnyUXEUQUXATa11uEJjlqzDuMdqXO8/rmeC5BvBOsL2ovTbT
5uhKHbbFIltyq9w27cTUUof4CCRGx/L94GaUBPgWNQvkGPo5nBHas4r3QHXevOJMXffXMA/0/NAS
EXoaPlbQm61asEvUuxjOXoYygYASW3TNRKYeh8cAPbAuiO64Xgn/BPx8JU2OZ/f5emcRPfRxKffP
i8uAgXUNZTc6qFCMKZPzo/Il+e5gBhyWT4u4PWTW+ZPULcumdivNIJWg+7X+WlA4AUwBs7ckSZrb
VZPCJPtNmIILxwLAaJISGoxY7F59e+YzSQow5hoTINyuo2eHp4iei85aDfZksIqzbOWrg1lFub9/
YSaXkCvThz0djWvQvwRpIJz0fZxuVObNZ47UDVftLjNMBanDvdmSCIs97yzFRdt9TKnrr/24mIzb
64zlJO1Z+6Wc+hqVQNcFc/qtJeA5CzTvGh2VRl6IAfCOkGtKDXN5JIGH99T/+CXUdDgntOVfCyEa
lo53FejkD9HF8t9InjY8Nyhj7AECBwkvl0cpBrdK2XtvItunLTNmlwqzUKo4QhlfFGQ8GtRyi/Pv
I64ws4HmR5dOvjPYruCtZ3VQid30dVn5/ZQeWf4SNgaD6BPw46NiRcFbaa5Kz7o6Eu4Ihc7ZLNc0
UPN2q/uQVQIu+0wU8tvc0SiVri6RtoPlbwl0+SgSUUdxR/OLlA8n8tGw7SEHHxs9r3JsujzrYE7H
b80T/DSXD6xQBRV2UuSjui5sjxk3COFtnlwpN0jLkQMMO+bgjdlQTsHT0uqyJ2tGtwJAFk12zGxV
3280YfjBK0wcJcFGMbTHHJ93R38DdGNhAv6u2X2aCLf0zPM3ASS5iLjLHk0b13gUXWVxVGsjnUCi
sihZdYgnhExhDZy1BGQGemnntNfCjx03O6Zqg0lu7BuXKOHrojG9mP2dODp2edO4eektKgjnQ+nk
azDbAECxe3SHV+R6nqMFZQ+bKfxuw6hoLuxLDu0MLfMGscovV/3wa9gUN0Tr+d/sDdruiGQfgoSH
hze0zAII/5QVo4iDTZrqO3FtA9RtlgU2t192GgEWL9w2UyQ+ahuViIUHrUViHgNCFidxviOUpYjL
NFO7rkRKh6TBgk17E2O+8fBcchVHxiqksrZ9p8uBfuWnUeO7ZXQ/38CvtLKtEyyxRweeEEZOmKZw
U+cUnyil0eCSztizduTDqlxHl2TdVxmoomH0hyuJytcK8MYGlKmhjxYHsDsHvW5EXYllqOaIDJtt
yLpCGsrOzWJJHPCs5LWGkyMqo5gzQeh4k9ZpbSe83GeSfdYnDTuLMEovty8OTkP5SDeehnKRFDjZ
WxMkYsPIUn5AC/UuQBEpShX4iqQfIoU2AR+4rWuhGIyrJpHuCVHb+/HxPgBBZeQWtwyXFY3a+SG+
1brwcDaL5n8/PCk++U3qQfMaEZNp49snvvbfkVQvwigxAohdIY9nnsq6g7b360iZDdhnuEJvZDju
siL/qgy1mPkzZh419Z9BI++7KQTfohmuM9Q0ZoeSXsLgxPi422pjZWcgkn+2W8Hj9u5huourg5ji
DTnSTLCUEVpCzJLYP9DAEzoOHY+e+TWWGxp1ixNlYRacsEij0lGmplkcHaHXYRUEmLJZ35iKA4EI
5+vMsui/G9q7AOvKPE3J/ilfvbY1mjCmHroA/WDETeGcTjMuZyxB0UGYnusSIojk+kzcNSpVgTPP
/HJNaWYtrwUTEK3J8k1FqhH5BEdQd1wIhXICEaqndh9hSRZZl+HOp1YCHqKWYqtpYrzvj9E6dLfZ
lC8l0cIMjuqavtdowDGTiejyI0nrUof5EBsbWwQJQ9IW+LeSQSlRiVzLIBLKDbRkulTuADKAA8t8
m1FKN11/HSvpV1N/6ra307dYPwPISydU0ssF47bWJL+B7aIwulU6VBKmhjBFEUwXd2GGXOZ7QR5b
VkzCML3Zu6meDG+fE8tL7gGhYiZEAx1TFJktsmStIMts975sTLzKy7niaH1gtqLK8uwfBZAy5Jzz
0qj+LYPktZm2XAmj6izEIMyRe+fTVepSaxj9HJKXSFIqFnhakvs9r2rhMfAbhnm35ore8gfdZ+K8
6jvvmu9BoIA1+iBqO/EUyrR8ZDkI4iJrsxJwwPJjHCAWuUzDfC1qBIekEodedUhtONVM3ydsTRD9
k/gI686ZhQ7nLYdXXPO663aEREetWXFVqb9rTN10Do1tNB/FJY5w84jdhWjD6Q5yeVwj6r93kyNg
POUEb0KtHyu6HpRb7H5wh/r0ZVFHMY5hSp8BcJg4TebT2EFqT2fLgwIAfQ0q8kKlBtF3FmHQ1DEb
gBT7JmGiUfIn+nIW4WZGxCRttGgI3GTZrs/bZE5DvF7Cff1K63LaaC5br/iGjfVGG6AH+Pkg8g/s
X28uqhQXYeLGN69QlMnL11ar77d+hiMlbehWwfrCaDlsbAXTE1r6crNx8rt0MDzOJaUd9hX1A/LM
Rl27rtA7FT5ZV7xChZ5tPJmy3fq0h6MyZSr2FT8Dm4p1ezQY2zkcUuR8llHru3ARRZywrJLYW3P8
BluU2651h1+zjEMj8BK7qbEVXFvMZyBFIzE/vVRVtcc2j/4ba52PVPGDwZ3pbeW/l0k4KvK7m/w0
0d3gl1LxgY2hxVRGIk3qxNVao3QfeouD6bI8z74RAdGmMouhUbqPPY9hASt5cgLvGVazwGhN6vpc
UlarFbiU3busBau/qmJvxE3iqW71UK24SQ/fMfqpOM4iOplDmyRnk+2e4jb8LJeZFzwCQqfIa2Qh
de1pm9e7xZIgIWCRdiF0hNPx3BzKcg3E1XZlFIOfQlh0WdqYYch/lbt784H3VwgXIUm+iRbZ+HDX
S3440ybgon3Js+lrXIOO/dT/6PCAkfdJydQyPtl2O7Lb7qvUdWkIW+Clr1Oz8w6Uj5VWuoCXTPiA
xkbzdO06logV2fgoTXzmkZgTyeX+4HNHZOG6941fC7HcPyH5xxvyNMtNbcmwb0eW7bJ+bhWAJ/tX
43gelDy084wJmZxBAhN2SkkK1UtC29fiYQGsTRhOI/XwdChhQGGq1SdU4Z875yABC7+yGFP8+fU+
puY5DPadjuxzATH4M05+m7p466vFlUW8m89V9wP9pRjD2hcc9724cUf36aOvK8LlPmpn9docu1hG
rBlELa2VbAcj9Im1126o8vOd0Io7JafPOTCPSVH56U1a2frP1fALbSlsauly1RZ/AJSDGU3zWrKa
uGO7fG6297YEmqCIX0CtNMiRFK7jYR0uy83vCfPWeYrHBYIsMioQN/XH9hdMbi33vZFitPCnEaHf
YFft4l16cSRiwUaksq5/WGTWu6lcSEqZeHvPdHNPWXkYwFeYhnjDyj/uRJBaLcU/n635MuUZ0IQW
LdsZQTLrytQ4w0CFSlSmCbWLdsUEqhPLKDrwurPM6dmSiU5D4U2mKPMAqofAxA1S7VUX6lh1d1FI
LDRahoV0BrqHvHvl2MuawzP6XgO4OQWwUQe8bH+pGs8SrU1JSG88jUMeBNMfUUsc7Vf0flbtLTWq
jgnS4mf6Rgh9d2d31GXS4Eiy1MjJadKgdrhuz3V0/0FS8XRKnUv0a7NtVU53p69SKD0q89rs1xtO
hC+sDarz6Si4ZevkSki+NvhfeRzq8Bfk6XGAFZ41F8SNY+Yn3qV9kjuGnwl27bi0ZgoAy1JgOf40
rTg/Jup4V/gyL0+SSmenZHlrMqulgmTCT1p4lySIbP4XxMSaMSjq8wlnr43f0py4PSuEUJ1xUPP3
gw8qQYP30im1b3acDPRfeXZn0Syh7XRBRk5XlvO7a7dlVQTreXBUZsvNLIMAFEXUXI4en1I8Vo2T
aKPbVymFfY8HS9egh4x/HLeOxSzOd/du/LpYSOv6CVSRWEsfo6iy1jkhAdOdfA8qQLsquFZb77dQ
LaoXkO/fP+WMx0IQ0mzAV3TpAVRkwnLJMdjkYTK+IjJX7OE99mvecGnaR7HWBS8bRF40um9+VDJg
wnOOAtDp5X7il7B41PF8MwTp3EXADd63Gn/H6eyKnTHreMOFy1oVIHRFEiIRnVZoSaQDR7/2eR4X
NyLVAPDliTEIUEJ3jSypL4QadNSqp1TpPU0flJFinJfKXDS14rPNXAYy0GQMAqN6eIq9z/6jAeO2
SUn+EnETscSgG3/yqF0/eDeAb1t1X5KyGZCNVHYQpFjaMo73INBpka/ue95UNFX5WtqTvnfgPb7I
/XRKDBXbgjMqsBDDUmMRYiOHJhEnoYMQLpXsKgW1TgUXjrTlcJx6G2nf7kCsE92RVXYHzKbsK+8q
B0P5XZumHVaH0LCLkQnSrGvsx1H2BIIycYpgUy37W0tarRJc/9Qog9AbycyMHO2QzsxLwRDWfynZ
S1gM32UuKjbC3LTmmLPeJfDjBDibWG7RcHyzTCveuyXbliNXjBNm5MCGiowxRLmCk3qqwO2sTs9M
HUWjSHFGJoClvU6M86JcO24oCn3A2LHUs/zOkUmAGt6HLzE5My8Wt036LMY2CRg2Rz8b2nAXKj4X
1uoaYVC+o7HkUbmCPL6UqAANdW5IvHLv8QJ/6kWkeven1fMKMiq0lDO0f45Y/TEmiCtaePMBpXvJ
YsIkhjB39pcICXW0rIo0buu2AlskdRhaPVrYxpLzsvuG5+nHu/VxQVxiRwOSVdHvpiGkMcA2/Rul
abuilcHWNrySvpPJqeKUnwmpXAGu+yFZh98LSyJoxtXnnHdEH94xl7KMsQJBboNZ+8W+WpOfcSuu
YNVvtrdFKT0o6dc4k+fFiwhmcONjsXcE2jql1qf5zY5rSNnAdkjui42Fj4fuixSuXYu+xAWJ5eOW
pj+Bgk+LSNdOoq61gi/kRYuj1iKMmVausHdnF7MecwxBvrkaUbCjvJpesBTpuXM9ETdnV/IvRkdW
Ohi2cq7/T8roQoY3GxVDQC4q6cmGDRVbIvKl7z8BmkaeTnnjUvOELnCpm76zYBDLS9fldNrayvGs
9V62Dldtr9EoXFAGq31sBBiEYdFTMNlqT/wa1DluzPztc7kKGrVYL+m/mrwgJ3AnlET/LfTExaD8
u7ggzDNDy4MQfXG8ERWG60vDbp3ExCcJUT37KJbu+3Ot33p4RJmljsB09DWu5MuVuPNFQ8RDF/RQ
6OSLIw0KNgQgKJgzxoJsDWE41Az1ZwwXt5EkN8VELeoMzwYa1Y0gZziFy7zQ7OknCfPFzRovGEOT
ZRYu+IufY+DqSFFcHo+9VP3fY6w3NV47ruyApxvxsNSpQkxmAT5hMIXw7sa5JqIQ9VkeNm2euD+a
phtNgyjJLHzxLDOlywKYThP/J8U55v8sWxTh22rqzJDUMvmuHGvYaDbwqipkjlA+7UiPsjCXAvTi
oJOM+0gcbPeGr4POSOdBZ3+PVfyVvOCZHzfuKvBvMyX/iKvQ7nGu52VjasPC1ph2f4oN3kMGKPS5
1OiMG+r/Tv26ovVanAU0ITQuvq7ToU+wOC8URRmgR8Qc78QofyrowxGYMxQUztP4WiTk88JvYwVx
MTVmTmxP1pgBdP78Y05NWAE8u46NbtIYg9/Y6DU0hsGm0Nco+G3CgkfYb3bt+RDP/BuozHTfbH1t
4JS3fjPVZOC9zf5iI2DnSGlNb3xSUZFurioJ/tTVsdwW+RNrDyYSv/3bWSelg5U6y7FhqePIkS31
M7ZflNAzYAjCJVEHpqh2m0m08YOMWeCshtwoEFCuA7MpXvk7V4tpzNbFbkdjO0f2wf1SBRGUTQBi
t9WYnbVmdiaUU8tIcBPVm7O7MIFB5tnWZBPtHvheDR5Sh+V/pJaRRM0/aq78R3vjJXIaK75ha3+U
IA+bFkpkSz7cXr4kjHBMakcPVFZY4do+YhQJ5cViIhjou8dJAXSH4UrEWe0zaoH/KBnNVsErnQxB
LrtUrM5T6mm5wDMVkCZJyZ2q12/pAW1D9Tl2PV5Op4XEPatGSbj8EH5QNFFgqhm/T9un8s1kKik9
ZOgwmWNBv1X1KUm1TICySsIQfOfnhgRvhdqBhS7Dmq9mI+P/BKxIExiYkK70IqfqjSyD7Vn7tzum
v6uHGKzoikI/98s3Ou/Vy1EkGXxWH98ekuyhZ9kkU6i/HCcg++hZXEz05PPe/GVGoHpAynsNyCxA
nUO6QZ8TvxexggVbqI0Ptt8DCAtp157tLId24XdgoS3iVlk9XAk+UDqLVaBKhQMq+LFyHfJ7KgIY
hp6Donm95NR+pGB8bIQ2iptbSwV1+wtwAHwcpmMv6VpTN1jIjUmyZY3T+H54dpq2nrrmKF8FZoDn
v0mdYeMKMAKJpnYZa+Ddw8v0tBF/QxuNJ41MBaK5aatuF/XgTHHEewBTgo2ds6aG5qKYmfIQ209J
K4vsEuIEErWcnoAU7dZn3+E//5Ipre9sZ7bDBS4rTlttpDdI5jFI+J8ti4dyWAkf9w5AJzIZ5O3R
X+qDSK3kuTC1vzKuGN54wFv574OBV9dYuh4y/dZuyvTWW/+VI3vHi5rWIoGIhJHHyny7Y+4ctF3D
7F1NJzY9VtqZmLAVhjIB77ygno6xjHFeZyOy9lJ2r13QYxaLmOkd4TDD/VHUHOkChiyx7KBSMQyj
+olvLRv+npRRU+HbsTaFvrzz1aY4WzIxTgqgHJ7JnOIYgiJ9OEwLEcM8/bCUbW+wlM+ja8n6MUMg
HCcfNkX9MnybTjhpT35eOzWz2VrUbmcT1dg5Qu2avKhhi+rhp6lHTEzWl+DF4Ggmlr8yY022TRlJ
MFTFQaMFkW+EwQhjkc+pDs0HQftM8APsYVhVZuJxj7Zucaa3YZ8kEvbZrliMvaV5K4+uS1sqCCdL
ZxoI2IjJAOiIA89CDeAweASGtIcbkejIbN+oDnt+xU0j7yNzfi6378xRFAx7FZGPXpjX5bzjRNka
oaqPeM3XVwkI/zO0HHrHeY3Dy4GtjXcOM4pbyHp7tYHDPaYZibov0/A00C4ziMBLeagk4ZIMwDiu
2X+ZYEG5/TF04hb0XyV5LbWMUNQKKkiePJRtbU3YFuv/HhaacHFNuWTdBWoFZK6GiJtE14surugc
4EPr47nLFu//i/D3/GWhzNnOFlJWoO8JAjft5AuLtA23Exv+aRHo9U2zYTzeo6nEV6pdGfppNf6n
5EbgOSiWSedvKzymSODek++AZhnXM1olMk2qT82nImdQ//+lQn0MRpnK6aanKtz48FuRJyJvEVmH
2gn2trUukQzRISZCh88aCw5I1E78rpddfbdbIw+d3aCzlnKkFUF+vJG5knxqFh91NmoAmj5/KowW
ufHc/CVNYVg5I4T3kZtrm/iZQDMyG3iAyHUxI7/2hUIZvSH2aQUTJP7O7rVtDxpTkukIhgxXdgES
zts1QOo4FLtra2Mc8O0Bmz8BBTdHVF9r/QlHDpxR4hWBwGwXDsp8okI2fJKuonjAq+6/IAyx0ceZ
R2rtciSdCXzlyqCI2fnqTjiKU9ot5yaA7Brt36YxtS1s+UirUHnfzD/6mp1tlD3Qdy8XSb2n7ETc
1r2pA13uGm8cn8/DblD+tdAk2WxHWos7ogebBIEiuNcMYfHGbqk3MQGEqzaGbyeE6Nn5fG6jT2ZO
s030VEiBzPttbbvglwRIsZ1S2OtlL5D13LRM901FWfC6TCmsYulgRiNQjxLF2XHWGelCL63S4KK8
U23O4BxDuKXKZwO7dpOCa0J9Y6AwbreVx18qNFTPWIKg1aDWddc1x2tLJt026hoj88VxiCkaco8j
48ZlMxxF0yCsAiJ2NRUu5rAU7/xnOU00BvMPq99zVZ68/d9iZzHFga0uCD6HUtgZ+/CbwhLyIa8d
qhPgsu41q69DezAy6+khgX4hPmzf3MPvIP5c8BEeMYBVG+bMkxoFUruWgM4EFfyJMeB+Mux4SvQj
R7z6Dz52nWaXsHhbW+2hMuXJFz2iOlMdTdSIlhzkT4bbWkxshelsJ0/2g+xwmKNdrxSkOjHSedII
gW/8Xzeh2Gfi0V9gwFpkF1KA33R1vh54k7zy031h3qTDkpvWLXucTj5GlhrU+4bd/lqIrbbGKFSE
COjkQnpBZosgDD3mHLuOxCUZfS4Yk/fGpIvzaGxEONZ02YTD2H72Pm/saQVADTffqcpKAUJXJt1O
TVDPRK0rsPw0kH0nuwFqSNV7Hweh+p7D6F3PXACclmNFjoFQfFMDoAsrd8BU37iXa+hwaxtu5W89
jLsWeOrQog+hUi4InfOEeX6Tx9fHMWbAZdyJHSET0dFWGn/ZTM8QvpQWOAcXhCW5qQVTUtbj+/hX
PbC/WEV8f+F1j50YQkpizgTZx2lDa3Qdt9J/G3mxXjMsScv756JV/qehojmaxOl5v2MbVhZNMg1r
7FdVIdgfe0aBAm6KbWcEBGzJHaZAK7BCvIA5t94iyQrRxW98EYi7N10QvY4qf9ZVXMrGBcYx8Sey
r0vsIGmMWotOPRA+FSiaU6A+BeSn6r/nm/2tZO1gKDtJ98sVkHQDrAck7uAviEY0t/lj9bHKra7x
M+HXVVfJ082+Yhmy4GJZkmtTvphENUI0oyUFTBQ4ENL33/2bdWTO4mhFwrUmHYVBAS15bZHRCXLF
ZF9tF0sWaTmXQ9YpKSxcyuuHBvoiGBh5yLIXrTdkd+CLEah1TRvUzQuztNvGkGA6OOgu9sN/tksj
gaZTJGwFO0rC3Jp2BjFEsdKzJKdOi/D1tq7XCgv9HGfULpFjyac78gk84FyTZKE3G1rnWTxlFgmV
MUQIw+ux4WZ3ISFGzScszS7ZAV6uY+4YayACP45WJd2kZZ/RBBVLJqQUxbOuxzhyH1JXsnq36Nzf
ywXYMr1k/6mcyrCVJYVgqmSX6mREWsNoq/U5XMk6Lg9B/o3qpFyIoHm03LjWl1Mkngzt+d6O9hag
uLmfhs0TjJbX9GRJIeOddjm9vl1JRCw7USPspO/PDhdNjLFKCnHIF/5PE87l4s8iRrlVqUI6vLC2
AhWKLWW9bg4CX2J7sn5wa2UCMp+tsidcrhEy+OC9jEDKeJm7TkW48HStm9/ownRpFAlDk2BEd9Kn
D1sO7Rf69+ECyeoep1j0ZFO7LY1ZjCFFpWKPrO7bOP6F3EPEE65rAuW3sQnup6cqXSvDZPT2fJFf
QFvpP8OAha4whNya8TFlY5cus59Z/CjCeqSb7GDY8BFVCOhi65u/JpDg99RIJNvGoD7d4Q/qRZuO
Aj8sGO+7G3MJphczABLcMq1Hcj9A0XaKPHvRVo53DbnvarymhA9abIPJqpyK3LpqJJYpCufMEd0e
8zj1+PKm/1d40sF3JreqQhnUgUMAfeL6MGj80Kd+CPcGLvVttt9lydq/wJcjCo4epOc4s2ony1Uc
wv06R9NmTbJFnRUGeN+frI1ocidrXbQDBteie9q/LD6V3TFxXLafDW/Qzmi4pmqmVS3eBkk165Tg
3+ys/M5CdaLOO0u0HjNSHo+FLH85m6n8JHsgncd78GwrlAsbS7wzMYV4tLJeiWiNf3pjdQOrsDfJ
1dCwxX3fowt8fZCKCRgxa7U14fHiXITusHD89Bv3daGE6ii3+s77T/DVrfBuNf7bYmsj6fMkf4Md
C4gexWqAgt6/3hbCWmhvBRLi0Gg/T5LR4XJOhh7YormBwfVz2CFvHHQREjtkvBlTMwM6yySBqxRH
xTV+rDVT1dcWeKefyNYTIRa6tay4XLlELA4rNTiIMJL3caWlS0wPzPTa0mJgYwhGHkadOvzr1zZ6
NJ2mCiSlVwZYW7Rk/wS7fK9kS4Dz2uMiCEfUd0F6g7yKEef7tpDeHD9aOJ+5frAdzvj/GZhVyN71
j3eOpjth2r9tQkDZytSR8arGPuBNqmwh6svpB2dZ7FRy81wx3+hiL8s68jKzqQrupTLeGB/oPPfG
D0KrpsTgfj9AFXL4CgvHjgMYxueg+hkCIkhG4n+01hK9P+ueRtQDvp0KBxUNBi5n9YBI8z6augyW
egAz+TIVivsQ3NGDg696OycqcHRKGr+SZtV580XmA/c1HYHLKm+UjKtNfKMPiwzEn3yPP5eP9ekk
wgq6SfMyOEMopN3XFlBtGNgWPrJxvHrs46jVddOJMZSjtuM3rWZhLk0cpq4MtQMIhqvc1kvp6WgY
TZuvv07F7LBlQZ0CFg5jldr+K/RwGSba9HabNSeu+n+4PUkKQwxFUYvHYJAAkdyjhsZo2SVLbGAL
k2Nbl8HZe4h2HryF+PRT/vk6731FTXGIsDjJ0p+J9Y9OnLRTKZ4rSU888M45yaUofrdrrxjKWurX
JNnJ5/k3Kxj/0Wet5hlbFyS0x41TPkfUSlcm0kyu6LhiozEx1zX0MX1IbwuDhXOhcPIscQaKLlVz
Ac/MHgZd3Ex8fJkyEfl8Gjum0Gv5gbbirXD5jVKdEftWJ9dR+T+wx94lDEUxC6BYbtJKaL7sGyNF
M2lvlKj7/0w3OG1KIyio4sFFxvwm7fi9xTLtFsQKUuGaKN9fppALy7IM6kNURKW2+Q6WjWZahWSn
b7rBEEy7sj5xW2Tg+XbKdC70smwuP08iP7ElRmpkfAjSTwyRNeWyXrj7iBK8DpXxW9OEQtaaseF+
h3izUWpiPO9M0Xom6lsDZwUccKYJbMoBsl+PGw7UukdX8smiqSjRJ4I/wO4R8AHDcjt1J0lYcU0e
BupmCwkqrOISytRxDV22eMWCWxkSVQu2MSq2G5GM7O4/q7zmZZc9IaU8l88Qa6km8W8/0EZw633s
qzsLY3p90cZvC0PaC/wCx50QwCjdubMxDBS7mj8LaIPFYFriPfUMMV0RfET2pu63X259i1AP0L8F
sSyAyKXR8/Zbt927eiBpOf73000PMoOpqLyJj4UQ+IYngnGji3FMXExgLe56YSPjx+G6reVC7KoD
tOzmRTeyaQfNsQDTPkmoxkoeXZrmHYEEkGRPG3HbaeuX/WcTZ7SWXI4YIXWok8eXTX4HAFvTcuiE
FxPJCFu1dxbW3umfrzP141trX1XjJjhXkB1fW7m7k3mdyJ5QAdhBIxCdo9SqPLjOBwRlCtLaUVoT
JjTlKQcGMhYJi4JQDpbK65u756uBcVpjuPnO7ZNUGVGuKxg4jugo0pQPsgfsW3Maa+ffxbTkJ55b
EFlLE+JO9LkSx0y0e4f+7L98eh3DjXojLu6S93TrfEGoicRdcMu3BFGs0kQ9f/RXJGZgdGMVfkzS
SugR7pBtQYaxIGrsJzq3gKmGM/AgxoHaDwJWGUutLkabCiXmUHKKCJ1wkXtuEgMLkgPbBMLya1d1
nXI/l+0bGdNZMoW8PGrNHfhfKd8vJW02XUFGWZpFLerL3DZKh3okQcGPVKO7sxnWsyqE2DPpD0As
1NTvgXA3uV0OMR4RdnA5WhXEgeWglqoyFVz9B4L/0Ls8mA+16eQaEtCspavkBRC8YmgyuN0n6GAI
iqmRLTLf5uajT6CT9gGidk04TPqSRVOaJ56mIkaYKDUZD25c8mMhKQdM0TKFZGrnja+W9gavL8wO
j9ss/xEIEF80u/U13FJM/qoUNTsoQmbUjABr0D1WKYQzyCAkzPSMKboGprIpOB/lBML7XKuHrapb
EHWPBvEfnqdxM8N389zhI7eUHSHWnUR11Bfvmqp53veikA8VUO2A9t84UHpdwZ4w35y6uV8uzz2Y
8yOHuFHrhs7mAydXIjrN1qS9KSH8e77KuYaZnpzi9g9lrlW9z17G3WpZHOTVjwFo+i3v7ngZqBX3
WcPlJkE1M/gfcZzKtsu4mI9FMQ7fKnIqdN/rb1OHZD09dqnpiwWg5/mz+xwPlIQNRnI5812uulOH
W5c+QBtlK1+8lq4bxatB64G/FHRQ+2Nvl/JQbPh9fW7zjY5c+mwlLFr6Ncfaw5CIyLka68IktxJD
rTr6TzfCXcF5I2OHYoKefTBgNf6WcOskm9TheroEmlj2Tl74+/HBu8UWirZ2t8JpMiFK76BDU9av
lc8QiuiAFHiKd/LmK/Xt8pfEW4vN0/y9Obmpwyjtj1JVeRMUG8iv9QsZtA+uf0ShTeZmglJDceyq
s84bWCtekI6jbsYEbW/NRMu0KfRv+yYC+oahjLDQYbXjQAOqQK+yWiravPd4LXMkEyZ5zxu/SPyI
6+zj9hK43PLZg4bV4tWYyr9qC2NfWQ4UTQqeiaiZ+dO7GTIcFLDb0vG/w6oozfcL3GwIeyEDS2IQ
Di5V630lBVstmFAxoMXuweyY3/VW5ENryNgFTw0Jz5+iEDocvFIEJEPu4BDXBmbhWyKiDQD/oBj9
pTbnPlYSuWzj+RFsvhRKLkSObCUUwjWq8j7xN/I52MsoJbGQ8LTIoYn72uXKJft8g4OP4FMVu2xf
vmfj/x000coNvTkp+FFZ9Uyko9AetV+MfIZ9Oq1CWCIbQQbNMaCx6SNrsl3oE5graS25GgIvkTcU
w4VsmQHukPBhDmB+cFNfbVdMKWINbm0zdAseKPvR2bKt9ZHHojlyu1Ps9zub5J0Juedjj4vx0EUu
t9fxdMbD9KDRdC6ErfSyrDtetW25GO3qzyJ6VUo/WZPiS5psoiri8VnsSRB2jAJET5njdcsjfIFW
d5i2okZt3zKglHzSHdwNwPPyV4ne3mtNU3eKpeF7RyZ533OtxHYBx0pQbZeWircVBibFh+J4WyOn
PjXTu6WihFuk6AsI9Kg+Yt28d5dwQln5B3w93MR5oyJHgLJK6zOJ4c18PHXKGT34Yi6ayHUvONnM
Daw/aMXrLZINPwwM63Rp3s2QoVMreDWEaXtylIxcraFqfqkXfmhaRds9ypY53XnQIpbgoZveP26a
FQB0+iIh0b1GQ/b38dAvx8nwdXVX5lENHTSez4tJ/yCZt5ghGuU3GgUJ0xop6OglS3QfENMDi+wo
Z+e8EWBwMyphf99HX98MOUQ8RvvrpondMUlIQgHDx1ymSDZpjH1edOo+G7QHG9HaJkCj1QsIbvmE
8tGf63k7ObePYjLvip945iiWgvuVdUG5QTJmEf0Hh9llKWQUw8QyONxqpanjfAQ5RfaRAEgsfzbr
rmJZPm0sKeO5JicEPL9KPbRD4He74s4uHcrO9T06gb7kw5c+NS4yDtnqjbb9LPb/1mtMQS6yCDO9
zXi5hkPcSNAR/nO/A/IysGVlxHbVpkopaQQ0ItbFi8RiddqAnB+onPSrv2J8iKI3Wf/jm3C+zYEj
bsnU+WTCOqSLqghoVRd1VZgutdXvvtTL5HlWaurmyNwEIgRwM7tCxdJB/d1dqoDTAMkNXAJObSmx
gaBT1t6BNCDt9wL11TzWJobK86tZ3CsNFdZOPfzuHpM3FtjCX3/h3J73iqwId1UlySJ/XX6aKo4z
Or7PyxZ3NVB9ytAAeSuJG4PBSORz02PYCBuFwYZ5b/SDLlAh2k0yQEscFeJ0A/nEUg+puw89YTuX
1D3hQFRfPizo1NdGqwdHQCKZOXpqgWK168zNoYmT4hGeqD2WzHpUNVtIV8X5zDUBU0jDqIvrEELA
ymhe9Z8G8iLjfw3MBb9OpHvmVn6X/fw875LBw8JiakOEBKkcGwHbtdIoQ8rxF/6/SQ/anIUt0l1C
KdLM3Ixae29QXXXmECVsLjRUWE+jVFj3jkiLwNqTvDCpQJ6R6PbZ3IsIeutMZqbSD3TPRZpqu35g
IBcB2K2rb/LwHNJhrcs+f+wWwOn9jd1/fVEd+LvAaCcI+mIBC4cRlz+1HtoccLWArph9b47TYPSS
iimM3Td+kCCddbliMryM5eJj3PaCRAeGlt3/St9Vz6TN1z+pU+o0Ti6JECq/S1uDDOyihxHziJ7j
bKp8Pxa2ybFsaMejAPSvykdByEiZg5/vOvBYCx+9fshxHEuMnzW5PmrYjhdoFqgWQy7cML3ZlHjV
v8fPPJrUWoZ+vE0RLQHUgxUkavvTgiMJbm2f8z65tNAjKB6KvLajcEywq16SQ/SY8OyiqvFlfCs7
ixNsVKppk87LzqWJRW3GOi3+gPKLNXuzLIBh4LKYOrQxSw7R0mGc0JdACJTvTIzwO/6piNJ7W4pF
hQkx9xrEwccpRbd7nNnGnknH0PcA6enP66Fn2DKEfE8MLLxdpFhhSThcYzuTOzZWMleWfJvyqjgU
NFUs1nDbqXSQVjmcU2WTpEHlYiNu5n8ZRtWy3EZLwsl6kH8aUd5j6gHVhz+PvTCz8Z7a6cqEmCzp
qDMNLbm5Qwcw9AFGXvZxmN8tVa3YQhAPtd+WNHLlbP9O7LmPQpY3UJV41iQb3b2dHFx8RGLXA1Lj
jdNSusZm2Eusoe7iHeN4giySm660DJs1CmOYGPegAVV0tI9rM+ghpEk8kl8DkIazaiNXzbBv6Apa
MJ70AMX1eLByPp2LpzkQc3JURepvrJAXwiHeHJE2Z/v/0mWzlHNVA94rl+B/0iguNMWzet3qAueO
qfC6EHn3c1y5+wutrZ9nYUNVtamLk6SO69m//CgHzngmjUgvSlJQlnWOrgWH6cv38mt/TrGdd6yr
WI5PgxPAM7YIdlf/v+tNT5giCWIHSZyqNZ3n5k7Vdj8TN8dx6p25ZSw3S4OC5gpafrIr5mVr6lj/
KgwfZheKqFoKP+tV6F70gYvqPz+maLX5XQSE3chY4zx9F9+ltyBvzja1N6OZU0iaVjoVqH5YxKgN
LVN1nAeLo55dpD6mQDYaZpAXJBrWNbuWYzc9hEslZ9eFtwgHjAW5sUk9R2+RHi/zA9D8V+mKjK0T
qfsdYfTQm/ItYhtuyNXTV87i7FSVnVHq9XnxewpNTShJ3Ao+4d6ivv3RHLrKTvtbIx+Ja1BDZ1BG
JAOtYrIvQSJO1H6+IpyEH3goBGzk0kGo2SDHcEzdosuv8VbpMNxtQMotYZ18dVsFLnALSmE78tCT
PNfiNhSprbxAsyoB+1H+F1Ab8CNVWSNordBYEbdEiPlxvk3eW87zEhMqMlAVwlcgqlcn4lUl/jzR
AUoRnvUFaFaPEzdO1w7QU20Qq2oybvz+sTQv155RRcS551hrrfbB5nwKULnaFIMyZwEOjPXMmZe9
/sH6HsrE2d5FPwb1OZn6pll0LNf6VcdwmvgMYOAys7ANWcDUOLmRo0xni4yBsL5ncwlJgUXO4Qp6
8PMtOUUDr/xSF8f900cl5ZoZ2VUOFZrsTJwSvK3yu/uCbN5n9L4l0bTH0UhJwnnsnVcoR3cj7VRG
Pe80XxYpWXxuEAx3EDDhpBDLqzv1CESTXvJig9jI2fC5zhkxc4fVHx2ncEWrZV9QOAKbklD8idSI
L6gXbm5HwRVzIY7Ixrhe3/GH3HtHNh2ugnm4ZWWx2dRM1Tgxnofgs7psMX5zxCD02Pw+UBP9JJs5
7STr3xOw61ZghzyedtnYWDyVyAke+QgQY1V37KInfAOKJ10T5f48MEVTtiHF7RmylUcNw42to9pm
Z7ii/5grfbVQeVaRNz1rG3KuFdGThSg7hCe2b7qB6BCtQfwwykqy7iiT0+zlefM/uVryHIZvxYXh
wBknlB3bWDW1M0P5AotpY7bppZT/7DebBopU5HOpewqjXOtxa6UWmi+mDn7usFQ6UuRNdJsNNzM4
cqCuAt8uIEmaIhZcBKGWWGnIrwl9bOjxKaquLsN66mtQaz2z4ADIkZDbFlBhV8PEfU57VzMRbrd5
sgT0vs8ZVnQnNCu3iV3jELUhvwrJoTE5oQvAdRQfw1iqMLq4LWryHzld2e/qMkWPc66FQ63jHG3p
nEw+w7YfRunQecttS/00GNNzQZHHmJWBztR3L+JGY39GDpyE6E0ctwyZs1yiV2R08GaKCddHLOcg
d8kXj0WfxBj6zzLYH2ShAzVUcBOsde+xB+tkRFw9l2m17xhkINTFNnqTp1OeL3SGXNMmFlWV0udH
2sBSXYfkG5xNVfvQaxQs+xIKrKCIA902bBthGLmEi+QikU1ZarU9pusX5bJZd9iiqOIOldXaLKHI
6swhLJM77Orrw+3wDt6blnaKCSzUpGeAR7vJ9kPidRfN6HIMUrU2m3/9wQjnLafTgqpJMiWN9oaU
5tTIDNkKNeyOrL4XknlbDK5/hE6JUni6eCkFP+JE4m6ar79dhfLTsDgAO4NTVzQWJtZnGcVugdCp
7sjOYosa6XReWrbJU+KB9tP0NIGM/RIpOOui222LrtXoAV2QMCy+oR8Xv6HKXXJBgIrPGQsORNL+
q2CgoAIAANlAVzXI4AtJYKZ9KLgYMu/cgGJxdPbMUHWCxXiF3mMyZDS3/y6kS97mW7uTB3ZhrUjg
IUnSesqWusaPGQdyHOulf6GKN0obcsdBwhGlJ/80dNkrfmOM9fKf744EyVik3NY2IfkKmOq+z3qq
Tn1Kks3WNssNNaJao3wmzr/KCYVnhnqS7R3OW1MhJKpLiAsME6FgtyZBDy7CU+sywSaXAQMrQVSU
y8cZsMLV7gdxW2HXYfUoQIJkU0+gt8Ct2xmcU9WZdS0yqFEfSeRt1pgYjHDeseZFVJWkj7jSDMfO
794H6LY2SGEhfKn2wwCS3mJmDamQ9tzV1y5kC1LDpYOu9sCXz5eH4I2uxI7Vu1PcRMgH8MqqOY9U
bvajLyTxXV1ePyYUkLv8c/z0mh3XFTf8+8Xqi7lI+7R3rlZm3UHux19qNJKSVGCz28oNJNXqwJtr
oOIsT5jV//aZuGxqy/vK2XsBNuwN0jQVy8lC6RGi107oHiIR8+qxemUQrfjuo4Isbnv0PiXTTGwK
HjA0ZxJwMZ7fjB1QwyUogxcvchB0xgPpE18viz9nDk902ye45KuXsaKpMyL+FM2lzbeHHyB/fsMx
yktxDZ1KA/tVUBXxuSL+JKPnKyB0lxILSTkggjhWjd7Cq378KF1/OhgNzMsSz2FDlA0ICNGs21Nv
FBGNkKyzTgP1FbkYD/1Q5xozcwyry54BqN/l9H6L3sjocfJ774hotYSa1ux8WcfB39KnPmBKh4Ze
8Owh58R/I7aw3jc7pGZxEGC6Iu6rKmiX5Ob0pQ7xOQl1tIQHrB9x2L25aUEvy7jhJ0Uz2hs75MQv
DcCyPyLxi5fh/Op2ivw1pvjkr0nqkhGZGjgW2BrMDMdXLueliGbu1EEI2EKUgRpPCVvX4bCW2TiA
5BOKPu0BZJH3yCO6zDc9NPtyPgI6HbeRY3FwN2kWsOreObIizMV0O8Vq+VIAzxJVHkjRtyT2tdjS
wsW5Q/Wu6rMub9JgsKuIsh64UnM6fjEpMMOltPCWKQEpmaZscsW29MUBdILW0jwsxKOU6G0ltNM/
faKwSGJJEt//fLQeMAZ55aNiKCYUVE2E3pPQLR9L+vWbcaZXJWJ+471uayOyfTfZ1zh0p+FMaLR4
zNe6p/WpZnCSMmbhIK6kkf1msVF07/F4pgzOfXM9CQ0eqybW/qb7dHpolSyyWaQ0738kBZIsW7PY
QqnZoEgeJ7rUS/u0WOI++XT19AqRM3tfnFlxTAkjQHax1QreEizMRacH0XGvUIADU0KAHaeYEEjZ
u3xSz9dG93ULp/1hyDFBgQnBuB0n5hqqzo81Kwrzym2Oz/ZsPMak2ifbXS9B52YHUXXR5fzRBxHu
N4gMm8Ap7f2cGnS31dgoiR6LZJjSxhICMJpTvL7IhozDZcTQTIgJfBGbxjREqLq3dyE1Gf3OzQ3A
R46TzqPMSHGBqSll9mNQU8MrEDoZYWWurC00AehuGSJ5A1U5cp++ycgqPNJKPvP48/HMFHJL+arf
kYwPwcyo3rr92dVgFPCa0p73+b8hWQLSHe/VEZqhzd86vg6YXtNwo94PQ4Z36kaGh3JsCuVc6XJb
vkb/VNmPxzv5apvMIE0G3EbJEtZE0xyACk0SNRgJNLq0DBrzjQw2CA/dNepl+KIEGxMxG9Y89mee
6Dg5faJ9rhLhs+Vnl7gJy53OMEuybarwe7mhbatkuFwUHKynev9AMoNzbT2aQzzH0pMsM04RH/Vn
1CB6nrFxNaqw4IeDCexCvzNfa9bLXj14dkJM7Roa/kDfaeCNvcmEqqf/KGEa1NwmLYyj88VIFSoh
kNOiFszCsb+OmaRJeR3X8aW0IpmYbGsHOMtObjECP7gl8JlY6ZtzuYjoLHtowZ3vMRpAPwbey/Uw
2VownPndMmhiBn/s+PZKCgNx4FH9StU2d5HkAffmwcAiwc2Ec3FYtUNJaK6WevLjmBys26w1xHQM
Q04QL7xxcaudajufbm4ktvvClgpghUzw4two5nBwE3q2hQp2fp44EY/4TptsnKC7SgYa32bnOw9u
oHUq7loXZ5407OWFqDtEoOEEw8S5qcM1BFCoonIflZQlkQd2RxKN7q6FK4b6p5p8daokE0RFNIzh
O3+tUreAqb/pEBFRYXxPjQs4G6nDywK0Ldq4/UNnzwrC0nW0W60qdmUs7qp9IhJeWxAl83CrarHN
vwx9jC/gDqwONKz7ILqnD0qyhmHCSpMiIhoYb8wXwBBH/rr2U1FP4i2pT66xuUqkmL6RTBuk+/18
AUFTBd7y3diAniceLFdTgwqiUMh3mDjsmTr8xYf/hRNoif9hcHISYuNycuPKICPAWI7wtVo/sQ6a
T2ADpczoxUdUcYqgxaQ02Mn4HlL8kVIrs1+u/FrTeVsYXL3lZUi0GptaTF+jUjfJSmhG8tByKTXo
T/KjqlXnyIBWI9e+++2sZg3XWPSgX6n4UC5uLJWA/1FMlOgCSkGbx+Ki1DmR5pOiqhrTBSFzpBfu
ytJLt27dKvhdYwIv6T3GqI2a/bZlySngAOQ2HqAKJ3k855M17YFqiGxZHV03PXTRRnD8NilUeSWL
83nlkIpLnk4s4hfHcDseMSXMJ2bplFe5yKydEgkuASrD6Ige85b7JlqHrz8pAReq1ygmaV1qTxwX
DYlDc2/HRa0jbFXLrun6ML8E0CjB1LyKvs0i9AUZCbfKJ5ZwPh4Lhr/4/YTXcJJA/VAfGCyY3aRn
gJEsp0e9b4+6PswEo/G6CLG+i3d06tXlabosYjG8gULcsKO/A+519HVkqyo5jPDCsoa3nRLEy7YT
9l11nhsRvTXDx3XUF5ONsUviENqEHuqzhxwJqTa/qluuhXypMiXWe724aAjCatiqTZG143vjpdDy
KLXF0LnbNsOMGB/wXslr9BS88/iDO+ZuL+qKbdt/1HgZtIQNQe/dN/u4JYK0KbxAgaxoMxKjMLMr
OOTZNdRWmBOdEAYcpEMK3wlcyxQkBEcofhdqJUqwQi4jLJwrNNLwq9p35lFG29eHRYbUmVWuBAeL
ine7M97VBY1LBls2THOBQBDC4xOGHOUdHNo2O0NLi3DGRFejUKuGtlEGTMMt8hoNCcnN858pC1WV
/CWmrCkIGofRq2X/5pPA8AVoaX54dLEXhumpVXc9etCP0LqQgUhOCwbdmsRY6B4TOGJr3bHHAaqS
rpRDYKoZMvhiStER8JIGFKWtZ8g4iJuBwM+l3711hUcEOqF9zUTY110s00m4U7nHB7IAjYI+dhMY
h4LgGP8yHQ6ZuuUWHx8dVxK8EtKW/s9byytbNfBDR0kikYfAVeSzGKghZA1/TBwIYrk9YYKRFF0X
swfrsQVchcIzS4o1WmmEB3hcnwpuWsU9LB0pqNv1n0+4Tuaedvm/VQrwlcDRLJsNi9XNBNbThRV6
OQwVL0ixE7g9gIqYHAyUTvOsOHK19KMn2xgLcv/Xi8UWIjsbw2W9Oi3gwuU6qWGj1U2QPcUCLLGE
73yY7lrtlXe0Ig11umx99ikglwWQ+oKpz8/NzGIl/sSV7XtSPKEkAmWdxQ8purVUlycOaeTaNoWb
T5+EnrYvUR/9QNXWUh9VbpJC8XzAZnt4RJ8KHzfD2nF1ge58X5Mmt3nje1+Cen5cSlpG+p9nCdmV
cQ5ocRbA/uNhu3p8RXKbWaFYj/BO3HAT/kh55Okxi+X4MF5rlZtPoVX8fYJGR45Ts8ajUTSbmVRz
iSJGAnIcxx0K+cMsErgW71yrgmkc1wTIkd/HN2sHIBlkeD6Vw+pHeIlvzeDvDY9pPuSdgVghSkxC
H/Oj4rByZ6dpN6Rsbq11hcgaCQwKGQv9lbtlwX7w7DW07cvzlbmf3h1veKc2gFqKIwyIDD64bvXS
ugCKdH4Fl/YMtnooZPWS0BcfzMzBQnWjSTntqVO/TMDVsnAQNEjANsBgK1T0cIidr2Yy3OL1/rRB
yvr2h30j6fy/L350dnXN+Za3cJcWY3U/68tsI6rjiZ0PSDit0V/LPmiwalw3Lt2deqEPXyCbGYsY
hXEz+cIpoSftZ0NvjPLrWk5i5L0GDjhlz1pWMATGp6AJNcyu1TuUKD+F78YppSQFpOAFeoSIK7ej
9hKGegQdS+ZX7miUU+52blGBAsJiCha4AbWqOU8yJfDW8GwBngSFFQedmJTumF95eBWcXnFeBwO9
Fkb9o2Ab2/JdUjLlB9u/fkx8lx1e32qCgte846ul7YHlM6o67Rlx3WbvFVidqAjL9zkooFn1COVl
DO62ydY+TsQ/8T8977Oudh4Q0OOCVX4R9lbwT9OyuD6LVFcdKZThbsYWsa+f711nxLfQpbVdsK/U
+xAf6ZCTEdtLCtXX0MRCQ7Bf7L7Oel0oD//4j/ctU8MrkVyHAl/PiB6ZWZ5r2eK4OKGbokj4fkFi
D4o+e+pSBXpFEkTzDnQYjyonQ5DA/EmXip/VOGxr/kL2fWWgoAbcRM7ImUC8WSqK7r+SkKiaFsdS
Xfl9gwn3HzO/ITjjUeVOqe4E7HcGkn516/BE7eW3ErFnPnrahhBdUNq3RpaVWk45hwnKFFzQXxTC
bFTmorIpcuqtV0HVUgDP33StoIZ9J7UkBbw0mCL7BKLX07LNNAi3Y7iU48a2zPfOKv8rX0ToWBjy
XG2Z/wVHdS5FUCnhj5xGXqB6Xg+1N1yD8sOWlLKv2aMNB6T+G3hk6eespc7y8QEX2EyX1Lct5llA
cXhz2/StesB6zh097SzvP1miDJvOM19Z2wZ1cjaP5iHHOkNM66Bh9tdIyYGNw0PMYz6pEW4OD+qk
IUv6vFsgW7pMOshh5pNvD5NSsbxxL+tdnQsY+6pPavN2wOCG9+053oM16hSXx6SHXf2hbWyL3OWy
G5f8et+RNr4QLwAzGChUj9iENV80pvIJ1h3Rf5lSSTKOU4gPoIzu/8MOTAerfrZ9Gw4+xaUm5NFE
M3DTG2AV7It7QcKmlb5P8Qsh5aziTdrZbEMPmosapAlTrnywi9U1op9lO6AoWi6GMMYIbK8K1qFH
5YuPqITUyn18e2cg0G1D37OuTgBIcR22Ijwv5TGS1pXFtBCVqrWLqeLYlt+EyyvGPei6bEw5pEPe
eZyS8F0BnR15qiBy0EDoutrMScL9rML7Y82YXR+u4JVWe33mxp8aIvCifGddwdkUiZGQGZGVREUU
27dGeEQUDsiOSvEnpws9MtWhxQIUuUTirAB9JjER6t+16n1aK2aW8Gez69v52dug1PMS+p0jdKpj
OJgwn5HfqHhsqvHrsBHpoWW7pPlBoTyIemMrywW+MRcC+p+ghB2gS4roQa0OJFaMC6ldBg/3sPjA
/WezRTr8baqOs8JpeITfssT8HX9dDadZCIGPPgDPkYT96OFZPlTwLKqZFgoeeAhVE9KwgRh2Fs/C
rbUZQO7X57cQ3j8SemmDX/k5KdhhdqJij2gqsvLemfE8JbMBN4MYTQwoZJgtHCzEOiD9f3Rjbpxh
AKYY5h5+c0WMe60mR4GJhXgA7LnC0Sx1Y4wiAVZ+JPmQx7l2/+6NQPHVDZYJ7A1LC2JJwkIu3ZbT
C4NwZuWjMXYWJVNqFAcqL516woWG3mpGpukJGOqTje5OAidZNHpbxPBYKjjfUnQ0dGD7E6Z8aa8P
7ZoQkGs4l+yCD46/GKrC0EjyJb5mhO1Xra0JhVo3HjwkL0dSlF/cLaakFB5Tqe0moweZbLA++8n6
SsJxPtdN2ZiWF2PUqEBnWwhcFraK7NsuTtOco2nmGiW+AghczVFaDE+Tz33QK7vapbBpdd//RB+8
zgWLiNKJklsXDf1HUF8g1tU7o87sj96xMAN6zD+B9n3g/HIN+cN4Ik8elsShdAgrjLSYxf9lu/2V
ObVsGVrzO6UY9igE9VPxEYEkb/gKIYgMwlBOciUE6yvoUZ4FycykHqyhmCZutZp0UQsjdgLnqC/5
pHkGKa2RXjsWDMgwL35lotHfvPCOe9V2loFpUuIG7zCWq3BMHommAvQDkWDGA7S2b1ICyZJa3KyC
TsDPbZfw59kPz8QtWkkUjSQzwPfsIBFim62laHppXdmpeEdiUCX1r1YZGTIPHy4+Fxzkw03N7WFp
RaNz4FUN3mokJtcAhYvpQZnxQANZYvpFUmonc0drSj9cRH1EOI7aYECyS9LivDoQT0H0SSH5fVRX
Tn91WL1WMpt7rA7MYIYpA1Tk1VQPEUfE/74gSPguAqpSnUzQckxqp4XX8WZWRQyxwSvFup8N2tJo
z6+Q/YN8nJ2FGLedO3msodNZhoQhmAx69juOggGEfXUbWrtZ54KwTdT0WXMFhO637fJuq8kSlX85
ltGmY/ji5aRg+jjfRhJg7qjQclVLuWzwLGXdUoImXuJAhslE8NcEbqeGVJAKC1nJ/qZAYIq5J1JL
lbne7u64aa19ncyjNpCgNxExzMONXCZVfuQBTflVpHjlySmEE9KaFQC46Kd/xMzdfLIZenZIYX2G
MoRXyeIMyVaVamjyTfmhpjk91d5Vu1JCusbT0UM8mF86ZNwuZQo8g3XCQNRRerSvCOexGrdJqFV8
tL8NTmKDiZk/Aum6Ert1Oa5icNhL2u/mTihmamNzD7yuhbXwq9XnZCIxI+DtA8qYWEI3rFuW/sDU
Ucg6Z6M5gQP5eGpoMtoiOQjlfNjl1Ykm3ltm2aLTOqII3EgXFPU4ep2gJ5reFBlj1383YWDIbst/
PJHSD2dv6sK9pmi6tUG2VOLBCrcuXiavJXar37Zt+2osJ4SA6cZmqPeW6JdeyR2QAWuKeXMII8pu
gViPJ9CfFVJVoToPavP+7VhJ2ERYIE6/pRi65Tg2OyOOiZTWQiFTevM7tbjxmBZCPyKkIr9CwltS
pDlhUGJsvEo/zMIEDcKCQcUDHeVCbDOv1qjfJearLJLtBTh9OmbF7la20xHjA50HuVH6iRGbP9jN
RijfcjhhQD1c4k6kRPD3cWKTqddwvhir1HjAMOJ8XV6pi1Yjje/J17ljoK/fOuhzd/8O1ROXtMCA
6U7xAx9z/FsTv6Zfwq2vWFcUx0uJ/lKmzsNAIGvvA07nGcyVo74IYHp6XZI5SUbpZuZ7DWn3L/3J
Ex9PUwfLFjhQEFRBDNyjL3LOM0M7o5PBR7+8J8k0pPhzSXc14lM4RGcUBDzOgr9dB3ytxbYZxjwZ
vlt+gUn7O0JD818JHjMEBX4a2U0RsfaHrIi9n+OYHkykgWMSwABNM+1umfPxgyBxlRLfI648CqOZ
t4g4I4r5TaxN+vDEh8uCfesIWHTkMQJt1dXyRK/ILSr01qyszZRsv1dyGtyyKHKTYW0V9Tdu2cZR
cbtzR9p+8BhU8a8hGO1m5ZTy08kpy2PNiJIbHiQfozgCAaLpauuwygDJGReQtx3jmpGdNOKqXnT3
9Kx4KI/IbRcH2G5QUiEYGXLidSrqazRzr6URpwJkcelq7MTevwXeXVvRUFJXQBACebtlEngVrmjY
nI+uMkn4Z6bApVLAGBY86+JV+9AnbDCNifIom2VeX16v4pHO6Z8crbLBuqxlMAQYpord3XT1k6Ao
frAvF3jxESdlfXzWpygvF8jbcV/xA+K7IJ5ZFEGWhS7o2hmmLt0kIBOuhgf62EifY3DNPHdJqlSB
4jZgRW9Wh09jZWPBPlRC/90ZvdEHCnyYlBmfabaQKtsRUBEyE7A4roo/86pW44KvrlfS3bpR0kot
gHZOhTwu15EXipfotwk2Juno1v1geCp0ZFdvEepJHOHENXhF4d0lY2k2JlbsBcGxR9jvzAiSAZT7
4kqnnwDCsM93orxYgxJ/b6DTweViZzL/Da5Cj4w9F/Qzc/lYCDJOvd5EjZtb9w37dHZLHPIa/15b
/enTmxBAlhujpl9aAvWPzod1V3Cr+ksTosAQUxvH0jTL8JpxsI/83vR2c1lk9eXqV1sn3W6iL8ST
y4EMQNhntk7i0KbG3S0U2m1y9ozI5EGSbZTFMsyUyMDTad4nks1/BFa2eOr2D+NWYBs4CTXUlUeL
0+dGSj1gSBOjxi36Dz8+FIW6Kgi3L0ch2/Sy1MpHb2psiCP+Z6sJMiMt8MWhTgrqG6i6vxec70p0
RtpCz+1gHI0DgCCSuCNBV11UwDQLFGROt+5/+9HZqD8Nvos/PMSdjjaLPWISlxSSnLARptzBKIJC
mwixozfo6AP8ckjlriJMXk589YoJoTnM6MiBlLS5E0Jxq6oHbL9aBF94yzU7SdSPHmOcjP3DuPkB
Y455G93D+HV12osLTtJS+oRTim4D4xlBeSp55JHHWHkJXIeZkpd3oO6+PzedvBujcQtYs1y5RK5Y
xxBrkKrHuQrmdYjrGXnIZ8B5j8HrwAqON0xdfnE3geJWjEDCu0qDLmHmVyK+7bG9nM4IJUVkhonY
1kSfZZkjekybA19fPUHB5qqj9T9xHzHE1dAcqaXOwuydsHs2I4dZlctYcZDIAkDTTPMTaL4G0E5B
3xtAw1toGPO9cEbfn4puvp9/NImgOPdeg1m+xqGvBRE9hJ/EzpwEpqeI6x0STWauSEHmknXMzYrM
uHe6pD8joIdWj+RoICtDtpEWrXadq+zJMWaMRB4y9iHpJG5yun/xQJrUF7RaKi4lKUJr8RxO5l9Z
U+FTNT7Wv1L6RnWN0f+HrMz2150vGUZfxFEKXP2Fowp0AlGpEDBUZ88RHfN50vNrqLhCzzdMMzaJ
RnkZzdfQp7trx4QdIsAgFokE275qI2XCKhm+yV3B80mkbXCbidGpGVBk1UZjJ52794oXd077vzOX
alptg1rATyF/EKuYArX9xeddBV2TwRbYzcG9IoSddsHDzSP+/KBVRImJ90quZIvaTPFFx0qcc23X
fylaXVxn/UYGVo2ehCPxbJI82GQO9TX2SlSv7Myz3lcra9bYftNpeZjlnQFrMVS3x+4BtBrz5+4K
xI+wdCBcHLNjqPytZYooUtty8eT5g3xk8oU5O8PMJYG+ZvpbwFud/psIq0TpyS1DUlJJPVd24PqX
y1oiywGDN11AIrNMWmS04oCqN7/6FHih/28bLSU+zBvkYATVn2sVa0dzozrCW23/TPg2T8oV4B2e
GlXhW4ulmxGb4UaB5rp0nQNQ9fsE2aBaY1HUAllDXDsAWsmD2FO1LMJmHCC3gITo92yt7RUD6Flk
c5z4KkJxTfO0J0TLGwDffUKxWtVtwkfRqso/hX0P4dG0ZbXGzW1Ly0tSnkLYlnfwaQP8+sk27ZCD
k8/h7gyuylon4WVeAUoK42+B8kA45Ojk/Ggwc7f8TiLQXJpBfQGqrHMdZWHKTODBnXZtbFWN4XuQ
EzhfKVrdn1EKgcpAQ6ulkr1sgkHCLmDLb15Ahx+wvw0hcQNJLHN/XLlYL7FISqRrsQzzg3kgRhPU
TVh2syhwYhokF7wm7FmVOSRcLayuSbEm9uFR45wSXld0VpmQj7+6yGX/Lpez8iuZlj74u8mdVZxk
DPFsvwEn1R3DKilDqQQ3d4YTDDBPfSyhDntFjgIlsPUDd2m3HuAZBBZ2njYPg5vDJoZ0cTC7RKx7
OBXRGqdHBQpGVwN5cNQiYDBrf1woAV8FVwJCwwXcW8bGmcgg5VR271jTXr4uzikvrERtaaywCVBe
hSkSe8HWNYWiGgokyKyLMwJJJDrwFhDrY3RyiR30N7IF2okhHXwcfLMWiwea4uZkduq+xYU5Jm46
wkXRK+/1vTLWm3YDdr2mn69WW52Nvj9R66IHo166Z/HorgUtAUsEr4bhzB4YrclNJCd9TIY7WUaE
IGrQnRKSfEhyZnt2KrABAmKiuIMJnS9B+gU4EtDvvxcqsoOdloA2AZ10gXT99ZPr4PDafQK2coI3
+1l3z8xlPYIvhI00qPmGrBDyxCI9f6WVzwq0FwfaXTnP504NR2ML+3siDFZrk3GYYHK8jvxIhrkM
MRB0ArWgUDabkFSjiluF/UUBT31gryrBVavBUpQxLU22zH4/yBj+JS2txZ9ET4s8ogIzGpehqE2x
xGmiF4DMPnaeZYT9z+OUOqOK+kgSIvKTjJjxgUG3A+PCB6rrD+8L2ZfgpkoO4c9hipeoAYpNh+Hr
q+NDhoOlZJyVhJ5IHPY83Z3/JrtbPTn08EfuBJAy0AYMgpNxM6LcOJLthbkQjOQ/HzZ6LwTbHuo5
MQicuMjiY9qUGD0KhR46W8nNGbGC6KUqOi5oxZ0FbuIGaNTUHMimd6LAyFeTNxoTp/x6t27BdKna
ehG1ELL36ojjqSmuNbbmolCtuB5vHGjIXWGmXT06vUyA7plwW+pBinwjmUxAlxETGT62zts5scgC
4SgLO7x6Hq0g/MGmW0o4FahkLXkfDbLZkpzehd+sAG/MjTvEKCI4/AQ/7NTv+qcmyANxu1+fzjvU
pzef24M2OpNHr23Rmee2eVPF0lGEvZE5VQY3fSqoO0Mro48XwHYZZVHtJ+sSSXQApVmAq8xrCMhP
E2vl0EjVIOK1uZO6OixgsWYssVYDMDq8hM3J+BEC7rRU8U68FMbGoqlsuJ3DXDSsNEgMZ5CTmPEp
ypcCwOZyvyrBxFpWeWvUbFCeuM0KKHPa13sKyZyhfuUfw0SlG5qXTryf5Pv/ANfvpVQmCE2AyRyt
lD3zV1/UlaCh/mvmvxSYHCTpbx1Ppe6K0TwECT1J+xdKNGu2NbFEw7H1P3bO2bXAAaeCHd1M1ikg
+ITeGPWQx1gHJMCCezHeBt747Kt5pei2tVszc3oyZ9DqX5HzqEZwRF+pCJI4ntIgzZzIKZ40R7A1
o3kS0e4Yplfn0rrAroOKFvS+Wns5Q6KP6Wr2HT61VCZnARXyTQi4zenpSHO5Ed6B4x5v2Ph3t5y/
fRvd8FSd4RKFEZqPHVv9DAnlnE/SIKSkKeGjibQ280ZKTKjWQVrxzBOFh0atT3phh6/d7oRjt+U8
5BgU32JaX38FV3GMrO2Jfio7KjcKmO8RVB2yrfOYaMKQdcGbktZ7fdRQNP2Ju2VrxakimKqNKzqP
MI2nEIJOs4FbsIHuUaXhsomUF1fPud2ZJ+GZPcoGPkGmknhWVL52F6NJixMWAeYDP9talrRvCZdX
e3YrXPMZhZL1e7bnFgt6VV2NFO827yxcPqOGGy28IgE2rgKS7VePrxK9RFfu96p4m8ZqwHs10dbw
5IWfos+JFnyuYrNRKCzj/LPNNWTRQ5XkXZ5RR6KgZdDYeOWIf2WryWg81zADOYjHwci0KtQoopbW
lD2IBsjVzj3pDtDv3EEOaIJWmaCtXPc5aMpzEi5roZ/1x6U+shd1OfvsA1dsikiUupmyaYHUO87z
qypSOHhhefbBpcYsR+vxgy37NBA5bpVbrWl5wURWMxvXvaZab+q8eP4ZivTxFCKuq19P4EW8t630
Ns/xG75mGxBfIiJf5+5egyHS1MC2p5Ui3BTeAXQ6dz4X8tRC4w5Xoo76ExlR1Egvxpvlx85/e0lj
pRcyTY1Q/F6mt+V7KpMG0SgzkBmfY2/B2e1Aod9kYIItyPig6tVSLJ+6vuIWMQwWBlX7vY/VvK9U
/PEQ2N9mKqDglrB6hK4D3bCJH6Ade1EUVcGoUM+iqn4tdS4TYCVEnqTw1v5bk4RTvHPrwM2suWDv
KbhP4zq53DhJuYhgqhVhIUqdE9dJQhyDfHn+RJWi3cC5INhy1zs0odmw4MOlB5E+6jNgP7E4f6tu
Uh2pDoyCKVMC8eoAwz+QvHPvZ1s+2T1DXNmxJhmZ/cP90F/qs2XOHcGgrsbJPoYhcXKini0aSIZt
LuduoqVoNLp3he6Qekn3gxFk6A0e3O5phowmIPUA6LyVK0snsiCmgyufR2laQu3PcRs5r9QZljLh
Nzn5K93/V106KkPuViO+dFsodtjCsId2GKBA1jpFchJuafrU6C3GxgWxbzDmLsI5aT4fAuD6u3uP
9iOHwIh/F6i12pmFVTn3ufAlaXXLtUnOzco7oQ/G3JTI6fEElwvEOkHqVhU96NqbV0PuMTbQXCEB
4OItWkEcX2XiuCMEYB+ZjGPSBgvgYp03WhjAl3nR41aNRmurK7HgvPinWEpNn8ymYbUSdunPNjba
omEt7l53YYxiU1wpjCAlyd9OBML4DCHfJs7jiRnR/kf77pwbkEPtq4JpsT+NeSKOtW0tSTnL7HFg
RUNp6+3fyGQ0XzEB3TKfuBl5ssRK+JD3GGHsYd3jmdkV1N8jdGeHJQq0DQSX3vvuMFmwtY4/In/D
H7RKNNxJqN9Acf3O5+w3E6arkkJkXYj9z9+yLf8KAqxkYF772fF8ktsjd5CkpkBsMAE/y7UZcoik
sW4IE7sdr54iX5s15nU2DkDhW2yi8EsxOsKqfN4c1flWo2jnfTyV6cV9z9R/hIvy4YK9VganVQMj
hBgUiSVVcD8NxspKUVzdwqxbwd7gSWc/SUkm940H0taY3p9JLD64H/EhjrShEw0412qPYin0xBFv
4YF88m45R9G+wrI3Jad0Yhx8qjtX6bXwZ6A1F8lVSSVNRJNOYFnIpigQ0YUrAO4UUON26Z8IoLLI
/NMYILBTPbIKt8ZlqHAdiaFlzTmLjGr2FY3KWIz8HTGa+axXKmPcKFgyVdi9BqtRhUTMKd6Knuzk
GJKjfy8+UGU8M7BTVchALJ+KotAq7aZNOneotKBDAX/lOx2oNTjFsOZ379z9G6rCtShvedRfevWX
dRLUCZnnPsSiYfWYm+aDjtIHrcrvJKQUVNugHwnOPmWp7GkomHrsmeSyBJBVDnP4h9kaKkTd5Cna
hob/NGUvZ25f9/CyyIs5B9FBTVMIE0dxXrjH92ppUMylcT29MQnAOdCmMY4qDr9Nmpk/4GV4EsKB
dCnrGtuaTV6bMEH0XAyieVYb8yJOKAmankv1SHjRGQWG0gwuJNdRu20WQP+uSPa0ryJDw6cPVf+Y
Vn2gpfg/h9rNDDoN7lp3owRSRz+DYyNLh/I1Jjcg+SVzc7o+lwyTi4j5UETPrRaHu9xhhjlN1Hhp
mPmi9o+CZuE2DNcY4ZHx87zmrGp3AxHBNXMFdlzcF9B5BNXBdUhfEf2liNtrSkeZpucXrOwnCGYh
ja5pBX9nASFoqmOkGZyaEHarGxFsfg0Nn50W55qt1XB2M9LTfuOxMAlt8zH6ooQl3LeUWSFV6q/e
oMugU3hEHkg/zY9KXFjJmPOCXY7Llm7jcfjd4aQ7bLCZFHWZ8TyZ2NLb6P+AXyPTBnGw6H7UZtQX
5bSSpR193HzX9OPbcgicNSeO6fkw4pxsMfg3rWw0vcFcB8Sterxi1lxlO7BbDYl7k6LJ6dG+f0Aa
gtEjR82prR7tnTfLCvp9thjpDHXYV8hdrASKKhyyzK5aHqMIpp+O3sU9K6z2JUHLju28EsKaisto
Uu066X0Zu31y0BbJzI1TbsvHVJJR+fqmagNdl+7hDf9hHYSCIWTMj7vk/vNWLx2HabxXChsB2RX5
oJZ1VqwlO9LGcDbk0DSZcze2vJwrQasJxfX9aDSB8yZQL9c6uKUeLBKHTXswuW/14tFOVFZk+2YI
YwbUVGB9R19meK61LB/WhTErYqx9ROANscYpDLkMe6vEq19ZHE5ISKjgk0feioCjPDFe4jCtw6Yd
7QcQiT9HLxxynDBBr71AdJL5zn2Ko2qVe9qpLV8poGNwBeEzLHg7efNbXcEU5d+Piayx58jjbpxO
9q6EBOuSYMj3FR+qn1qiiVuqIAaErjddU4mHG9hCmmz14cT2WA/h4H6GM47n3YkoQwQ7M8FjQHYN
LvbPXoYksUA8nygAUHZQwGCezhlyEvdAfpOanW9iDghaxk0xL/N5piyUP/C+6iSRlT5YiIb0JlX6
gu1strQWcIX+nZDsZ4815ZuCmJWo1LYWqQa2GTPf6Ro63+eW8lNI8UgIB0bUlsMtgyeodXDNFHP5
cURTXL0XG0qTyhWwRoBCYUFUV6chfvlzXp3yB6TFgbvQ15XdLKBTb3GYVNz87qbhdpC0RkBzqHhm
lv2MtcIqN8Y8nlP17O/miCrO0xn3K1QvqeAo4p1QmM9PMfkQancU7THhqr/XsnNbwz/5RLtWIUTY
I55kAkD3cdhGH9RodOjZ9kEHkYqZM5emJ8VDxJiw+MXjTqZ4aXVOuoXfbboJiVUCvK9OWtpGOve+
iC1rJ/T8N/KgkDYtdw5EQaVisPI1wauMyGKHLj8fPc/xAcSjrNjwW0BTa05Z2leTtClLORUaaS8s
i+Cfx30aQZwyNyHyEQlJU0m5E5GyytjV4sjTzKKAw28P6Yi2wO5/ya+jANbRciX1lWzldm1f5aFV
4I8sOEzxFZD+0akHUOl0D/O3/ntnwSLBbXeBsrNpmHgNh5mSUqb5atfztD2cPVN2MBbU8AEN/qjZ
cn7V4d4SJL25VRLpKGXu955C39K57Yp7SQs7t0jMSRZwD5NVcWhxfjT6tdE83MVX8Smf4SgRYgA8
tFhcnkcNfGoPp4paHzPxN2CNcGBNZ0xoffPrC36S6E+IZErUIuP1MUbTkVgBgHIyxo8CniBjR1ay
buicBOOHe15hPYYMU7yB21uG6tnR+RZTw2pk8lKeofA5qFR8+mS+sZduerqAQvRAEIiVb5A8KeJ2
NXjBF03AlPOfMWpNRC528xAiJqhFtdLuy2fHFQoc4QwpG3gAxmX56owjBnNVlO3KPBPJNUF0kS9Z
HSZIgmGA2aXrrfz5ou0lPSlQ/WmpQ4+b/fwDYmvC9CLLDWM1MMD5zQoPPoJalMhB8HZOzKVtVObF
7HFMy76KAx6ipUnGyoHUmFB87P95Ili/0wwQcjoEMVfn18L0sBZS48ED1td/qwhuCsmlsBKAedAf
M1PUq3WTqO8ZlTUu9wODsoIFlr0P/FHx78Y8FmlObqVDCJHuJmzCseTmE+a6A2GIIjC2qwxmiP4c
SJ/bI5Z7zeounvqyTSMPivn8f/9zCJqeQ7joqqc1Nj+v83tk4BN31WdvojL3tDzRcCGGHFlePS+g
VJ2LMWFfAZf/SF7xnW1hFZ+m9etg8olNAwo2AXZyQ7fVDThdFXykgAUvrKFmyOKwe10xgtLlioN4
OcNt6CDNnnOAuVQJQ5ChnZ0DHESWX4GwA3a/QVkfxlHemtAcYivuRVr3ih7lrOk16vQ2UuLZvtV7
Q65Zk/+dcJq/N88YKW3uXlgbhbmo8TffsEfaMt+ZmuJj+C5acr0t744Q5PupyUeRYzm225ad/QWE
tUeMLLW4Tca2dnhhaimUA0DMymzfuvJhByzzC8DZIBPpqrOL5lp3sa4ybr/iyls11BhZNI+T0rjN
OgqD+kD3JKn0Ovg4bcBTA2tWVberNqV3KY0GJGAU8Nj7g9dfKogzvZUgkeARMbjn9i6KSLVDiDh/
Hc2IBMglShXDHNP4UYthKobKyRdmgyKwZPmhMYluHffdw8c/SxnFjAJZn9asd7A+sgPtIFi7yIxc
7agyaEl5cf9EKAehV1PXMItaNhynhappfYy/k78c6DYO9iRatqgG7e7v9nGmTpCWDJKkBJQCF7la
YD0+V0oX8IrCBXE6nrlUcblngM/UMxvBxUYv2GIkocK/vikJXBzR9JQ/iKtL6CiVYwLBTuqUlNnV
JJ0+9hVj4tc3R8ZeeHPndP+sFhXsRZEpQ4ZAUggmGWvDzINy+0xbhZNWVSRjsJafy/qHk6BtSqxs
sIsSRhqSMlqVZu0KzML2BUK9Hf8M5TqvXvq8Sa6pGUAKLjbP+urzCSsAQlx1gSh3JLojInct9x87
7ZHbktpPqAY0VG2beX4UfZgy4y2BvTUznmuSqx98dUTu2w9JSU1+o/n9zsUXHBrIbnsGIe9XL6Zp
TH4tjWKgzqLuLg5WKlyngBTfqOwRB5qaFyDwEPtY43BPZYsYwEeHohROpbbsH1W0nuuucodu04Av
YpSX2TTJ0gLRth9fhbinbbmH7/ORStB+AbpsYLaXtCKH7QH7DGOpHIaNvtnyRKSWXxx+LKBl3Fuk
XMlQzdV8D+OvQus5gREGqw15urysLA8lwNyxmsjHeBEMtF3+p/l4BG3OHiaYX8PwMngFXW99YJ5e
L4T1ChJSg74wxg6CR48PuJTRt5QNZ8ktcchc0uI1XfBcem21PV8WOFAu2vSscT4PxIaLMH9ZslaQ
5CgEGh/I1ShB2nuW0Nsc/DOpl5BOysVhAHLf6yaq72I1OfsNsCnnrKRL1U0CkQpK+ObSb/NjMGKk
pOXZXx9J1qf4qJS/Gt/CIQOqfn0P96Y260fg4T5oBhVNRbSblHnIqKb1/hNzQwwHYZM5gHRchbu4
MdlWKweAMRlVSdrmphIea6F1A5ag36tp4h6En8f8AZiI1ixsc9a64cQ2kzVOCx/3CIbGE7WtlAzD
YoVPcpj85sS9LliuskYwcNjuADWJizssq0FlkMmx4lfKuSrxfwp+YrKnY/9b7dpgNCRd0ivbjcY1
w31xR52bhc9kssVbvNrQyPBh0bQFurREToksCNLa2T7rVRdbzX6Vkzl0Jo14oWB9l7BDk0zVapvC
94TeIpvA7uvvCx/k2iXvfwXA19yRKPC+fAxqqU1ZcqcidRPI3CT4Tln5/gc3dYbvsBbUs7RLFPb0
aktCItrphceWIxaQk5Ih6yvgPIJQOA3WKFL7Ai8jcPsgFCAYiNcOM3gpRDrFn0Pi09hAzIfLJZ4J
xtlKLZvis8zUIG3Y1+pkyTDJ0t+y53JIm+AbFEKxSOGFTtlqX0luLnvUWdwuIOHrrFCDHdl8njRq
PVLFD7Dg8tYoUE5crSE/EY0XTAjlkgjEsMhnXTx/9pIov6nCJDLhJ+7MBszrJA/G1aiRl8+V3rPi
W/5y/UVit5uLjx6uVBbrC9wI0tanKpT467PRflGZK7L7UxHSTFZFnQ+XXKTAAw0XMEFS65o/W0Sy
gnbhHWEkeMd2XdcvBgNQaLLX1vppoJw4mPRpYvc2VZdELSKWagPp51rRAlJH6cYstzGlYfXDSjPK
eqqsb7pJ3tCoTw7jJHM1tdT4TJccic6225cHXAVwha6BEYMGMbNp2I6rLq48uuY9D1TZqq3H7LQg
62I9VdSD36eGR5N42jRj/vQghHIFiUF3ppKXs3MadBDMMPTqLD1IOKTOJb5Ji6t1cKxJqBKfGpd6
A58xheN/1WrpToNUV1AX5ih+KidsD0e/RIwj48ilUlL5hn+TyagvsX9x5qFBB1Y05QriLhfBtBUR
8jTgUHfgNiBv4hctFlWRtFDQA0p9io+jsxZ05wsVZc8pOTtQ701OK9Evipa30YmbyepNYjG3TMhp
XJ+wJUqtU9l/K+Np4eRwLdBC51zirKtATrhhk9qiuUimoLA2ZzfAQilhE2d1gid6AW9NgEhtHP89
vtEU4LP7wxzX8LypoWtLnW2s+tzjGmfaB3cDXoNziXjQeSrN0KagTV9DDrjF8S3K395jT6FPuqpd
/6liyQdQYKKqKLn02IPI4AwA8fiHMGJWGnQ85C3OUEXk7fBSMfueo0JM0mqE6ZhthcIWnUp22BU1
RTXLb7n9c0ii/R8zyAmVm3xEdPj5C9YXXs7SvcYUykktSZiMxT4cVvwFht0JZ6/SrGZkNJUx2skZ
Hy05+uDqnO9VnLHfBIboUGLIg9N5PoBU8/P0ujeLLDMHmkRrGTacwOXPO1av3vr0OXmEzBinSDT8
bwm+R3DyuIsHGlZ0OejDZnpeDKi/tX5TQQ0kSDMQ5V82t9AOENT3P3JTFPUZfZaUJmu/yYQY2t8y
4FswY/HbAqBzYNWNP+MjLKyiDesO4lv7qF68LJNS9QJCCMfu7nT/dG0RLU4teqTTiGqSbHYOaHj/
hovAHoldm4tMWRrBshbOkQsUBDqY+L/YqPwA9D9U32EYL3GLGIUM0eC9mrEna0t077WeUe2+zdR0
3d4j2J58QQqlsXibtHWpabyWuXsS9CthSIADVFM8mjZ2BD6gyzJ6XLHbUOvfTiMcFU5cc42qutLc
mhH+h/VPlu3wyVcxkHSl5zVQTMfoRGI9w7X/I9W0TwKlWu9OwyJuzDhsH5NH3U6spsA6takMXEhp
qP8OkNI7porl2tkN6RgQ5MkW9UOUe4gkTRWQdVF08D/UrQkWXmV+pcs6MsXQL3mJ9ty+3oFp1848
E/fwLFY3bGZZ02oeseJh2KYN3g7rbYwFHwTDcijY58JvoaBmMQKXDQCU+HqsTbc8HrfsRGdMknvi
Kcz4I0mRQDv8FoR1lsabMs0mlk+YEiRLE8bw1780YlUIgW33XnQ9CtScUjltNZ4CuWFTc4ZzzEPM
Qxpe3h24B2R18zcWjPr0OPT0MIzj8wFSyBJQ/PIIe1/1d3XI1vbYxmGl6Nzlo09ZrYsgBW5fSJZ1
4FwnwT+4McwfC1cc/UYCGVCRzoq9H2lqCUxJpKjSFJ1KJPVcvjh2414JswnebLNNfRb1Lb+M1rYU
+GINK8T7XzNE2e83MIbpuwsZ03BjUnaVcUtJt1my8cR/VIkQNeS+C14S5rum+5fUUH0HfN479wnt
oeNoB0Aw0aajrt91DMqdaZp0XcHNyqQNnlvGMFuxigRvOjCBE099nIL0u06XTlEPJeW0j2zts0hg
MR4xM5c+ZvVgTkXV6b0zwK68WmFrlDXgub5gG3F1mGEePVXUQYBdzkJGHxLoNIQcZ0VxvEDebMH7
GeS3ZSbOvzKhhK1hIYFAi9U0/VRAi20fc89XxH0jF68gFYkvMqQIwR5GojCPMl3oFzVoPT2iAUtA
UMSnfP2j0CKTLwXPt/JjnSIsOU/ldwd00XRPkldEw9XXh3yybF7EIkJR3KltfpV4NUycUJYSZ6Bq
6/LAlat1NwqdShFMQhOB9oE7Oz79duJhnpwk6Q8uVqIMmhIo1/LP/wIu7CdcEMuCNwE8SQjOKWk8
4uu0aMyU9Gj30JWELR+HPhGnO1i2s5GQCTfDH6qtAp8KdmVOFN3jh9HQWtghC55gfrJnjAc4O5rU
55SgDsbMZaZx1iZpCKsJSvxwNkKnDPk+Zxgh9jLHH4IuwuSk2jKmqw6FbV+U66e1s4NoPFX0dPmB
IKhpBF1cWq+T7IpFS9URBmqjRhhdAaUq11WKIylHqK/zdZEKGYw2/yr5sDJSwf9B8Ao3JFtdBbir
WUVB7w7tsdvbXunHqFSJIxfgJpUoSY2jzCdEncRMcWe9/uHPwBYag2+EyaimxgomKFjhsHwZTnLq
7Ufr5djv11kKm32SvL7kelUrF8cRbXnAxlYE/nv3RB+VoRehsO2YKFng8b+mDvYvrh+43KrgA5F6
mZbdiXytN+GIOcpdeHYZpaDIytftThi4cHN+itoSE+EP5ZnHXoAEZmXec2xEhVnwqitWAsIn1hlk
OIcjU2eQoQ7/yGDQkHc9KwDBjrEFH75PBK/KdOblqOoStgbspL3I1bTSoA6ptw4CCQ3MdSDQ12Hu
rTFS4R1dDjzuN6j9gMdRdm+Nv8+zVAtc5Hrz0FsnC6ZQekJMaMYxfAkJULECjM0fWnIJHrKsrf6e
cLeUVbQQvxNi1CkuP0k4Fqghipwn0WzzqWvm5Ul57/Vog989KI92dY3bbIiraKe7H6XcH4Qzfykp
ploa/9Msvg0rLdGC4O3tWGJL1wXPn1eyKjAUIEA3e7UgFO2dovayF145CaXJ7SYirdInsU+8fI3g
AV0F8/eEHVQWMTZdxwWUcUNYiP0N9h3X0oEvlyP5T9lbVFhBYZnPXJ6ds0EzZRSth6aNcisgIlQF
ReFxszIa6uMbO4SnmniMBBFiAxSGR8asmD2y9n3bUzvP2oNe5e1ZsjDaxEx256oDHi0bxZUe6Lbz
OlY0ftWIhFhpcmDzQElVPqGfyMMHh8tIQCMIH1SO51Xv31dZT4ceryvIo0BmakB6lNAWmWPqJ6ii
dLHCQDpE2KD3xqj3SPUMc0FaeaRhSJd9oEyw/IB/dLwaM8PMLGdaB0ALxosJTt1yAteEpApJMJMs
RPXvDrQU2kDYs7TFpmlo3Yhws9vC3Ksnw8wUT4tw6g/lIs+dPELyaTQRcTu0Alc5P4DIMqPus2Od
ZwQrqTO0f2k+rZPNBrj9DAkVNsyGrKRaS4e/niU/hbjyT1ITHmVHrawPqTM174dB6dTGYiqIRyVc
AhFruwtoVN9TA2jVy67cCMDMkTrLnSy4S6YN68lQygj3O+t7D2Wsa5Q3sjRTNDB1YcULgSd08q+o
QTjf0DUCsWMJOfR89FRlMjda4+HR88eS8QLEDnRrT8IKwQcy+aQz+gn7sSLd805AFjfMAtBW983j
xcvWsIu2s/gHQiqKsrW91vBltI5CRv6p8pXOyhlqQkSLbRFpl8l2ooMO8FGB7IpizSdML+g+2+JJ
/g/Ii57SuD5zOHGrJhStSFcsaFpSQeyIgJ87i2Ds225meKUyQLfDIv0qOImIEHFA4hDkzfldUyfj
sDfdhMbtBbu1RqArkbszvqrGjN76+gqgkB/A4IjjwX8TRTt38S8YMstQrAvSmZrAL/0oTvSSjyEE
w+A6BFe6ktkgA7Oyk+nT802tQDtXoI2cgkziy1PsDZNi9ghT4nYFG+yEwnWwFT0bZHHlmz/VyKRG
6JIVxo+7g/wDT/m/7CDDdJW7y1pFtxCZ3zzMXGot4HTs2oOBoXAcUYkQZF3LLBPB7k9HVxV+BenY
Kr4C/7FG46AU0Dh3iqrHdLdAyfahxFJxm+Rbz9a5UF8aWb8JWjDbTpH+qhlV03rTQBlj+8IH7yyA
m4xgcN2Yalf4w7aOvaHaIaL5g+02bOdsI0AGEFRG1wVTuYXs+TBIG1UqsqNdBfu0niOhugruja3q
zhuSefXWKkCGzideV1yGUhEEBCYbYZmfbj9pE2FeihjjhG15mjM6+sCpcUcM89wzfax72jPz23Og
rOixPz5fd/g7QvTsmaY/3YYPuK5DjEre5GBKeo7hcHcsnLzHDEyCG210NWWL+O3ZHNVrFO8mk3yg
WPATd1EuKgifvcYjzqPl4fAPZg0WscScWqJGyC9xmLf9xOX07E/iA0tmHgu8UEC1r1QyMnGtN7CV
2kc9opjzE64G3wKPqbADHNLdf6K48EsskcvE9FB0LLZHaZY9xXTr+WORvrpc/J1vnY9zL1emAGe9
UYm2VWB280aR/SDwL/Hz8g84z30DrsDmR4gN/IGa3JHySN7PIqD3r87350KY94Tu0Wv3Xk74tekZ
/wQrPW+XcdFxE/Q8V70OHKsKvNMjSa26lx2vI1NgDJDYXbtjkpyd1BXGcKCRhSOM/tlUN2srPA6+
CXGLW4WGT2ZpUUqBnztZab6CPixmLRk3QVB/p4q+2o4SYmjR1zAVaiNCX8lWmUF3nM/q8kMANBNr
Jz6dcKC8qbqTRo1j/B3sZFRGrxiGk71fh46/l3MjUFFHsDN5gUIq6lhkhiddBhLnGhh3NFXCSOV0
yt7YNmhpIi3A+GMckf44wIUVrOPGzye+rAHEOc6fZUgfXwl36Lsc4fVZEXXUCRIr5EBrly93PdpW
O0TIokGj95dbV+XMSOLa905Q/LdZlgUthPpT79dm8bKCbDk8cpiQeY3xJdsyBomMczfr7ik9fDxY
EMiwxcu8yMnRNUufsuzv6KJmP7syhLGC9gR1nZTZdCn0uJu5jP8USBlshHMutQzCW1Hsq/eIh/PC
Y1+Jaf85vnFCL5x9c2pdc24bX9NQIH+o5jXd0Bn9bAXXcadvRdWALLFwWidmbyrLQXxC29FLgALH
IeDI1ME34UaGHo+ywNp+ZU0Av5Dg4V0k9mu0JJGWMdIOnvvnnCROxIdAcqh7cmRNjLzHsyEjitgX
jClMmi52ysuZF8hZkgcjII1776qHCERgYelqEi+ZIs8dvuWRhJ/4uFDh3nUez8ZVqgEtm2D+ZXdH
6DWcnAaYl5sUhOFtR45NHEFDeP55nh8fAfStBvakWTEq+CGHvmmUcuE9Mwezl3uYyv3h+AXqvAhe
/oEd8T4Wr/n1CFAMM3dT5JnMMIhMCk3pKzwOPQJdGFYoHGB7SXXCv4IW5twlWjrdWimMHsaQBvxv
A6kWREVkHbs+ybnj6F3T5UxkUPiAbPNYkrUghbQDGacnH8k1bT4Hpm8Bvh6CeZQzdEOAT+hejxW+
c0bgUrmYi74kI9DxNbyrm5OSaXbNm9uxpykRcdl8KrJJ0LKU7MoqMxew37TPYUIgOg9CoVzPKVzP
7roYqb4egAiLJi19t5NUwmqerGrGr2ZH6Gdocy3xEX4HS0Jq9M9vbV8STrynYA20S4nJJ9xTQ4+j
qBBV4SlhGTVKIiBr1FKqJR69pHCjq20TBM02/ahHYVAv41uuyu4ckSFMc0PZxar4WTvM1nCJmxNp
tivODn3IEholJ+JUTiOKH8fKgq7t89fQGAwna3tsb+d/NI3CuADUxM8ZnToiwda6y/4d/oTyxklK
uTZ25NJ/t1Z4C17O86IosZiMafqwDyrIIzmyYqLq00yh1qPFD7z93f8lI6b2rNkH1KuF+sZK0SFY
ldrtkB7iMobCeSWrUC2Xv27rJXNvf1EfM9NL4BW5bXnDUF25rACavrO07YtSrcmKSVcte1a4xgJE
yVSHFb66ngnDBFKoJsk1QX2wcsUFUJ5qYa8f86d7jTnDzYeJFohJdZOLi+dKl2aBdPd7O0ourW4G
7UVpHsGOITASr/H2JZV2oPmP4mY1zbuA1hxZYtT1CjHtmn7s7kxcdxqr6mmSBDfI9O03I/Y3+jCc
vt23/ojmg0StEBLNjgtgRYRv3fgOsu8453EdRfaAVu61/ZqxIHbfbbPFV/jKAw4I6Va+XfB0MlYI
fNiqMZjduMQBEUyqzIArmxHSQ9nRy3AoiMLOFOGJ806L3f8N8y0K+DI0XQS5WqMYlFZcEiL3eOlo
V6tdtKj710237QeKXS4vO9pOKlj7WVbbkg0PZ7AujKRFs65cH4ht1sfBST5xFlAsZLe+7OxrEKly
t7HunqJi8VOuNRQRL7IXbAWYZeLiD9UpF69Ys8q6xPKeZHC8b5sBe9Xr9ENpX2rERR/ONhwJsjDR
La1Rl5g8YDcQPMGsiLFFKHd+uWAt2FV9ktpwp877T3iw/65nt4Hoc4PC2HDu/ozna8o+3SD7vlEd
F8VLDsj8BTkok1zFrYq7k7lA4hSdbs/eHQATXzDktJ1GVjY2w472Zwls71RRcLySBMUCSj2c/GMT
mN0Wo5jQJYxYcwHwBPmu4iY7RZnnHWKQet1NwF1xKVJKGL3HGOgAO9LX1V0acpPzyLzUXnwQBvvG
loj8X/JE2L6uWO4GlkTMv+QdecpGfkaOGybD4mozCL4eVVmSXisf3oaTA86ydLAozTXpf02C9e6P
wS8e3a3bzekSwa7vpNvNJAms+UAn3K4+uXUSFUvcyMbfZKAIwT966wxL0Uffg0sv4ebHQnhtFAHv
ZC1OQHvQ3sN8pKQZdAoPWNfEEhi+x9GQZXvJmv+WyaZ7+C3OmVCzFzUzpqJMKDG20mxfauqaegN3
5IxtLF77awqNT5i9/H/REGASB3iDjmyVZ1fe8SQdczkBwxOETTfne3KSiUqxPF57RNVgTkjGpStL
id+7U32VLO3AI9MiUZyd19XM4ik0lwN8HtCiUtubIOzlyDeONQkFaBORQhEMfMks5g4igrtICee7
0JJ/Kk2G6xkL61oi1izQQjSmfJQKGJSCdJYzQjBrzRJJ50FRiwr7/f3d+YVkMgsXPF1j6zlDIjBN
GQ8xQ/wlFF6M+kBQ1tdfkeQjQQ3zQB9Wpq6+gFphBNeTEpghXFhNp+CrzyoHZbfi5I6Ck3Kkh/1Y
XKStuI7zA/aQO0/O2JgMZ5GiHplemdwgV9OzZMb+WkGlrj4YGE/ViorWjBQkwc8v93/UEi/rhc45
ouHb7O6QT+iQrKvP/5HIy3rI35jqLX0GxYC7zwfaJEBSpTF+NTWoYQ5Iwk/WuZmneKRmxVU9KYqR
5oloaN5cr1ks10Qyq2w0gjfOJD6/pHr8o3F9FIziR5MPiQB8p0y7NK5cr8WwiZZ0PBz3CCDBwR1F
88qNylOSi3Ar6g7zr14UVd4qnzJyNEb/QWVAoLhcHvbqhX5tw8iBzzHLvypB0UdEPQBcB4O6zhOL
LRqpo8LpwH8ONWAOeoEOJlDsXXczP5y9m1rAX0jT1Mo0ltojGXkPLGIu8UKUyuUAnZcUsc3N6RdK
iltwwFe5VFuyzmtNXLtyVR2r1eljZypQ+mzBX2P5zi5ptpyh5xqB47JbPYdB48vzzNwXNLXi06dW
0ojXZb7u8FEMyBfB4cbknr0LgmObbmp4EKJty03O7EpyOynxK6mBbImv7Gvkoo6mZOYBW14UKOCP
a/vcxV+0oMggZPsMReLVdvTIX+O0IJr5klXuDA8omD0Bp0+fnOcEDKBd7LwHmPc4jk/FZ0Asvjae
gd2clfixl4gkgz3/qZDMGez48dbR7NT/ny5opdncSjrpqRyOHtK+Tvk/kkTgo7VrvPVNAUmpYGJr
Tr073RBBIkOMMWBqnkGa7MKeRIip52jgylInYLzYBuy6+4zRWlXNbmp+eq2vwUQtOGixmo2GH7z3
DDq5gUct+pdlPP6WF7nVKq56fywhJMCpfnwb8n2CdXS9xUcUm6rqRzkq119VKPhvm2Xqpwkh/yQl
GQ8WuRZ/DXwk+3wGHdL6EBdlgevW+KMystQhJ8tEUxA8uInlnsCLIYa7Y5yjoYfRDmAtfJrQB3Bs
ugAQ/JST+5Ma3DjGW0H9bXnHElxKrbxhOoQIA86raylv56Svw3Log/t+izAlJotmZjrY/VVvdvY0
aWhQx2Ze13krLOXIs49fIXdvL5xuz2fUb9fdBzJOTRgxp/fi8bdt7rgu5/y4MrLGvMeUHbgs5jrd
XO6niczQyJbRgh0peH6wATQknjJxnIqgjqnnRTERhJBeS/aX9YuCF4+0FwRdXYhuUDebKLshzIrI
J69fJxL1dHiuGd7gtgXDRXIKFZ08tkGASwKF/IbQSMlqceTR5KEsAbhQd6v82XfH5cu60VCA93g8
hypiHUa/AFA/tbpHsnyrdJ8iOxnU6NOwMGSOs2bJ76HcmUDphZQQuS8ARfAB3q9h4YVJo6wDuBC6
4vOpUEfR72hKl+SA1JHnJO6bpgMe0gWxiX7dAnZNwwEOLaIrWL60TUD5c1C3eCg/RESN+4/7u39h
nlhMvlgG8NqOWneJSO2EhfWqXQKXy1CewU/JZpxZXrmEawyX100L+STvkW6XcAjTqNBGBFFz3FEm
/OcEV1Ofds2WUBDEQzMX+FUP4AsDGUhOXSReIoP6LsrHFBajdZfXfeDLmba5W6bSuVKut60setwy
I1oKCM4duYkSDx0Fy1LXlYljsgyuqYeQi+4X1wiy2yRZZirev9Te6JEl2ZQAbbjxprjQZljZxn1L
LgmFm4HxFxG4HEeJt44DPXs4MK5lhpF5V8H6Gi4QZmwvndIIl849dtsH+rlDoDKCwQtnK4XvMZV7
fSPGtcwTwdtV8P+cMFFP4Q+LMGQqxC2prwaFcvTNVPYOUJMefIg7KX4JdbWDy+yQamacwwF53hJC
571K0NkUQEEFcyIhNNY/tKAaJIHXo2VnCxNClv6E0cuSocGCxF68itG44gnQN8Ktfbk+4Zt0VIBm
0wCrMx2BNkpOHK9YyNddqUNorJz7u38siHbQRSdpZz680XRCXSqPonljKs3QHVmO14VkVIFKF2QA
fcqeVVmIH9cyf5m8kcPvehglUTDGjaJr9l5O+nluhwnoatFoGUotGrd0NDv5iR9FwQREkUCv5jaz
Oys/F/VUvnhS8r9LEmbwxhFpHp30AUBxaIJ7r3Zrwkw/0G+USbBvLtkihJ2GjDPmhF3OkmnDpq19
DArvYqVMUOifdH3FYUvhIn9qavLtfXzmJWBeOIqY0E+Jz2maikkYUVuqbMfOVwbmpHhN6SCFx7BO
dUkMLMtmt8NDXkr1xhOcN/3kPAIRKoZRMeKvHF03plWCiDxDBN5orQpDca1aGMZBSOwuL83St7GP
X4kyBn+ZjIhsc1sHQokTzpY7H+gyqlHyx7Etadr5cDJNSBH2VKbz0IdGFZONpxdPc2PjfptHdfLI
mtB5LH5aVz1v3IIgXSk4wyiGApbnzxsK6FIIOwEcXgvklWH07yFpt3wrhxj9AJc2a6xRTJRlORRn
JGwAOQLAn8irSYaYD1CTp9NFMIZNBOdKC1rMpOHXHoKDkgr6GSX9nfx17qMLm4X7q9dNj9sTq2Qc
gfm6zcLNn1fT8CWIKBRemPZwkBqCBBirm8K4g0Oc6BEy94KMoYLo+PJhfgHwphsjLuo05xsT1j0t
V+riHyWp4FGPdk2rbyfgpDOaVmPhXLBF7+/Z6rnawVNKRIis/i0eu7/VwEcAHhEIrGdjvJbNnLiI
y/DJ3xdFhBWZmLOHpkV5q/nd3LeWs5+ND7ncSLheAYKw2PAw0oRPfBe1xOI8XPHG7Q/4KaR031Ew
cR5I5+vQzbv18y6MD6ySGiGLOtudh3nkYnzSXGcnh0k2bftYgk2aWC1oasFMJWIGO1m4VqD72QLW
/+0WGmHSwgemQnCbOIZ/eEQcovmS2gftLyAeniFymZfPr3z2PB/BLeT7Gdu/sR77Bl89wgjk/UlA
Tgr8DzX+vqQDp24Q49ONqYJxpfEM2YjVe6CnsH+wW/CYwrxWLn4P+tywTYbnzgrKbkQwvwJOgKxn
v8fydXhWovWwF6mxa9Jy7ps/YkEl72lsSv1Iil1pn9FIoHxBHJw4SE427tEg6kv3sdLODECDBljm
R7IZWVkDoy7cF/gqMxiLY3J+ycJE8VpYqZnSZyx3VSi4omEaW6EhAEY+LkdH0Ffs6wFu0atN8Q60
uj9hv/Y7G3MXWtFMWToWu4Vm6E9j19DfERB5EmqCs4ldy1KJcKsRN9FEWocEi9mfQkYrttwxVbkQ
Ck4dUYhGw+iIGpwATa+eTQLJ/WjTjuAflJQN9OznHtRrG4Qkit0kCfR9Ls03IVWABl8ZzlR6gRrY
4IZawntNfXfg/dFnXgaA5Zau5X3ki9Ic55BuQlFt2Gljkx/LKGbxXVoW8nKRfMU0w4SP6iBW0dGt
JBRFCo2u7tY1MLI//0nkA1yM73fXe618My2IO2hgox2GLtpXPbVkvKtqlN2aRd/FbakSBk7O5YBS
kodhlxrhIsbSAsLGBnfi8ydh5xS9vjnt3jCmJL43T2Dz4IiJnsOcJpC8/O7gQ/swPAgOoAwhmzl6
bM6QlZkCAZTpPNY+948XMWeW6cC6DAzRSSfLnvygz7uA+fea1phfgAyWQww3Y43sd/PYshkaopFO
aGoY9ZjuyCuIQrtFL45z83AP5er8QvhsmQd6YBGIPP32LuMyga4AY5aFhV3nYhDiTgBV8ipz3/io
Gl8hXeQwDe3fUEDDXl2c43cvKBydnHTtUe8lp6yFthUj+ctjgfk04hG3RfEwBGhyDwEqrr1N2+78
ww4jEwra3w4MUkkp4GyjEcAma+/Y2veHOChf+nTFg2PQ9Zq5pSdgIcqg2DhDEfgO7ic6afo+pdLv
e7VRsYYFjulgGmDFzxrDRctVhHmTdzEBtbOoPpDI4Lnn8YKbGgQhNBrDk7hb9QANIB6JmnJ0coua
gK5MVcEw4XoGokaF1IKuyuTHOpMzl3USytRBIgtE6dCrfzlladg3jcY33c5UAbQqjtIVyVQuJGci
QjZp9ijhdD1Kcvxqt683ZH29RxZJ6RVQHbkKhR6ckGV7wPyFu2Gu0Bn0RtcZpKkiFsdbYRSvivPu
auV5A0kcxijp8a8Kq8JrQzCuMuQ9zUGXXUl9+td/f5uHEe6Z4icXXGmiEgcWySI4vdbkku6Ouri1
6tSHUgP98wq/w4Ei/CiZJ6D5HN5Xp1nGm0KbnSQFIBKan357zkZGcQ6vK6pm0oglr+Nu1Tq9cqqx
A6GNHmzF3QCKk2GoRGB+4Iqze/g2gIJmUtuu9G/q6AV8qqHeM2Tfv0NPQ/jOHUOQFcLCHlTuynZl
8dZgcx4lK1H5NSNt74LDXLayfwakbJRJDfP2ClN7gScbczxG51t28BUdzd9pRxWa3YnIWe5tapcz
mbkoW5waXHJcTnjA9+37bSKpE6AsckFESoTu06Kz1s3XhftzclFG6G/WkBjiWK/lmhs/MWnSeziD
//GpFEF0yLYYrF0l6+AppCRLOFoXrNEKGK1//tjPuDIgkzQ/mffUTKj3xzDkuadrWjWKfGBmzTjH
fKtGuoMXjo/kAqTEUf5LRW3Xr9rWYTRt2YXg6OGxiUlIoFzr8c15IOwWJ8CQcQYt+Hw5JMTfYoI+
ZtsU1wsG4Q9XuCdO78pwe+mCR2NmoLDwuPcSEOhcJfQrpzDszCkHX56zKEcoyr+YIH0fM6C0+zVQ
/lGPpFtoPsDs8TZJWmnqyOllXlplt2lFfcyzM+8q3EdjI9OnpNk4PhfGNZr/MwN4ZOdzOR2PoNvO
og5AEIp3TQxgA4GF05UQCwugbHuhVQ6hq7umLUM74c/Pmq7+pLAl0dyjPvQABcgVZCNPL6V1IkXK
3eE66f3XY19UgiDRU1x6b2sOIYXNIG7b224P2LDJhMxByRCysm5NUnoWKcnNOnMCrT9lEc/qyAfb
WM+xlYfOC3tV3HT9dCaXjjKl05S2rGrKhaXnisnNrMxgOwT/FHzoI7O4xDzFmQNdyoWcCfFk+h1H
eQxpfEUAPqy9EdIWWRk3+vJlBshIpojK3knK4oyEZb96JCnWMLRyh9v03my2wsS5tyi6ro7tUOGE
QGxqASqkGarOJ6PtuNFvzdukAC4DQWk8vvGrHCD0CfbMFBlgQGunV8ZaeaVC0512sTNp2wqn7WI4
dK30ugJ4WOVvjmYG1Vq/QkXjf4TJx2dXC56fqf+qG1uMCibBdbyC8iESFzJULV+wPvbzEOvcuOiD
HVY1gJD9bJ4SDjcCIb0jG8XC8Lt2/NaGEejnHzQR8jPCiMDe9uFFFc5lkK5WIFVtFEug2kQxjwVh
tS1p0U4Q4V9Eb4rhOCHK+KbvfcaDZlUzhRkFIFWb6sX6q3+r3CP3qC1eIZucL71mqCxTsmRepAe1
RM4NfkaWnK0BN98UG9uFE4ihJ9LQPdf8wn7APoo1+Ue7OqLFcDJPRbY4CLY23rzgg7bSlt6OQ+Z8
eg3Id7uHUrYuki3IUTp5apUgj9q1PVnvCx0QRZ7SQaaXL+v9LKPXjdcewhSZcUpt6cOdKuxSur3Y
PBhZ1u0mg40OVzBalJA8UYxPkoFS02WwkGkoVuwEj/ICWybL3u7rLmD97dGCR+vItPc6SIZbZQVx
RTQLOucYG81YnM1RUMLSYz0+wtAjcEmM97GU5bTTj6NxvHn0DZz4346fMr1wvno7QXjfF6OYrCtC
ES4fwQU+/Cp9MLSDLpRw5YPzjMVXDHewIE9nCTofySISpUeHTdOpUlQqjI1FNsYJ9aNmofuKaztW
4mG79QvQNi2sUFj0hFHW+kCyj9icCymnWNbGOwwq0sydm53gb4qP7CcDrniynEgPpqA/aevVoEuW
mDH6JbrRFep7GGKBLLDDaIMfZCM1IdBTsjEiK3AiSB8Hx7H43CFC/H99znZcmI3Uu97Zs6IN0YZJ
AaoWbdNrtoKsEAoX+bUaMiaPJI/wrHagK0GFLnfCowB89lIBYv9R2ilo4NPD7WTwMJ+SgcDi7rHx
i6oJNZHrZudtcDJAS+QLHQcwlH5jW64Y9173kc4QWIyj5xEB+et60+2YTYecopCQTnYMAzur8J1n
HScn0UPsMslF33Sr+wRUqlispAINqnrsbssUgg5ctQSy7L+nQG4yRmvCSir2IhkXcvTYIMDyrbk3
6d+NqaB2Xco12Kzx0sAMuY8wpO4/bxkDYxnpH+aiATrc5yKUFHJA3Zdbk8CUiWqsrPoAfMt41ZQL
f3LNuZicWaxOJt6EUeo//oH6eICRdx2i9J8aky+k8ZrRP0mvwxg0itptpOvZ2Fwr11ymAbeOsntu
DEqZAdVMy+m6Yi7yiqIvfrx6z3+mJnD8Yk2EmCcuOt4KqCaoTSZCDVkLfHrgV3O6osalCOOY5etY
6zVyMsZYoMDMeDD0i78fELsmQOM9WUCT1JvAh+cJuHnOQUAHGIa+b8kZlNC7vk29X5+ueLNfDL9A
DWi+XtjqNx0E9VuC98ZistGB23P7suCrYxOXFcT14SJOc3YG60v/Y0nrNz2pHkdXqN24+0fskkr6
63RfVXUnEc+kYEUMPAy/thSyEjwnbmLt4nauGum0/P7YA0BNre2Hox3+Z+5XGIE67P1Q1KeNVQYO
XbeappF/c0yNQreihoReBr6lhAUJfzc4GmM9WMhAUCRj414lL3ULs2S4a6QbWgqeciSip8JI9edK
afmQYgT4WzC/6qRgQwtxam442SBoPFyg7U0wqAFj+HjG46aHyLJm2dl32IWwl8BQTuKxelA5vJ8q
VF+YKhZYmb6o4o/EEs9fDAVPmyQt4A8ZA8FDstWCo9CC3cMlax3jawotPl+4vaU89sqHp+ws4Xc6
jPyp0GSsZcaVi93KE3ctnCrFGou0IOl3k+a+oIz7Pao2vP+jeXrvdQsMxuy2iyKYX4Tl6bGFsf5h
Rc193gvxAoz57lEBV9AhwregNJXF7BsC88hg0/eHUpwKD1a/2QaF73ZCedeWsv+lx7qIcHRc8AwZ
BAOBeTKSurrjNnlEnZ4X6xN0Ybn7BfH/oLvPGR02k6qcGOs3UmGNLekma9gU9sVWXiskVn2UaYYT
HfaYenBqWsAvBu/8bQiUhCtGQFHqBxz8DbZhm58nVWhOQH6abzG20e9F+U+W9nq5MPu1htxz6RGP
VNvVNNyN7GMBKDMkKImFTu4cYEDlmZmFDlqecRD2SBBtvNVyrXNjvWmQ6Mxd2Bq0UtnFsk/dK/29
bbEqrVeNAZ0qrcTjhSDokkheFIbr4Rb9S69wEtIjJY1G2qnT50LIVYHJvgtlClUeMlj0uXRK3i7g
i3okKrPtODSHYCWhVxfCG/JgurLaFcRQKZ+ENr8ABNuNzivvYl/N4eOClFgGYEs6PIrLVrGmP2QU
krICpw6lSmX0goXa0fTU2YL0UuKtS78RF0iuTcdABWk+P6A0wMEi3/rT0DK71LERxXBlNbtE0P8n
J4sVNjJpzSnQOTIWE1QSNS8Keb2wEnK1SdzN/hcUpak082wJqfA5vvi7PD1aoaSYciOUaZdnUAG5
YyoLLLsSJg5ftB5XFzK+7q73fRYvzdzK6ehMx+Iie0LRJYfIKyyOGYSdqsVDWCLhOGv1OuJeqLrT
9y2Bo5Empbl7ehInGFa59HuCamJBNK1pp4WAvrLwG1YWUz77YVy2nXOoaNYo2CxwNB7/S9NcDBaE
hjGynJxqqRJVniYuaISYosE5mSqhkbylZ/8ysEGJdBFRwuOfGOP/pHF/nt5TXb/Rik4tFqSAf3ZQ
/HUmBklpFMloqE7ugVRqk7C1XGNE5FNRdVSE8H2vED050qfSwuYq/ezCoKSfuULc9Z0I2EWvX13m
EY8kSvxJ1A6/ZxL0wFlISAqSnp3yA6Ji6dYRMasKalA2y7rgJdh0E79clBjBNiuQCAjvNLBJNaiy
9IvjehYS0PZQpIbsdDTfifFlMjqYhSV+udDyyYNga+rr3gGYBBYH9MBawcqg9YGkdQM4dJkEnVJb
GaGJSkZh0AZLuRMjt0cnbmejfvVMTYRJ6B0MNRgMOqaJR8HeQCcMcYz+PNC9NifnyFlta4qbZS64
45IWUIrdwlR/xTVlAXC7zBak0aWWj2DCdNmFFjndBD9LjG2e0Vpg++31eVlsKoCtPE5IxylMZr4G
j2BKLqVL1K97E4ZziLwTp9eaK1n8jEnZZfbUuLMQ9LpVJKr79efG8gPaBRGLDvqRRCCOYZVVQE1O
3Ap2J8uCM+p6CACebJx40o6bKkTEiD5xx578XaofGJHiXF53wjfyHzMUch1sIxhO6XBMiW+VmSDh
6QmVD2qEEAOpWSnpGGtviFjjJ39NRgh82FCqQrEctvhV+oeKPAfbk/A4RQGnL1JdPxTRUh0ieFnV
oMRJViMVTn4JKX1jcwxXc6hBeugn2wxhI4ig5dDGEPyvkjLu47fGwUHrksl7tpKFS6pZHcKd0Oue
F7NnlKDwaDFSykGdzn/qQNdjwbXy8juL03T0KM6TxY9gYf1g2v7Gbh/SXfuH6TT7L83YGXpZBRru
U6F6RoDsYdV6olJ5JPGj7PALb+ysbUVxi4w1eg3aTUnjLJtH73SJbxUI31vo+qplPRVz2Txr1dT6
895yrOh4CrFDy1BuzzfYW+tgxIOxO/Uzs9W7G98pAD/rzJNvmbnJFqCTmRgnXmta14VjQk3YjcoP
Uk7b7DDhxYZRz8oNG7kjbB0XGmBKk+v6OCnq9OK/lfdjGuHHr9ByAgtERNTXYS+o0x4eQK2ZrOrp
urnwB6fEOBwIaSWkg/lzt2ZF4T9d8q3b89TYGOLeQT/BDhmX0dJU21jOFR6aJffSY6j+4HXsnF3b
ph12bNd/tiiG2NGH7JBFc+s42JL/YEhlED1q+FXwHd5VJWB0yVl8IACxCc1zTFsuJSQVMmdJR2gx
KF5M299hQcqwh6gl3n5Ye567Q3oYNs2jtQjeg/WHR7d5cY1NI1dWRZ0k5SOVB9ldo03Ijr/4nxBs
OdM5IRIfd3blkfkJaM3AkXTbA+clkXjjHLRqrWflVGL4w2HacIWbX1Kt5C+OjcDpsSuRLq+/s41o
JegVrK/1s+CLhY1kMuBbSokagHRgcsAwNIqGWvuPE7KnYtJ8vk39r5qUJt3gDpwVBvJ5ngYdmMnE
LLy8skgaivgDEvg5B2Yob0Rk2dewg6ISKSrL1coi6HxGKzgphpAs4xIxP48fVYVZQ4zgfaVRP2iA
3eBMSf3bgB7H1Bdrm67enIsYMpeNm7LGszUmv9Hno2QOhHjFcixrT1lawZkGzfBcbHGAQIBNQscy
7Rt4Vl7dO/2lxN17keZPMcInCGiqWH7zUNvkDlp7js5o1YBNKlEo4E1vtTJwXzrBG6BflgRzebDv
buF11Pni7l0gALDzti/kL0Kd9Vim2EpQVO5XsLcVO4fJzH85kR+/ziW+aVmY3bp6QXaa35xunfw9
QJCQHwM+0Gtaa1fwRxJg01dWaaXKmaf7Rcg2kqofs2bfcocUEkbI5+G8y4WESY79ZPvaBYV6lkR1
92r2iGAuCv/TTsPnBBneiSvEBFdxl3IdLJnJIICQpVuBoX72YjwlSBFjTZ6gTiKLa9X+JwraZu3P
iSiHfO1pVcKSyegFo4xrZAUkJk82Y6CZEkLW1rNB2ILfajLlzZG+sTZxFtfqnBh15/xLwqTTeFg6
2RTXghTu01Lji0cTM+Bm/OGfO1z+JdxyUSX45t4wu8SWZsMKbVrOjVZlqccVSZXf2w7wcxBDTDj8
lP3R7vPRCfXjG8R3CBRChLslXL/u4tkosU7RQRqTG7pwPAa4M0g2ZkZxuSWNZou8uCPHYdYTnjGW
8M1KYQudx28jM6Dq/yUERvUyL0Dqi9GwoCsh7GSSTAojyMn9Exn202I5aN6KXQ9cfDNQH5pprpzO
P/5yhep9IZWIAgO6PaumbBjiRIn0/DN1PX4G+ziaiPmYjhurpjnU0VSuUsCmh6TkwZ1qHgvRZaW+
kUydjGQ8TpqI40TcuY+XkG9d3VpzRUqBYuj1wpmoYMh1cnusSFG9XS53PtN+V+5cQtJf6teCR+fz
T6DBRCmA3tY/2OmU9/G6UiaKJULxL0Mbr2SlLiXNWCCxKmfW0sX6DDXnm1CclWSMmDaW8nYNpIWm
peODCVT1LLuX0sgRR+SaQ8NcqtjCggLVbdwqMIO6/mJLpSy/uZqeK62f8O/uaAaDBDABUtiZzfG2
kQ7ec23lgHAp8hF69SBqrVU4lAoM2scAaIy5cEt6baAT4W5Wn6YFC7VqeciiD411Ynlcxjmq6xW1
rAJap5bdI9+8kCD7C8ZkoPXdSB/dSERdk4PkAO9HktN6A7ON77wlx6GAnm+MB+dphuZjjQkumNzU
cFmuojWwHUY6lLbG/vESR5QxHKe1GleMAzliTI7RV2uerQwMt/SWGxKgepqCW3XvATj455G95BWp
Za9DsQKeMHOaGv3jm93/yuel7dGieLEyjZ7uSx8KojaamHCivXDYWFJerDVO0/399ET4nHpTvOLq
5QhBlOfB3k92XIx6MyphGVrVjsJjyJvm7MAgrm8wczO4YdUI/MMpRjeDSJHq1swCP5Y0j6RPlyIZ
jzTxeYinXhlQd4ZY6ALfNKGhVxB+2hSKNMwBEqyjlRtwgpAqy6eRM/fn918nNHVc4gFw3qlBgxep
IbeRqV4rmrE4GmIc9SbRx1c4qeWqOR7chmtKE2nNb947UZ6tJIDoMpJueanftJ3++/j/XExWSi5H
Oo+rvFvZofZWUMSWngcHHiSdEJ2sKz7ApDo0oYKIw5aaLU688B6CoYPc6dhFFatz9DbjF0fA+gXX
1cJJLQNHd1qutQMisuAOc9v6gJcaiPvI+HzLoOjBHIU0dGMcvxj8AUm+2Tis9tbhiwMHbr4Hn7sx
UlLHQPa6BL3pDsY8T4pT/pmvpwK/VYMYmsBRg4chVbLt/l5ttwGrZeVaC36kSNEKz2XTFLrnBwEq
n7pZE/TYXzvEccl2/PF8jzsOfCXGuEZRapjT2OhheU4s48/enlCdyvRkpS8imeA058Wk3Z9T0rWg
8+dKnI424t5D6xlcP6GyylrrbyYPow+Wf4Gav9poyrmyCi06Ts3nYnkyXmw/yVSOETra3ay2+V9D
O62pOVzF2nla+LttVAgf3jQuhjZ8dJkFJAH5eYpOV/6Hxxf8IUh9h37xVEfht638h6H1dD/AFziI
Ri5e+wdWuRIa4eBz3OftKQMPn6FdflRDto86SPrCB0woqG046XM5fCG20mhxtPytEqexvWNt8jKp
CO56DzlPbqB9DLPa6WsD8OacMAQkQwuGuh9T8FbwIuNw+nIR+4FoAKQahzPee0qXpR6Rt3XwHft/
MRd8g0bsGoEmqhhqklHJiOZZrn2M7t72DZFUj4lsOX1xij6jPm8inHl4suk2jXn58kuiyRCP7VDp
OPDZ3oPVQVtZ7uZskda3kijv7+VE7dwqS2W2BqTq43LMD4JW+zCdnQu7dHtTL4i8x6gaIFKmIND8
KgFUNxuapB90woJgRBIAhIF+zCLeeLa1X3I3tEG1OxJ/CeJA/LKSpTGzaj617KVD06ghmcypTenn
rROYzACEDPB8uPTx6TqUy0WQVFpMgTFsb9dTnpF2RdYJEmUDkxNZ2XyRjHPPu/bO+MbSSXX2aRFr
OpvXAGKLpd5NJPyx4LS3IPVFJf9FmQ5kGO9q5I9q7QIs8HTRtsSjbDKH9mYfJne/NVTWREsL5io3
n+SqIskQ7GEmKhGsmWCO+t8REFLaVemYMXHRlCnG1903W/K9EO2hxC7wJpK1NhaaOkqYhNnnA8Wv
D35hf6Ee0aumMRnQrTHb6UUftL+bMebKXuBVHFgnG2JalJcAOgOcTaykIVBlAgQUPh9tN2vlOo6E
AQlKcQuo1Q1LSJUS1ac7jy6Q63cAoVuC8fWn8/Oq5nhYShtI2SfNjpQkPcerXihjIfBsCPt0q/uB
4C6oUFu55Vr0TDvjLHa0ai/RSZcr9M3V8017awVM6RypGWZQEHsw1Z7AI8lsYe0/RpRhqTfyhdwB
WvIGB+IpmgE8YDNy4Mu2ad4/oG6sfiio4dmTBXIeykvcmWVVFpZnrK3XBl4NfMhpGcAFZvNxidIn
2teYyK8n5F4l60HvJ23VeY3xU3MVadFZC8VjkOK7H+5oAKgFNlAVD1M6gAkcU50O1+JrbpBc8CTa
lkgtC+SOn6NvwSQr38zNKMfvAjiXbUeyfV8r8gwdoe520C5y/3/MX61NkuKxPB7tAAvDcuFuUbNE
lhaYM1pIfh0AjwgpSkldm8rz9ZkGEsgYgVHHAWiXl0w5R66h4FMbReTyuScW0hTT+DotG2f6bORD
MyfxtL86bBGrjxRyuYnFF6yYtnDdOrETJggPrvxangFpfTBPuqZrYp/InMmG7T5ZQiQf0v24lc5w
e01nsVHro0WyMjR7VVIFoB+PfWR6m8+eB0V3Bkgdb0YxNc9cWgMSk9AOijJs54+m4chA6ESO6pC4
6E2oCRpdgZpuxve/CHrqIqufcIK0NVvDLinXUddr2vX6ywNpEPmndnt29ggurQMslcBRjrk+ZqBE
uJR+2+4oHdA1WSE0SSDx/ZpJXk/STrb+c32PL9bmE2tmYD47ZUAPpAa08lHvnVlMZ39+eGmW4XS0
7gNLpHPOB9KsOJhVafOiRVsEvFGwb999aTsSFbLG99q7lerZq7N6K2Tst2ODC8M5K7HNSLkxLina
aanZuycp32wcy/M3uQo42LBarhC7T+7cfv/3mIdRQU+ynj+TlKW7cl83ayEg17oXZPjAtI+9o24D
NmT/dY317q74DBZVySRwZ2p37X8zDJkEdmNuoa2SamHLwAf5CneVctJEwcOghCDGPPoPlZI+Niik
3rzY+RnC+7OG82Ojbpv2nTcpoly/QAQPKebE0uEyDXUfMsi5HHYFzH4EDgiLdaj/Hqfeiuv4wOD6
+thfTGnAz/fsXDyaH+ljgXTGUllNGYLko9eualKsYNNI4CJag1MTJFyqDdZ0qA00eHo32F3jbmzE
GRPabllA1zUjATLWgKaLsY11wyPFlITsukxPLzonHhTnweqp3sjpeO9+C+RftKjzeu/ds9oINVzJ
qpBMloyCegWg9hxzHXUUgPN8KIKgwpN22vFdYZ1fHxrYDQv9svDWBnqZDdv65+ShAm/PEQNYhrue
l65tFh3sePTpbdyNFDEir6YPs8cFbXpzSpR7tKkNErCciSOTRacZb7MowLZZZD55P4WQ0IHi7n+M
gMgZtHSn4qCVwoQact52XtRnjQ+ht7ncKJCCtlskbCdmOf39OLCch87Vy9dtNyBvop7nd/pQA62F
0EGWagBgcakK2jOhfDtOAyK/ajimhzNToA+yv+BAAKXlqfwDXIjeL3KFHwr+YLR+X1xTiNZTUafO
EFU45U/VNGlnPm3ZJLwbtcl7PBQOb8WTdJKp6F3R7NPKTqaMiRCIbwT/VWPAAsn5iJPyvdivSl0b
yspBXtvO5m7+DqXLtS6vZaVc20XO9rbJEUlJ2m9BwZTAFUxLdyHdw3AX1Lcr10bhiMWq24R8Mrxo
KL1kok5HAWBFd0TdqfH8WUgF/hWYp+HcGE/xskQ7tZH3KG5BVd26aYo2ms382luxpLCP5s/YmD6x
MjJXqUNKuRW6X9enue1N/P1Bh+O2dFvcA5q+sYJI4vI/lcXexGHevSYrKbX30XeYuYK3tEa6EaVI
nujWOg0UhglP1AKDi74wzIRoNrfJBzk0EKTPsrf3oiODWifBGOvXx7P5NcoxbjIYh2fRI5uaXale
um9bWftYJQIQTvrapAQONQaG3UsL+IxuUH4FM5Sdj6RX3tybDNai3C/Te5jm4QjlnNerdkc9QNca
D6e3fJ9wPTquFk1zIDuEiEPKUWerKcdspaxEfcLGYwiWEuUiVzPW/ICljUgWzhWgaLOIhTOTn6Jy
ZwH10dlkg8Vj0Dy4gOvwNXGb7On1sCYB+0LELEhUSpCfYhU95Jwk9Bo1l/iW7l5a4sc3Ch/h+k1n
QnvuIBSM80+6JdHE2qgD32Kbbjd56ZkvQKq9U7zAC0yPn9OpT+fSXg2KkDQ+CzQeVQAix8jVU/aY
WpvM9tOZftFKwzpgw66fs7CcJ7IlL6FNbRaJlpQNBu8V6zO4EG13MMxAT85EHERsWqF3ZYn6copN
ZJeFdIQVgD+0hiDKYst6EJWCKtxZPGbPoLVj9+Et/2z7iSjeO4eLqUNuhiVN9s7q3dlAmHYqeq+r
Mi8cg/Zmg6pfSo+vfNT+SgOxHS0QJRRCU/NHcRGv04uaWr38AmlzhMsXHq3SPYlJtLWomJZFwxP4
klRqX97oABNLKMbN8dWwA7TGf5qEVA8Fc3FEFGPFvZ0V9VWiEmQpkGQf4ldbAvBmf98KM4gKOoe9
pBxJTIbMxJhY+na2AbFiuZTQdBOZB+1FBBbMptB34nA3KtlJ758Kl/9PkaowXO+aL57J7KQhJZ5b
QFWkkyxz/Vyp6K7NZeoMF0Q+/p7xnxrYRv9T0cV7wayGUJKVqptoTgpydKsTZwZYzvOUUSRySEag
ZFOgc1UCNVAbq4/5rPaINbT28ku8LSt1xgkssTGbbSJTwj3efOpd0f4rAqzvtHDckGQI0xwslPBm
TJZntvULv0VzFyvd1rYNR2TvcfKJYP//akaAI0McOnDiR19kzHKZXQRwgrwZ0rKF39nvIZF4cEpi
+aye6jyHyfpg/rXVPZWCF24kiOsuaLElV/iEVYymfsg7PD/TqUr19bP0Ud+jHO9HdA82i1i6Wkvy
qAxJvw7qTvRhK94ek+InyclHYSJJn7EzZCKhlj2aGRrh3BWtvOftcaaU0T/dUxodURim2n08m5UC
+gvxooGubJCE/HtMIMlnQmu1dcTb2aZQ0c3rLg/v1fTwR35zHD8I3oMli5/ysKFi5U8SgJNsGYVk
o93B6miEoOhDnCLH32Yh+/FiNV/leqP+Z+tW8vdjko0HEaOLu4HbI/8RzL+jEjJC0t+eSu1A2GM3
yM8FuH0bQFIJM/If1ZO3/5MvQGjlG5l/ByHRRt+j5VNNbD7vRJra1jt3ucSnRQQcX6oqzUaAHf5W
IfDPel1qvnuOLy7vqPxBzafIcTKSObfkFagA7pGNQ/cC7zR1haczp1OVaORpA/DXVN0OIwRaLJxd
OgfbOwOdkT9P123/6q9U87nM04gIsbmxcTmQNYKofZSze7Jcw3e6uL64oNMgyjRmOTYdEQs9/nWn
MBciiA9X3ZQg+WJgO5FhIiFbb+2fu3G9YfoG5EBfeCP44JgKjBpGR0uo8skTKyTkQxlxhs20aDBx
qlKv6n0H7LBE5vkF/SanelWWDnF8tYJDNvrJng96757IcUPLKd5bf5+mXCMYH+H1CfV6RUjlLjnK
jNWi0bfIruj49fO1hEqFl8qbdAV3o5kImidGT1FM686KdhQOTcUzPFoAz6FjTijB9boGhSdkTxOv
CqqeVHLB1nKvLdnqrA1vJaUXbf6kQep7GfPC8iHzEU+je1RPLZIFOA7SX7i5FCntvBQLF7+TZf5+
gt+4/NNL6fmGLTN26FzWsyaAH6eib5qJOqVV/fdLMzmwlFuK4lhxcGxT5TwCsNFTOFEHLVy/xUlz
YzWtpTcdRuOSVHvXpWWts+TOV/Ht5ynPM2Gc1g4xvs2M6hO6zGvCyK7dQu8heaTZxDymP75Y/yTi
1VITXRJ5wePxmiGE9GDVJodlNgdzbAG5qjVNwe1qLm5SwlvaMAbn5g8kFMKmLgl+9VuKYugHCLrS
Qi3gCmuGbQ8mIifcO2PpFh7FGi2UX1n/G5OBFGWONeuBdrtaHK9gLLwnMVJYqXvqvkY7g/HvEgOs
DDCJDFxBjJF6yIRN3LVh1KmM5YJVq0hCJ1L5MKYWKiDlF9ogRpYtOeOB7UeMzNic4Th/OHo87Xx6
4jjRaMYh/mHNa7bBTZSjpjqMXbahVc99JFvHSlSu2izD9RbVfYKg5LjFioWy1p4Cej2waYek2D/W
rYqsFG/BN0QhwyHOk6cmhPPetea5MyrIUK3+Dj7xiOhIXcbBwgsoluHiQULG+tbbHrugL+bWvw7S
PYTXcYAUu9ZH+3Tbl/zh0oyEFt+e/M/4stqLlgOULE0RRigi+MTwYg4iKq35ygkm5wJFhAAKjJvZ
lX0w7XcT1WNakB5TzxsPGTeLUznFcbgn/0ycaOmo8gSr6Lp6gKy3Q2gwBSuVmcXotYDctdFhLc7y
7R0FpLLvZHPRZQBbxp7VckOhrumDQxKqOrDPP8D9FsgXFwXR2U9kZa/2D/mT0R6/nIdv9ioY+9Ox
tLcGuw++1K0yU5Wo/ZOu0okP6i9g0iMiQZVvz5z329jgUMGloAbaxQ8DXXtXVPCt+wYm2iahV3ji
sC4pdp2N8LptoZdudGQnaaCLDuyy6MDxDeY5A+HCCJDkKTdMlHPSxjiUVJflja2auGpJjuEngEDN
J+aMBOnCR7eqWAIMLpF6/qJ2G5ioqiMqWkRYn+JbBqjayLMKUxofw1RrnMOWMKnYJhsGjFAkR+BN
Gu8nns+UYcL2lJtIze0Yui2D/qAVYeM1lQwxZUmrrWwd30eEgJd4lXzHZFd5XBub/8jTTJGbqHZo
9qf4v65kZWvUnsabGtv6X4WMbwEnlucfhwcJy1GqGRmYMNHtKa/or7AFVHPq0DgTp5bK2lTK+hur
Zkm5Edj3h61/QqUxfEFKIX1n3dfAwAZ68GtnVcM/NjeVAP8kaiZggAh/SI27E5Xqxt4YKNAlfBNa
nOF8J+La2As7y6M6FtVdGz0H2LiFEE7WxqZy+Wy7mnaKDXCEoMGMLtELcTyRrLTSfPBQMBwMu3jO
Or8xwXpFlZsKBwrori3pgOJiZMy/LYph0IQ0NrT0VEUAu4HFPan3G6auqnJEbxSF4pgoSjXducPY
0AVs4jTNRbslGkmgTqvlUA31t0Gsyxd9ocbs74XU3r4/BPQXSQPZMPCz5bIWExwgbMOaPvpWt09c
dTw3RTVdRwQZE/Qo8M8t/AbedXtlrLzjgAPtSFcrkB01IvF0rebUq6LhLU/AOAh7O+oEEFLy322z
cU8rQ853BlCyn+zizSx47RZdSRaAGCrNdhhy9EW7oxs8PpK2/luTCD0I/sH3442LKpQWA0HF1pJy
GJrp7UYEWWgs1ekOzMCIaeiJrQK8lIPoxl4KQkPfPnobw0XlTnTynTHEl6dbi1vBVQDcF5SNJYmc
AdHNC9kFZGiynAWS19Ttkm22xoKsPx9+LjQQPIXpshlytwBt58i5Q+ooTBxBNeRolbjKPj0YEqPg
v3wzC94LyURd9DJhwwb8XLsG3v1M81ekpkIY3Ul/qAB+Tu3AaRDXixbtfP1CIH7nhw7eH+0171x6
shWzBvoe/6d/LuxGbs4CbmhffcNMkflw52rTJReZ9uYHRqdNjyamKSJg0jBwTXxpAbgufn2XR+NM
+OwtF1z0HTUZk4wd4xQGCp4Iy5VEglGqM94bNZyKpjdOvROVCcMkVPJ332HHVgUdgHmoD473D7+l
Tk1EVIgXB8mwbuAV8jFKtQPtP+z5xhHNAwrJgYWTejlJ/UEqcKKSJPMq8XEy5mpyy9O5gS7NgxQA
ooqqgbElns0/1+mTngVWHQxaN4StxQ3r7+OfYwwiSTDqVFPvLRxFhbwNCBL6mk/+H2NUd1njpdbb
dGbiebrc8AdRSmRXuTcLUaWeXGzxcWMHhdEnqapeQhWCXZ0u3DtvCplRuV5DGCI6Gv50oQPlCYyf
PFfEV84AIMTpUekLanMbYN1xp04nxrkCchxEmJw1TtNOiiAUTB885dX4c+bZbNMYGi2K2ei/fKAH
r6OmSzMsuovSPEcyjRDa97XWIfBvijpfVyPKSt/s5e+MoFo6XUrO0twFog1nHJjMI57uBqvQJ8+T
iK3y+ywiRhq71zox6Zc7hI4miTSdZW4HW5JiKf1bTOV8Ahvh+2sQr1dLOWfHlHC/Tvz5Ftlb2I6V
sH3T/ymjBfNc316eeWfLevE1GLYHYcNzlYacboVn+R6ajzLc8phFCxqHfMA/nAqgEpDjgx6FpO1U
zRfudIzhxfbspXF5BAk0gnPo/u9MByqRH518HbXksNC8f5vyCC2Z32jNARBtkujU/PMLTT1FewHn
XJJ6HKPw8Dj23no+75xOV5oCdCFAu1Gbu0wUIucMZ4MUl/2wnHaLT6TBvI7+RbVArIibBbUYcb2N
D3Mvw1tfOouZiMXzJ9H5RKVEuIMFfvSu1ZhU63d+N+E9S/MRWygG3pArPAPbDErw8mRspPFF3jOQ
yOlq3gVUvh8xW1tBgaXKL/YCXCAE2Kk/jqA3PB7OkgL8LtYA3Pm73OFhmaHd2ha+fuvTOKaXbMu4
OeAzNEMcXNIjqy7BI6DRIj/+dwNC2f3w3324BqO9wM4Ai7c2xlAVFxYutWasy8ew1Im5Y5/Y8M9X
drvBNGI8opqTFVLQ8epFwMEQb8U1cKRYl+KuP7AbH/SUQlD/NeWCON5O/6nSvcF67mjS4+aNEqrZ
pzJwmZKkwAYaKDmlAXHwU2K2iDbFCtM+tad4zr5upHpKvgRBh+b5OR1QRiYhrG7yA/Ha7ux6tyBk
AmGL2ikr8KM8cqrAIdY3Gz5h+Kq4wxkNUrK1fPAERlIppWa6tpPJZGo6ORWz45TfpxrjGsaVMq9g
8S0CLL3FjHMeF2a18IVdh8pkHo1BTz5vJnih7KlixzBIc0/SeHXwSImmlPkkg4xwhnKlRxJuLsng
kF63VX0rfPQaYmn5QgyIz8Aux2HnOkd3qyKDli7AFvm7IAnaMv4ZYHTj0VnXZf3Uf6FdHIIqo/CN
jFBLUDPCmCp627G690Y0iboIditnMMgdOFa0w17/DD1aW9B1/J0hAD3+IwUwtQqDnvLF/ehlzhrP
eGmkD9gs3iR2oLXp8w4WS1do4tSC1y6XNY464DWdAzftgqhoFnESu0IQIrp99nj17ds+j7TBWCSq
EUy3ayxTqqTdmY24UvkPLzjbx96QmEmOcYEDmrWn+DND+LjOb/LjcoTg4ao6sHfIM23OCrIsr+8M
ncLLLP/nlRowfbWohobxfYBW3j+BUW3cJCK00MaUzJKDKarPT6FiiJRjMnvxIv0Cd7MZ2/Ho79sn
s0f233wpQwRWwZntzQCALl8cxu7bKPmgnmhuZE9zo2MDZQ0QjKN+F1VgUAOWAYLvnxdAlWu45hBw
/68s1fQHsTYnEznhLckeStzwCcjxmnCtgXkUF6UZQf+gDubyDr9gr+xeP/GtmzqTXbKHjjHRWXn+
FwF5/fevteLeBIo3nmh+f1hBUBJk6y9Xz6MlFA2v7bdCeO0VVU3tr/Y51+pdD9UaTstg1AwtPpAB
+g00kWtcqC23tnWrEp9sICMO9Z/FPWgFtTMoLE13n76jELYrU3zQcHGF0YVqi5uXGJ5H4W4MJUy8
i6wd/Jzo5H8zK1mb9RRFdVJ8m/d3yQFx0QbH3cWlxcIWBsFh2RQysbHVKRXkcIAzIYsXKLm7R+mF
DLKXwoxoDqGpLMnI12/k0AMV/AETybECdISihSBnD/Vo6J5P+99+zNb04Dhc6PhgQcCReHVsPlqi
uo3cdolyFYs5gczWoYF0l6J+rBI1ZG1V3mDNZiP0CafK6R5woPTLZ5P7T3QBn5UsWVUhEXCcndaX
G3a/WTtkJy7ilru5DIVpmEjMpQPhsRpbefXBRDnUqQRz2d/hxTqHqd/I8SOOd2u2DzP9i3mYkkoy
AGYZs6z1lZOU7zVLxpMU7DwPNihFZsx4zcUnQcdxSjCY2FarojglxS/5SQYo6IvKtEg5rg9ldz0r
sFK29WB0qqlyULLLlbSSzOFOFVl0i3JA1Ih51C4vlCgO/vm1vc9WcH9/5v/QuLiZWVltA12tXJvv
XTA9e0LDjNwEMXyofxAVDS+TjPie5Lr0dUVfyKGqrKWMJyPF/ehex5EozZEUPgPGVoZckcCxcxjO
I01hFMhgdNMoAWk/b7GTYjMuR+2wh+9NYO74efCbpNSKpHuMIeLkfzYIZerxc5qT/Z3+tjlCX/KD
Xp/BOsqAF4RUiuQAQoj4oCKEybAkkBa1ssDyyF748V6b0XhgwIA2enZ4Eobu1SKxafGW6GMVbAxn
XFsozBgil0ZcP833q2G4aqIUtymbetY/7pcmeYQ1YSTzTy85dwG80Cq/sl2NF2w8AwLccVbHrwo0
i19wbibOEYUy0SnopuNazMIq4A5RvGWdAdBA2QCgGt+UJm2/eS8dVUssPCj4P4ta0CvZTeXP6J/e
LGv+R/WxLfgmMkVJbLYgmWXB/jZUpMFXpqig04je5a7+rAJ9syzO+Z+RV5cpOtJVEhMR9RTWiT1y
Mq53EFUif6HngfMPgBNN8VjvSpgcbZrZ5Q5f9BUUQxVz6JBzP+enmtEKTwuuSyB2aPF52rDIqkKe
q3rBV8x5cntl88Qxhmck9EBUs1+d2vWKUOMr257Y5EnQ0LR62ieAAR4lYNyJc0ZDQoJCxX3pwITU
FsZEy/pZlFFXt6PILp0GP0TgPkujNCubeBEwyq66MG7RDShsspFJ1A5aGv+1GwM4CwTEhMYYkryj
2jw26uSYy1PDU55stD0BfEHRG7XuSa3hkuTEqM05dXdPGP3H96l2dG2lEFdczzaAqPgdj0Rt1JuG
vOITpgG1HOICULo/XSIqJX8m+A0Mi2NRW/i82M/DTGzEjz0mwhUupAy6lNuynmYXIdOkFjzVoe2r
ac+WrRZM3nUVvPHPejs+wKa7l+A4OEFv9o/luCBOcb6saYzXBDrtCICMCEcqDDrzxXgxA/ZREsPO
0CPoUmA+TsRAWNethc/ci8gHkXd2uvvn1JGRiyGKOjmxwV0fOWgNTvrfw4oS3+SP36cVXtRpTf28
aAckRM3d34gDCQ0CaJj/6+fqYFddbvabs1ZnVahSHsrp/oKgXU32vcas9ylsi9HoVqV4IJp2OPqo
bvyOQyq5imUiyJD+Fh3WO9mWAfQGE+ePYsP7YzJPqs/0IScuQV97UbwgIjow6G4y/fw1SjxusC4r
SRORrl/uOXP8CXY4cRyjzTBW8JCF7PDFXmXWf7sY+2MEISt2XP3UY44maRMUgHubQPIYXlXS8pEL
2h+WbPPajSVnKo/jmb9xDvJkMFlrMYRiAjqK1LVuljLrUnpehVAIfU33HoAgc4U57+0+I1DgVUVh
feedEc4kIrb7NWI7o7RcQCiC3BL8/Oidp6u8Sn6dJ9o0xeOxN+U4fEsIroehcCHF/azdT9ii9Hfc
2fGNOkT6xgOSFJjcQGi4QLzFIbWhKnVOBLfpAj5Q23cY5lKhrbOoYVNBWzuLEJ33pkAmmXZg/RVR
o1DtfmE4iqkQBkUkNkwbg43qZqhSquWO035ueTfasJDXGrGQz/7BlJJhSNcV1SAd3qXLPKy3FwBH
nzrP9cFksQbgKAlLM0D02W9dTcGm3LICxjZUSIbsW68ar2lhOUI3MMKXMR98otxC233+5X0Utazz
mUnW85iTAsKpSWsbw/MnFcx+AKAAMVjlG0cFsoKdGgqM7VKIoUd5dQS8FAaBOBn6edfH//h9F9jr
NJEN4HZ4WPiVvUOxzl4N/DtHvyvVYFekyPsXyDeuVj8K6J6wC+rpzsjeD0B51s3EX0ms9ilqptPH
Tt5CZQVDjQ/ofQ4OmpNaiVQe8RnJMdCI4PveDJKGQoKR+5WGN/hydhHJrnZlXP4kVU4nygl9MW3Q
hC9vbI4VKwWfpWkpmWOPvl/kBdQCpOlsgR0ew9gH02TosZKBdSYGxQQLdHIUZyzymMXr2ZG9lTQH
OU21gjKF++M+KNn+tigLFVlUv7VvMU7bn+EZ3EEkmSq6TMFcxHJBQ487t/UcB9h/zJ9kp7t/QyZe
2agwOO+WvzXu3ezzVcEnqwLL2+LVcrpCNFBfHTSdLUzddOUFmUNuQ+muU+jayHGssiGusQKKbKJO
fuZy5aHgz842/rQQd9+oA68pEMMSTfRcvVv8Y/+2qcQZxS8nz/YNaINA5GFQmEVigcUDYSZk3YKt
xj0DhMf8Qip/dvSnVw05MokbBjVgavvDZOSBktFFIpQqTgxMhP+vtRG9jYQSolwupGcOh6CxJNqL
myBNQSNiDkW7Ps4G9VtO7Fi8I5we5LHJcDn9079iojOlwsllN46Zr8mN3Md/yITc7ZayR8d2EATj
00Jp060gKeAPx9tAGm6YHlObsW3Df7enFhyXRJkc1BvNOGbU/Ru1vFxXcA3VPhJi6QSMU2ek+lzN
uAQELCw+JrgbC87M+7kd2PrdlZQWah5vPF1Xqtrc6fvSqnP8ycjMSnJUMOmEqJ4/r/uGSkEtFQ9z
4YXBIJDNtR1WTBlYENPHgXaTZrJDbQt0ivQ8HnnRTv8S38Lsu9J7OnQ1uFdjnFmGsH++pf5lCqu2
g1hUkkYt4Z0DJ5HUxdkvytvJ7riGmturJ94VrO+dOhurxGtftJ9fUH9hrxgRfJotKdFD6OF8y27w
AZAg9OP+LVLHjSKs5eP7BHq2u1o3KIQ/4Isub3wF3qo9ogIkA6Ix7jZYqzuESQzfHPI5t4sgNq0o
wGlC9MBtUH2Vd9YkzZ6Uc0ObiQVtvpo9XcXDP/aasSZVKjDAy4cNJISCTmWE2/4/nfy3W7k5Ia/a
y9opg5UUNab2y0bMi3F9MmZoCy86XVedWKdpftISE/4eXllVQgmPn7zGemUy4BS6NnBVb6vuRxjA
Si1zFhZLydy95hlxV1boPZ62Big0PEB2km/lwUr4JnyxKpQTSjsDiVjUCm8hIbreunRGk3iIKwQB
kiFQfDRYCdJU9CLTwcTJ3J+AKu1QCcjltTSaIGqB4cHp1cunqge5k3r0GhU2m0p9DyCmCiYZDvfg
2XgiXpMX9DjZ4+K0SA1kaQj8sueO6UMXMA/bD/lTYryhF9kvz4exu5m0kERbn8xkf3z1eT762YGn
iKCdiorqIKYv6DJou9ig2QYhKiVQvN/iFd4sV2FRDlo3hv/B5De1sccnRpAkYxYrHm5my1ORLlT3
wOe+UH3FokfJeUb3FK0G3Ho8KwXa2IvUPd23Spz5ie8lY+HyCNzcYOeOm0FqkrvsNC9LSpBvLWx/
p6YSQmjNdreQej0tin8XYsf8VtOoZGoNlsyr0LMUkUL+oW6NS+kBPo89PKPgqJncbEpdk+jUi7f2
LV9kuqnEiIqL9d1LOxG4GhBt1h9YrcFS1Qz1a+Zjask62Hxq/SBGmsLHLqvZK10HzMx6d/S7GZXS
k0tCm+Ptbm15IxNQkp1GP1wZEsf9kDR3Kd5pZpVAEAhZ+FfBgVq5N2bg0tLXwpVcbcfRw6FWOcgK
4vVsP9ADw/XMvvS97gqPxtRGBZCpfIRMMiymLaou+TMik3ND7i4X78HDIt2G/3ky/WAraMBAEctl
vxykP5I0iVvrTVHQlOIy2j+KtFgYYYSJrgpy1c1CdVpQY9vRcDydSGH+uMTmiwDylaqoS6eXHDTk
v6U5Xyzbz9kG2wrrBGct9pRitYWe6LAHx88H6gDRH+Wkvy3ucdynzZ8vDtDl4opa4FNP4HxxyNpo
KTPSRZQswaYFCoo1p4LRGxZrcxOEs9oFBR2MPycX4bd73Um0aI8oGia9nvrvXTnKwVdBM/g9O6HZ
xBMcpA87Q3CcT5xgF14ppsk5AZaBoXl7Dva86L5ezJ5y+7ka8OoIEOnQFczcY4JFtwnDmwxZwaZH
SX71Z64H71tr2b2pr9d0YKXwczpmhbYPlvOVHeWVcL+sDAzn23Zvsgjz4xd1Z693bLSEke05nSlU
goEq12cwzYXEWzz1qv5XNyzW9EBaknXZp/a7gCvgoJNWkk6dtYKQJc7BFtyR3H1jAsNzRvTDc8dh
LjIQBu34A7tDHkX2ddcrfuzd0uioxyybc06skPehkh5igI/gFxOWcrzjkO7BihuIxu8sh2XlELmk
+YZfTzUxK5Q+Qedr7nVplu9amDBpJtWK/BwtHTYHgXY8jAk6lDeYYitu0uhiQT0nJy0JZdI3l+Qv
wYWk6JPm1+vucPL+Mj2Wn86JOZEdt9t2MRIj1pmhF4GLZnoJhMJecs5J+3s4tZZvRTj8U2dImi3P
ie0ghXHPKMTUZ9245r7Zbkw80LG2j9Xz0WVeEbkR/w5MQR5GOJfUcewSf0rk0cPIz8+Iz9T5d3Wj
RfYC3mQkJJ9Nq7osNBn+dNVt/VQc8bh1rRlZEXvY1WLljEwAEoyDrRU1wl8sCL2VAA7IYKfO0S4e
Oizcq2ijKHQtQsEXOGju+xQWZCfBxb+leXAkW3mJDSCiLF5e68rHBaQEEfAGsJEAt3gDTN0BRWym
U6HZZ1ln5A2QM/HwM3PTwFEK3I0XF9qbOkcgBcJLVAG4m2FNNxM0lE6leoCV6VGD7BP5SgTY/gGX
DWHl4vreUOPw3ZoAUBhEydVa1rHSr//PDESrMgfYVygMiBwQqSZ5XfLDu3+IS7oPW3rg9entymko
KG51pRyoIVdElZYECF+ktYjP87YB4nuXSbUM2zvjpzEzVvNg4h4bGKzfZhEN8I3k7KAf5wMbekYg
xUEWR+R23R+6bkjBY8YmJj6e47cFKGRGdHndC8gkeQP5ILRMTXJZBdksXnkekd8Q4chWiNYWPu/l
5KhG624osbhoYpyWzRi+OCfPRk0zPTlsK3bX0mQlAOLEief2iGjqQWJrutLjqGlvsZgHWohC88tR
CUafHKqJnz8ig/kirgijXQBdTEffhqgQVIdycsMLyU2/9bugIX5GNDaNwalveGGGlS7C1w3rmCKk
y9ldMae0v37n0x8GEjU+M1Ch8PIa2c+PTdP16Zj3+yP0tbRFgN7scuEoYYBwTG3sNOI3PlOdALE9
3EoylYEceRdzJhRwAkSTS83f8a4IUZDdqH9pVhz6AP/FHhcV6Zr0xpGh6cp4zlxPNbWHqxmQyg8y
IOOxhKIosYfpWMJfRYfUu3biZKtGEidlFJkpmMsGYlaFdSsMGl6AzZ16tK11zbPMERvYP/L1NrMi
w5Eo+HKTw9IdaXKhp2U1PiKxUj6Ql5U9YBvdAzcNJ4UBSB+vLQ8+xFxuD4SYPqKTEA/fJSQjUvQi
zb9GgOb95v8rX/nV8jHMPJ4y7IbrgQFRFlYlolmj4+musJxpIjt6zz2GkDfcWnrgy1K9WcqV6L+l
9JSkIbJh9yptpwL6NQdRMla6pSptVUKnhzV2udPcDjsm0iuzedO7fYgsh9VOvdt1jiv++Fqc2i9u
DsS/n+3NYP9r+QIx5VGiGkvZPW4TlU/+P+YYAGBLzVPrlL/vm+khzA20NPN2D9nCpsD+HkUY8D4/
NRZ7j8Z7QdytJ5TdevEklJE6gkaqrg4APng5mLo7ctMbDteye/v1sgUyBOLt7lOQfSiOkwPsvNoK
nQbrOxCj7KrVueYRVa5Zo7e8I9Mhv9AVOwlzfxD1sd+KUMZz8wL+BJzA8Q1LS6cgxaJBgCRSXYLx
JiMzlEy4mG7NJMtWWqLDDR3/oDnJezKeu9RISvCRSDgt3CfU31SmFn7P7oCUJvH4EmITLzvnITq8
DvYPZmLBmKKxVzsyRwyavYFi829y9v/Kx2OgWVwH80RDQ/rPEFesU6ujGOHs04lrBgWm/YLulZIJ
aJbSVu5Yz3R6aqy3sBRpIin+Ua25MWh8t8d0Xe//ZOOqxhDjKgmdU7BQs5LdK0OYGLR6SvNLN01o
zJAdUG3zkov7NkB/yi28REB9Zu4p72ZHjgOoWtK1TMJpab0w397m7p2cHlswCC8xA0sBE0SC2qfK
YBrmkU3+Sq9FJ/pNk+R+0M6YUmE+AD0jhEtrhFy1HL+v0Q8HZnilQIsNf1blg0l+VAcWkkCceAYm
wtI+isULJYQfeCPaYjf2FgzNB2YS1+4vyFsexifGIsV61l+SbTyfzCAqeX8EISHnz0Hitd7zHpMX
5gxPM/h4/ExbcnkWuC5T4EPzO/jdXjv67R9e9Ba7oZZqm5RgRZ6Ge9FN3gBJs9QvjpnsA/BgKRfq
zTgxlSXJ+UmZYiDNn/R5YcfNnYJ9WK0Hj8XidpBaGBhM8GEWVZZ0MmclQZAJEoCa9rWyhJbhLUFY
PuohFMglb9AxT+bQxFr9TkgpwT5LBIBsLB2uugw51ubKiLtuPLB5SrPU5TDHOxBmWhowR6E3SI0K
BOdEnNvfx8GP1D7XJaQ6q3m7iBAS660gSUC+Oed7ty6XzBOZ5uB93XTI8vI1wXRoRk/wcwmAsxb3
rS4Oy7UiCDXP5pR/fyWE1wk2rrnzsbudAAhenmm9geJLqz10xRW0yQRLNGZfn3oVxv6hgwN/WbZf
a8dYe7ywDR8q2+HWWNHLk3nHxrbPmrveOlF7bBHO2LXK9QTUU+Lnm+cCzU2Yvt4wjOSb5WOOgEMP
6Bbt9iM5E7zGkfoI61JD/fror7bbJqLobkSH4g4JVAm/xly3RYqOdW1878Gp/TkviY8bSAP29dIm
yNqH/dLs/1A7bS/YKN9cLfeptifSjJ1bhG+VtM34z7ndI7Ad1o1EWtczhfRUXNPd/S5DCAirjKaA
lEjy+NuHZ6XWD5Mi3+m1VrkibDCaSsKtHi7FFyOBUIvM7LA1K87SBWMhwERG6w7fv9QPBwGPKysE
JsXoSNAMCbkhfUsqNLZeUwGe0jZtmK1WG6uWotk28CXf5yfWRKHWfdDi7xsfZpzoKsVLLVRko0rL
QgsXC12HpaIb4vESH/kJOJspepkoTYpl12/nzuaSOp5VnlADO+u19z8tAZawve8Q44r9JbwfDXWN
mLafZozTsuLSdNYQNNiegxJr/WVjlNIps5izVK+nKaQpfm7LGx/PjYRvZm6xn2ouL7LZwJIGg46i
OGXHGruAolDnDiKmvRhZJuxQCxy+aebSHocqHF5eHuNzF0+L1FAeNSRMzWwboymUmAZFpTZXnvnX
e/xEJtomx8L9yCGQ0SISg+F2UqZwtIzkUejNTQ2PJHrcgDAHoO57oKKKSUMG7SlCNQsEOJdlJa/z
7mlaO2IPgGgaBwP6MSSkKltt2pGK/Rdc1lOdfyyVZDZayM4dfmIgDD7TytS5fFpEW48xUb+CtxML
/lQtZDWTnUCcCbbesX4Fp1uLQk0Q2S/JUBkysrwudTKHlMextPA20gmBGIeYoDwAoUxukeFAck3v
aOPBMxtSogj9LXu5JYHlrWeFeFyAPH12RXCnUBkVA9LUyGT+uDP1OgeJ8FbABCdUrJY0JASLrN76
Dkog+gJniJWSVp/RQw+vgL+yetE88Nfn4O0jHBuQzFlIBIxLDb3996OZFNpGDkN6JlMF8yuTUWqB
fM9LpSoptBRWMKVH0SrMXoUxb5Bc0Ux9uXCNGAfhXqpBp44X+FHYjxVQIw6nd7UgTWE8yYUx3KH/
IX1J4VXwf8BwwlaD2jX+nDO0UlazQuu4B/u944C7nGmBlxJfA/kNYMmOVK/Poi7xkHPxAmtdz+7L
pFVHwjZCtoNEI3Dxen9o+RZ322jOw6iFtxUOcg/s7U+Ul/c/Zzsyi65I/flpLp4VVZK8d6LSwBWM
reRMLJ47d67JsOT7JyRQHDgOpInYN8Q9Q9PF02dNCTWc/Rhh4mHdJF3I3B+K86d3XxgmlHXdle2E
NPxWwtwNRcXxDCBLCmo5+KD+UZbH+hO9Qy3+Pzi/MnNllKt68CbGPtTrprdILk7C6AhB5BjzQrYM
CEUhqn705uXgqoTvCxg/SY/DUgHrPgrxyvv3uBbW+meOHORvrIKeTKr3/fhiTuO7lXsD8fKp5zZq
xv3u0Mvrh3qGdz6CSGZXglB0C+NHk7g759Bwg1SwLgjzQhOcUL/LpK1aTL1do3IsQ2VNbzRJkyYS
2XalDQzoWjjbX4yw2+V1mbCoNQxI36vT9PMpnnDv5vZ0VTyPNVTk3B3dmRFhqS1EhITeYKUK+ZR5
WNT9BqRpzZynOUZljWOGsRi7C2SOOgjbFJfr4Dt1TrfOssKQAW/LIDEAR+YGlijr4IxpKJaN7Ebs
Z2xelT7uqT5b+qg6UzNIgH5Tyvc056gePmf3HVq9IFX2ZA8d2BIGqOJlD257iYg5dgyNEFpM1aJn
6YG4VE/oU7rEPG8cGg00IZo4/VUsYPjZcQArBESMS0U0wP2EucohCKKNhkOC8+wYTE7QbYlohQ76
OTOZRjiy7CkmnT5c1jpqnIaScPJYHRUaq8K1vxNSXxyf4izcHkp9dPXxXCL1uyKGJZ94hIQJCgUG
rZYpMLTQrHQLn91JO3jENHZVnVFv5OZ6AACacM1Sxu04F7ASU0jOrRKrB1Iiu9rvhotX2MHMx3Tu
SMFp0TJ7Mz4RMp6x1SYqfyfgfnOSt3BZ3szpX9gxWBWt7Z2vE/iMHK2CywonVlFDbOPneyiCTbP7
PqWTQrP5jop7Bl2L6EVDeNnkEgiBXHoLvHrdbO2P7whxKMKQ7hJJA6nn4gx+PrNYFCRyucQtZU5E
Efk/YfpXE3ZNbJjHifZxCpHY9WN1WkpBiMTrEp80WM8wjWt08K8emg5tjaYfar3Iwp9JLHOTTfnr
KMMElP2jpwpOMKgukJuv4I9axJbOmc2srgBz7yq6Tb7UMR6dzJ9HN3/RCkNFCK20l1EAj+82I79H
T9eHpMiUjK3F1GvfPebV7CQh4OvjmKOYx+FY6SqvPEs6rPLT10vJq76+bDgakbPvU1NQUqfgPeY5
fuXKML8FzjlgaE+6OvjxkL6ysDMFIhww4I7bfJfXopKgDSW5ykBgW6nMOlQCgxBgBo2T2UxKBSdw
4Cx3QAjX2DBernCPVGtcF+m5PWARU9jTzJl8YRQD/DA7DY6GWtZv6FsxkHvcUo4Evq/RNPDMnztz
sMJMFzoyA3y77lsXsvh6bpepGyI2PYAb2y29QW4cfYOXeFWkXSYoDjWtmie3jaUwHgj9MTZN7qSa
CvHO6XvhGKKi7ztWVg6rnNjENNtgEee0rfSiGK2pCXK6nEBJ3vt9QuLQkfoUn4qC0w2TeL2Lv0Pk
zDuGk1x5DlmpnEv4j0VRNHYIuF/HxiPmGd5wz5KscWFdFvNfouVg/xWZpj1V6imVCkzVkhAAHs44
kh1PBzlU2y+QeR6oeOcrIDJDZc2ol3BDvZHaQ6O3YkgaXmRPU3/dhPoEX57BhbBJB26v0TA3LbdL
Puhpje4T6zTTfHroYijrZNrn/Bob18vEz/uVTZmc9I6InDF71VVqm+df4mD8812VvIMXuebOOceU
cz9Mg+gjWJU+Xn3mczU33PSOYSZjC9Wy5IbQ5+4Vn5GEbrTtmDliHnXCorbFuRazClJNoA6bmpl8
lRoPKFPwluF5f5ZyNenSWakFktXj8tx40IosxHN+9UR8DVNJdzBUBqyCKmklUBc71EinUwVWgpUN
daNdMpLSoKQuyczGpncXlUpzK0ZRWyLFKtUpreP65iExnhRTrOhZ58mI2oDSNPJLMBA2b5IJloKb
nxB6plOR5pDASWp/2kBHYSKEuxCs2yIeqjenP7ZNduWEll39B4F+v5wjqtVJvpTtXDkLaDaQRTpX
kguP0NsUBPmjfRWy0PflmE9PosK0fC7/hApW+VSfHqbYbS7Jg+8r7NP0K0B7N7n2OJ9+KAZrie3b
02g4PyuzeG+pT/YgI9NKJ21AS+Cwoq3ofBReNbwmMFX2zR1n/Qh1j4DkTN5orFf2ZzsI02ILqO3f
fl7Vi8Dkq+mzEjg2dZlmphwzuPLw0e3ldNR+wV+gTVRsxXsntDDxNsnYStybrPRkWh1h4LwlNbpH
HCfk4y2XrYNCwAxmohR6pULvdg3iNvf6BJHWUNgdhXu3Z4QC708j5TSf0aTXy5UyyRZ4A/GIJmnR
GycyEFbipWEaZ7zGwWrkITRmZU6f2v1j9u4cIXcr2xEwrV7ABgmb3JS1x3M1s/pEWJIb/O0JZa73
ZABOo/GGodO499zQ3cgFPF4xGK12lQtfWVR0dcC1a9pCOoLmOKEhyCSraJi2kLdRznNmXGi77LNL
wkleIkVq9/OVkFe77NCm2olvsuXC9jIdu2aO9YzzZwlkmuKBelvu3f0zso+k+huRh7mbRDy9dolo
cEce2sy0EBI8vPPiHes/tA9J+N6vsgAPN8tUmNKsxAwLIETCScLNI1uvwSrOAoW4yfPkCUe87KL6
r62tHyCoXR9OCIKgxWMQFQhf9GmCq0I6tqRUAOVwqPqun3+u9BeOyMHm12p0Rudib0OoJcXzuqys
+NMFFy6iMjewTO0UL3wAp98lIkFkz8MtpoiKL1rxO8rPO5Hs5gMnuWEQkEkqy13bOGgWyRXfMjQ4
DD59MMi0aF+oD4nY7IsoVQZ5dEJqMe5RM1YWEpCr3jJq0RKu/BgrInHp/mgAnWGzX25VNDKw5p92
OttYxUQg5+Zepu6EcZ+n84VwfYx5jnG8zK/2UorLUxyo4nNmR14V/bwOijlvX1tCBg5rqkydRf7f
NbqJCLLyZi/6ZgiuWLdG/mAj9jREazhgC2W6g1n5jJCvLHMX4udO2YM3Y0elA7uyg/HtfLNvhkJP
jzP4v74r63jnf00aw2UiclH6BzyFVywbWTUECPeGS8622pNpu7bJLk6pScmXvITtdTO1ia5cvNgy
LR5M1NnA3AAGM/ApHY8fVJnuawo36hGGKrTM19Pth7tXGLgSdZfqG48k5783owBxXwY93XYJhZb9
bWLoa+dBVZoyZb8PzytBtR0Khs5KDj6CqoplPAeSUoQEU2N6UjL0v6AjQutCMZNHfQobg/KbJNlx
wsbGGgxZ20NpMkVNGDjfN34eAIqcbOZwB8pKQQprinYz+7WiCIlrqTYO6COt967n/7lZh8TBNN1E
iCUtd7BZb4Hj6nafuYRW7XQeoZL2+hFUP4nZxQxKvkAPYL/c9i3pimOwLmr1r4uSKCLUHXlhHez5
PrbqtJc8EWV/ZynXaWZWQkckUZ+Irw8+XkzJCAsG2Lh1tCsb51QOY1jlin0BiC5n6Z7KF2mSYke3
KKcbgbBoWQb/jEX4pu1XKAYZive68Q6Qq0NO4JjtYvgsncciT5RxU7mcx2Eag93GSQD4xb9jDIag
G9n43cTcYQ5lvRrjI9PjK5HZne9Odb/d0B71dh2utHeQPIvCX6JMcj9Ldof6/5pEnHpFixPnD8JW
ekHeqOViDwkhC69nWwtQkIcZVqLWGmtgGlfzv11wBj2RkbEsP+FX5Hz53XFOEHW32tswHjk7A+28
5YYqgMpvOak+TQ5tGt9JIt5DeW6jaevI114NZ/DWv/aj1QzqToqQc7xEBYwU3rm/gnq3hih44aM5
tUEmb+q9BHYTveRG+AB04J0QqFAQ2aqQx9tCPUyFi0Ufkd3voU9V0PAMAlI0mUjehiTclPN32EVc
Jo/3gsuLvLebw5c76qk23oJsGyduJ6Hra07hIBwqD+3ySYBwqQerDjFv7UqO2swEoIsk/rVzTML7
JMbkCf0zg/CPKCgKYaUPoIUuo3ZoxeQwVqssvQzxAdcH0zrQZCuRiN8mKwfWZG0cqwq7EM9sZ5DS
KsLY8VkvcadTSwCWfi5SW2kZlQ5WSDfNdI/q65ocYd30GElG2d8yed3KS/GF2eCPLtO8pJ2ln9j7
3B/Nb044V0nycJbkBCoNqP3ye0e6TdPiaV4fujQPvoyuIohR+dGzl7/7GSUcU3BykovSc6+MieZr
opglZdQ48jO9MMI2kWbokVD9RPSvJnrZQ02N64sXTre8qAlYyQLKH3NZJ1YJCi64iSc1mctAa/iW
BYFsXOCleVSz4QPCnfeEhCr7kztMuyKIeoQtBjn/M6fpB/ospb6X6EuM/c5pjPJuxvgYe5VhZyUk
vSBDBfWrcViZEPcCchcHYKS6V8F3N5AvPp2wcHf0WMxWgtsh1hbWxYkM81lJMoWlYBXlis8Empml
MPPqmBphANDSTpsNpIrQ553/XZtXB9UEAp+ZXzHFWFuVaj4tMrY7ADcdOPRCSNWNXelScfxh77Zk
efN8pNem0JDkXcKENFIAtsz82OdZmW0Bvf4fZuXYGdzwHqQMinRg+HXk0dSCw0+VyUdAKgo97km8
3lBq8stGXEIGdWQIT4oCyWt0ZP75kG9ncXYCFxt3ZAY17ZlfRro9NuW4RMtHfllwHiUrFvUD6Uoz
TMqMzdeBdUEqcTVUAkFaSgh31YXqoySxKC65aniw4h3FwNEjC0dpnLah8NDs8jt71vShQ803ZalT
/UP7N5fiwamqkRc7eJx+Up9wlsxBGjibX+MRx9orZP6Dek2SLS7DzAcjtYS0h9O0m7n7Zn3MbAEe
/aunpKnlcMf3VvLb1tlAZIn0rMhIysUwxk2g+Kla4Z2Qsh/P8Jxockr6oAbnttg+xBiarRwTxW10
hYLR+ABFzI1PByAOPQecM2jlO6Fq5pUuV4TXBNtfXo12XQenFf8he6dOvuz+8Lzw2EdwkrnAc12T
dtfKVnOmKXjSCy96WLkchp3oAdZzCiJrTeP261P5KpYV2SjIGVtXOTCF2kJH1Rvc0RdjyaxCbr6g
NkZ18+j1RvUzO9Kl+YjLkEU8Ub9rAW5vjzS+N7KS2uhmaezS+WfUcevNDzF+epTn6BqxyybaIvIZ
XnqFN01pMRKLzGqVYa6ux7V/AFWvEKZitYmphKtUtFgiTy6PhgThgaqJpOJ1c/Cr0MsKso3TqPMc
kXNHALNNq3aBBkNCltAu4uGq/1SVp3t1tsKddn7tifylbBBQyS27v9UV5FG2rnCLype41LgM7vLc
afGRPvArxubnfKs664aK1ir4enH99Ej2YkCeUKmSZ5dM2exKyekKgeZ7nhEpGT55Pi7PeIv0y7zi
2mzK7T65tbNkB77BWJn+mstcOruyBIGcZqHGtQdOaSX+zDAYKobJae4/SesApt1jyyZ/AoQgLTTS
5gzn7BDbfWMrNrklmDUH6VlBNKrlxslSOVOKNnl0nGERC5aQiN9pdHBbKtVpS38dslI3+CTK2+93
ge1PUxre/urZxhwegnNYHqJJ6V2wF9LuxgMbb0Z9d8GFY04Rgy8j4MBjWP3OSgeUcFXFWfSsvOCb
ULxr4y48ZQMEAKRZ+MmdjmDPCpWCIKQ56sAll5Pdrh2uCqIN9Ph+3V9fg4q7/QF10eXQKNxdL71t
W6t9um1PaaPgCHVK1b07yvvWSQtMt5AAmRpPDDQtZpCphaAL6MSxTSAxkP7DE1ktUrmEcPcir9XF
adlR3ZkKhtqWMoPgnmcJ/Agbd8fhcW4qt7Y/eetTTWtCpYQuG7eAyXQPQ1hwBRMZOU7hlfnBUf90
n7USQbvqNiE/4sMds3rBn5D/fV+7yjzlnEBiT2tNj4SF6OHif1sGfsXU3crW3+02mFaFQRAgbwqF
mkes9WRXJGiKJdoLeemcTj8vXpeZXW4tiNElamBRp0zVvKmM9Y0/fLfMenMOiaK+3l4rPJtZYFta
72MnEIU6/185hcKFg3AFQpgFjiDrruZQ5JJPO5NqoZQffcG+xsmXXBbbCHohrKP5VMbZUX9ntFM0
rdjC19jaTunsfj7ODpYFMn7+4bh4HFUzAFgCRm4W2Pmj4zhxco5vhiL0YN22GQObgHg67S1l3DKm
ZuHEHOs/3k4LhXDNt23a+qQiPwNAepVjfS6J2oUDWp9Ky6Nddji+KM0v0voGHjimMDY3xRZt2NBr
a0LrKPgluVgXKgcbRapx5xs+vk1Qhm9gHQKX9hxywYOBkCp7n4ADAiQmJX4t5pZc3t6zoh6K7ZQM
S3+xd4Wan5Y9Vie1PDmjl+30IMGLMNoHb6CZmW7r9TSdgMykzMzZdn6OVL3384UQE/aPHdjYqVWU
vXv5Htm6LWcY4rv5mli1MEc+BsBKenTA/miRk6684yEMjJgIl14mXz1j0+pxCOR+e8vlbqqnBdFA
NXF5JZjgXSBJWHWvefBt+Bf7fBbB5Ygg3PQDYVACTWP7yEHE6UMSRPvtVHOuQypjrTJMae6JZbOP
CTWmbPvP1rw/u5vfTfaXuE45p3lYDdyHeu3RtIVIXSa7gup64kGHuREXeCX2JkYVHbUJvYes2ilH
SImGeH85kz4nbUVhxEHzxiL5K/Yiwk7o2hmaEifuGO1VyTKY605PlCkcVaT0nxNGs9CCm53Yc/NQ
IC9/y/xsll8ASfQFXKvMLLYBiyH/Zh5KmiV/CnvNu7W0Qbh1lFVXazZmvTntcCBBvcUlk5cSUzdx
n7irAVfvqngJ5hd/Uh5ir6KRpw1EkZetyhPASAXKQgrGbeopaYp20pQuiwt26GgWNP0s4nOX5PBX
8BwDwS9G5U7S9u97k9iqMSq5nm3z5HaSG4Aq8OOTL6WlZTBFmEyUr4JJF8ugVLdadcSMEpXw/nZw
o09E9tlZymgSHTT9/8+cXCDZzvGBN/CrZRkqwTQnhsuAoXiWYToXst63yKOXGkOTho4SCnqJ7r5Q
mk0mCLwMi21jkFfLCSkZcd2jUp9qBSfvXo34J2O4u44ZqzfNvRNpymn7MUKenpzpGyZnyMPi12Ni
YDfppu/UM3WCNW+Z1EdMMCDbBkzVcfIZQ7+PXH/uyjlWBoEu5dpQmCj3Db8moSQoeEAeEqrcxKD0
gvKgg3CvIkZIjqCwzs281lIpuWoorqHP9hbRl9Hn4f/GMDvkQFmN0TdhgcavBhfBJA0yptxgju4P
nkPiTbJosdQciCLu5bGx67r0ifJuFLmEakcRQHPUjcTGMY9tC+Pr7+Fd0u6mvwGwZ8O45WT/ChiV
I94benbhyi/FC1fLjYnT6EJe2HVGnP/CvDez0raDagNVEsoc1zBNJjrYVXjsHghDrmIcQi31Gs+8
iZDGcBCHZmIT71IR8vc3ydqClOjlrxAbsL/OkQjmAz/EOQHfo6KBAK8buMRSMReU2n+jRWY7D4AT
kzwvwIOHNxlWIXDqub2kLWT/jV0kNRtN9VefJEoCW6oKxXTMojexPFKfybuLQpdEuvQD0LCSZ9LI
4cl9TbI9wcQ2YTe5C3QjcC1De2YVzLk3+pwKI5QxDfk2I66erIrk8DZn8HbEIbD6tubtNWKy+C44
RtdiyBo+DWfxmOlwDf172xwpS3YTb/8jdvt7+mdtc2oV5m3dRqlWur2FKGSxY4UmgI6CS7YakvSJ
aCq7ayyvZk6xGdjeRSMOlyP1XQ/pr0Vd0WE4rxy9gSKDsz0CtW4XOoXWgVfZoJopJjYdGeMM/wv3
jSLhttF4HgQZz8IuCxq8v3kVOvPBqwMxVIU4wky76nnP0PLXgSiKja9SvyRQRPx89tF56prnoEdb
czXDg/I90/of1mG6xxsYjOT6mKpm4xAWUCMQVB0KczIPOpnhg+8CjvytypxbPE6ymy1Ts6Ay6mdf
ghVteytT65CwxF1OHxRdkHfnW4d3XAM8oKk5B4GttuhP2anrwbeST78678nLmqxr2BEbKPZ7pnA5
5SGKC2+4iIcQjTavjhncHFwPdwPerJEBxWBc9uTJLBjyV/nC9dvpAHJOyUVPjQcLZQAzS1TOgF0H
SKIwnYvO8tbDl0aqKts74wqJfMxRbUlhterZJqPSXpeDvW4jisG1glQKE3WkHp6UCW+KQwowcfbR
4f5O3J3qLalhGLSPCZdK6Hlg0XrgZVsXFQ6ZUUXBaGRk96bwLY7wkjAmvWm66z93MESekwN27n60
/pXOf1BXZtagqdbtizkSVPv8wTLwhq+1KtEskqxiSISqrZDkFWX8Se+X+j0w6BY0Ijx99L6J1eS0
Bh/NK/O2vrvAnTmfSK58No47tu4KRNR0oVl29BjFBebD/c1YDrXOF8RKM0eJPegJSZWNLAZTS+xQ
oLp3Oqsc4JZnQzfAMJzaxL4zJC2d3lMM83Vpayfp8CwzFfdLdNAd5k5WZoPDskeuHdsQ58/LU6LX
Rskn79z86UQUPjRcNw6ohwEVTMl82IlHSfiT9LjFgEqMhHt+Gn6n5iprhs9sOs+dN9AGi7/ktePh
2e6bS89CXQVCPxgeib5c2KzwOxzlQmWjkFHaCl0Bvu4g+ZK8jbeSnkeD8EjnXu+cF6c/Kbjm2x0G
Vjm0tIOBbAevqi3g6MMJf4O7Lky5heRqVt8uzNUC+z/TrJRNX7pJrAbQnEb7x9lYzs60gakV3eXO
LaNlK27Q3rffawgvdvSCNA43fj4PCgqjFfSPBAawsYw4sRRtINVMV+9kFwZnGuaENtiRQg3cOr8i
6ft8IXlQhppNMlbbN9GwkLN0OOYiRnlvNfg74rg5jTe/MCJjFaDox+/g2Db0vDKLx4R5DLgRiHQm
0nRDntbU+JQqLI7fESMtQL9/5404ex7iHVcSZLKchi+fi5Iq4WctRc94yRnX6Q5VNuWJyXlbmMm1
VZEYSl0TIBr98VlyW947s/b8+Wm7sVyOHLM3hFWDD8WDCY4IXGvW6x0VG3obAEwB/GKgtnK9l+JV
Ly7s/GfC6RFF4J78V6jLN2LJewjKWBeOX9YgnEra88asRlpcrKDjacZmlexv1if2rItIbA/z2EfJ
O0413GRIlw2qqp0eCfBjMx7FGDzrStGk0kQVQe4zpGDzWwyPiDDk7Uk0DOmJd2uJlyrn60i7/vl0
86kQk1CiJN3AfLfB8JCwfo/QMUQBsHR22VicpYtHZHmEjC9pqCO7ZPqJ3iZdpY1CeDeeMXkHWMsi
leaW8gVvSHIHUmYapxI605XN83NylLlCLeR2eM2nzhX4eclrWUS4LHCJDAHt7AswIQFTK9N3MFe0
PADFKfzoVc+U32BCHvhF4G6duwsq7Q5ldi7yqoucUE3fxP4TpaMyDt2UTDeakfn5s2D75gkuxSC0
iwo/da8td+eL03mPoNbL4JfsZ8o6RCXLg2corJL4eTcHbOdXJjwagCU0vJap9gp+dKAoaKaptFej
sMf2nyIfAf4W95TVQywv0+GO20hpXD9dsGgqQLpDVZCNX9MZAfD8Md2VrnsPxSKTGqm2UH1w/t1D
z69+ZTUkCY9uvaicdMnbKTxWUPglQ9F69gt4hfPJVPbubV67pAcdEhDz+vFQzB6skx9SvVXKhQ3+
2osI9KgasH5usSsQEJcGwj96IQlShRPPknxDAQncTLj2Bqe3PRAt4Vf9uhc6eIQP2+028MusBAJT
sccY3hFImHMTKfhzJdepWYuMFJ/5pa75NJFssPPW6Ne9nGs7ByVNWGtvZ0u+eELYuo8c0jGB93UJ
2UB0VOSDBJEwXuT3pbwvrfG6oYgWmSaB1609MWkOeUsxlFNZnniCBjbl181hISfZBeAtHXSCDogz
qQMHulbDY5T9TPt2jJcvx5Ox/pk/gwvZfPqjWnQRw14xn/U0p2wX7AMGZsa+dyoh6YHYWueW7G6H
Q3lahKA0Ajd3QNALWqtXp1VooD7KcqlZgD4TnYgaTxGW78hZWVmhSB7y2JO1qWwQTTsZlW1sJnFW
WcAKDWLw2JgjahEDH7QlH7NQTZ3ZjTgV0kMTfUJp5pLWlUNlw99CJt+spC2uYNueMcDwZn/Zi+Kv
MOEyv/4fByBsnR+NK8f5XBvrXUnpWIf8tDH3wWPY+ZMHhQkYFchDtkUequVIwuqngZlgn5+3NIR/
fC7q7PMBgQgJjoc7/7fVSrbnNJ78nqfNxdKXv3UkJC4DdK/17wvwV6NP1SYu9uEzD8J0h297IgXl
UCziVXfJK40l/8uSzy48/lQNc7rSE4CKwp2qbm4ob1xUW3dAaw9uyL64y3eNBo319+0Trak+dVn3
dumNifF/L8IKTnzx8O55IoCrTTBJUdW7UwLAYWkkkgqulvhF8kn5/JGDCDMtm1e6tb8ucow3rGR9
LY3AN8O+1OqZIwP5kms1QoahDTRn7cM5NaoID5XWTjTZqFzLPVpklwjMZ8pPvs5bj8V8LHhnvzGT
aLfuZU+bldXz/awA3iGV+kNqCWSvAKW8Nwv7wRgeNERK5pLOPeLwV5dBPKQlVOWpyOcdW2zLfY6C
fb6od3zG1KCIoiCoilajWbhqCOIUDh1RrRBICUug0FKal8fMUnYjJxeGNcaCdT5Ruc5xs5h/8YKg
EpNERx2G4DxS3Ayo68eSgsbF1xpp1mG6hJ4REUCFAC7B0rJbxXQ9VjQ+AaPpTD/kQO44ik56lfXy
hDqFCEp0VKjt5bfZzmKwyS0BfErDIUnTa3fyC102qBrSJVc9/AkVzdwyV+pQLYENwXo22maaAVYf
4rkui4n8ht7zjwoi8qgalDEXllREvVZbkqq+kiIGrQ7bZ3niaWt5ylaBmpYhch08nwA5YYfHJELJ
ytBFSFClmAfmFxFMjOZb4H3JNm/un6lUAZMZLIV3MeLYTKjuX3lAUPXMqkaVFeDv52V4oW2NHz/7
9/aYghS/xC09l1NgKmvfvnroq2AutY03OB/BjY0/OKH1b9zRc/juQG5/e7tT3exdykZoPTEMoQDv
ZNCeFOpZVKEoawVZrLygi23sZLfV3r7KWjKu7ZGgIkBqV0THN4q/H45bKCjMMn7psTcN4KB+FYB6
kjyvzIhVagqPgDKeu1hTl9+LIq1Xj/hkFrl6yEQH1JcqKox7lkSEEf2wCmRtffWmvLywj0+Zilp3
HGUYFT4aHSPTxaHemMXDt8eNS62qUCS2pHEwBSzXvJ7pRtWlkEWEZ9sG+IcOC/E7Upapgvc6VujL
zCODnccCffhFeFr09DhSXWrshGAJCK/c7/jnWz7MdetMUJyv+eFl75z3arYaiGX89YcTuCEkAyHY
O4rQv7k94t9lKk+4cjL5IFdl9NAyMyQTh/pKmTxay5QMFZ+pzKkCUEg4iszaLFTiynproEqEsIbI
ne+A2pK2qEJ0DQOjSNokeuRohoUKKgYj4wXqytB87FWQJUMaFETpWsdy9t/ez7mi0W4W88QTFu2r
umnnPMtel8rB9IxIoG6MqyKudmsGBCCkq/nJd3WCOTTiP4O90bu+szBKEp9jTXWN51EERXY/ayR7
1JjESKqBdoXRplJB1qT7kuZ4yIo1uhVijpJW4CErNxz2tFmzx44QPzRyX2krKWLJ3DZ6va/9dI/6
pCcRu3wU6DLh3A5vkC71jCI+fpsAbtXsFJcvTrOb4JpVnCRwBuZda5up0bL3bh3ujZ75UqkDNdhp
KorX9LSSo1QrxfwsseQp6pR9BlTI6HPkTordiDZZsC9o3fejnvIjLfDOn6Of9woHbfQ77bc1WPeJ
OQX8z+3YcLz4OZByFJ92bCtVo9CeOjiR6iZSb6aRmKoz3hLvzWt97+pYE8BEChDACnDcf8rtlwb9
sxuaVXQOSk7Bc7fsw2i/p9FpwLFQxkzqmE1Dr4FFAWd0IqQU+5P98FFI3So9aeu9yGC2lpKEb6KZ
rHCB8UacH+Z54yTa2hZiVxCSZ/5jpP02LqVFmUUekJh/dikXHV1lNhvv71B0ecTQlGa2CMJoNrtp
7ONm1I3Ni2DPV6gl+5cnMvYcLRa65eIK9tSiP0UzqQ/se4KJjdlCf3s+RlICEYEgMPp2X1+QKs/f
XbvLIq0HrY1ibflQ3pFdvpTglbGZb8YS+hcf6Fzc5QrGmKbxcF7mLmxpVIFD2dhdGMRgSEvxyjyK
74MdIXu3rs+qOXqxRgDo8DXSGnLVYLXa16vUuF3MDv+EqdzWqW6yrkYCp2awkr0LwCz2aVExkSA9
yNnwhjc8rLXxjlfHjRspiewe98mgjtpWDM/GqENOyXrNY7yGRaZt7cPWCm2BaWeOxSJMNRvYL4Ev
fbMtXmbWHCRU/h4LeO2xmPeJydKtdHYXGxEupsGFcJVppDZBie6zSQmf2kMdrNeJqyD4eo3DDNEa
3Xy7MvGea1nXBTPtuFeCLYmmSi0wdoWKyjJ+qpontcPEcKLX1b00I4SzJipZUcSD8agGrokfafAn
XlwEnrxKJSkCFlrq7eQu0ki3wZW4dnpDpcuDfYO9CSNdTg/TnygYVqA4spgP5R3a5J/AQX+q3FRP
k6jcAeYQW+iYWlJ2NMXeCfcInUs31qDZkKQb+nrMm+tvcakN3wDq4HhtO2N3XzKxox5EeyOXZDZw
6bKLk7TT48sE1OVEULFoeH/23nSQyhxOWW4GVuW1NvDAko0bThbQWyvv/NYY93tIctJW4ZotLAA4
XWWhdalxVlQ7BoueThygBeyL+E0sz3STFRB1sqkt1HdtbLOH97x1M5RjZzThHB5iAxZJqIYYhLKQ
3IBndFVitv1kAf9s/t5RPnvSFyZheigdIj4naVdLMRfO5Z/Qe92167nVS1QinX4/QaARN138pMNH
PEX3adkq4a4r1+RY4dsJDLjKq4lhInkNKevJf420uGYyZgzR0NGJpb3E5yJwZe9kjbU2dp082HrW
MYeQy3LBK7N47BZlY8GhFbSkTZvPiA4TRx1VWDL8RBTwdF7u51EJOZZA4eJxtv2DnQ+3JwOZ4Ydk
13mk4gJAZDyM29nr3zdWZAIXfWW1Wjfv0uXPw97dFaXusoFM9TkKsD/yRac217AzDg5Mi/HsR5dm
va+fYZwiT+Phmfujrwu/JrhRVqV6iWXn+QilJtoC+7Gs5GgXN5nv7jGfdWIynl3Whj+Ezuf7+P9A
m0XFulbCO97NXNNRDHftqQudIZ7zV3RY2BTcLtT1fIfqosylSogxR9fLcOP7hAjnajxo7cistHLm
swjHIDgjeozda07FRPP7GeuwGnhN/v4mTaXqN38u0m53hUvbHlCTX6WDymhRFMte9Yy3PNi/x3zc
G0lmdrivn7ZRR+M/9N3Homl8JRjLvyyJEv6LMZgNlioRiwTvr3HU03q57vVUra+uzxrUJDXOyCHN
sWXndkML1laVGNJQkDqyZeE+yPRgIbeX04IWnKEjQd2LPITsGOkMEUp1YbEW8Wmv3tGO+kHvaqAj
km2HiC0ZfVDfNb5I/cKVrJDf5vAmF+DZX04/fA8I8D/QlSvF1/dpDFozRwA5MmiIH9wpeilICUWs
dDCcRDNZI11hAtzLMsnGiScyH1MV+IX7azxTMu55rsIZrkTCGOQjTvcC+fXAMyRJfxmgXQFA1U/d
GJNlQoaO64zxDdSARiT46a1eseScx7/eenkJTWVPkekhg08bHdExEkEivim/UByMaXyJLSG0YPDh
9bMpVD7AK/s2JbOAsr7W3dLwoOMHQztT6cqBEWCw0dAoRywnQB2Q0G53CA3Qrg/C0IumR3LMnLrp
h34JZMqfcxVP6Lhsay6ygwetAh6lqFHsg36kAqx0HKd+dF0XGqMrzSdB5DKXJTGk+MbdopZqC0Ed
Lpm9kDWZEpgFh0/VvBsSpCY8Z178irhO36Uy1qAqQszyRWgB67Jp/7rxO4hHSvBaH5G49IwsyDsv
S2TD0CBbC9+hxX4KpgXcPV7oKS9HfI4NAE347njlmPEExBbwVV17KfQCAq+shxFCf2X5sjilYD7V
iJWBMl1m3yHceb1Kbo+biH1nDXpwYePQ7cuk+MUcmpbRkN9ysgPUDIjjapf2RgWy8JADeJWGdMvA
y3hDahkVGGNLR7YmkiOyMRWHbHelTxF1+5Vu8GjC9v2ALwMW1gAjyGfe79xUyEifctXJ52aGnJyK
xZCYOx9sS5bwTZTsYoK3GTq4bQKPjmPIxnseI21xUi2CezNVkiZ+/JkDYcG78RJ0O9xy4QfQdfIM
EHfkIaShxQJ/Gx8XQp+qxXBQAOwj94rWNF29ddb26aFiJc5sF7DcOt4k2rLf6gm+RPsWGyYDpPrf
cEmMDhUCP9hTAaQUdysa+6Pxi2dRii5OLFwNNBg2jSVjtZO3C+7VUwdEFYip2x6V1F4+UpT/ECMk
FRjb/F9FdDHV8bVET2tUH1VejNWfSrmqNb6bdJpud66XTPEDHCOIcSg4KpgxWxgY+EsgNRFoIypb
U2n5TFqxrlUgMAkbViDKRFamxibFKmBTe8/SRuP9OCBpRhMJRM0oIX6IDNH15tFC4Wq/fBikkNP7
RgrJ27fSd+xTgE+34J8XxkJHDLaOqgwEP6UPUHdFmtDidjWghjlYoS8SaRfkK3IAMFkIlBQQy5aX
YNh59GjOtAfFgym5qM6DyxIIp6Dqta2pzxmY6qHeN4wPM3BS2wux9+5WpOCbhHoZl6emwdMVVutG
dUQerWK41PcFT7ZHOqRIDWDCv0OQVBt3bnyyn8Y21GWtLaIdd0+6MelqpAUosfMzQSvmGkUSNTBb
2jNu9R1pD35JdsLibNpGdJund15eV3rhFZWca4w85PvRoGc6cS+DKYQP7idKwOcQcZMu8Dt2Cc+Q
8YmkO1wO+/Gm61cuUJJ8jOIsSrPFIzDp8g+N86b66oeGaffVWSrStsoIhxfaqXVMR6IouqJ6NoL9
CimMl5K35GZ4raD+5t5W2LLlpZE+gIj7KHhhnqXvkFfVnU1K0b7hAwviTLX3raDgOXPZ1JIJU/Pa
omcpZax2KBrojOXJFvB7B0QpDTegYCUt9g9lLcVfPNY3y0r5WuxGfNzbxgsfrv8+jihfXk6v5xUe
J8bt9yOdt6XmyrvlmWatfqVfzHo+JtQkx8RQBpu9OkQLcjHnZSgIdhrUzRwkTf7I+SePX8vZTuqN
Fp289RKc1Yaa1HTdsD92TlJ9QpHLInwhRiTUhFfOXk/kGhWZqVOsRY1oj73ofFy1fsl8IySG0Btj
dnnVk03YzXK2r7GKpjicOIP2toBbSM9Hwy7QhnV0HlcsjkE345LuJkCJV+j4gfWke7fhQRAJ3ZtR
vt7fc3vz7MyMp/N8dR5f2KNAOtDM7nmHT3fwuj+kaBSsABuUuG5Ka+4JwcYA5XYWRg3g22ZNP+JU
5ud/oF0sSB885puwwVxBYXu/F6xBWTtdFlK7QEx6QrnBoq8FlhGlV14qGdzoniZk/tx2DaavPAsl
e8CRXCW817/f82N1Tyu9uTTY1pMD26ORoEJv55D0Bev2dqt89dLKOxLsmJlDQ95IcYLoOMe6/QwJ
T/JhQkk6rAwaxmupJehh09a0BzMowyE81iEdeEMkHGgMuFc+csJ3IeX3svrDoQbehfSP0usQFfZ8
WlLcqe4H42lRfRHKlcbBjSYaeNfFzhNEXNlIvIWJGWp7hfz+hy9UbiPR+OeMOhghzqP45AcikjwQ
I2XE8uJ2JDCpRssQEWIFwTUQ9zqa/jDO7oRCtMJIFoifurMtbW8G3k19BVFt6WNs3KdL7tMwU9QY
O4bfGXCynr9lSGToBAXcWvfsGNaLuSZabf6fQdR+ZmSqWFyFht/myxCMjD4+3OomVGyXbBTgyUt/
N57IhV3XjC+IxjUWJoDv8uMwujpy8ACdYrYb5FZxQb+4P3A5ct8cm6FRhdPxaOOl8xQ9lo5p0qbI
+nNDWtlJrr2P+SJLW/HjNBt2adOF1nG8oECXUARVD3lyyeWq6DrezHMa/k0CqVTADw0fdVJias4W
JCg5KgiAq0ZS6Mrk5oc69jDuROMxqhBJ0HOYuhaI1JdfRL87/03A2bcrqgp5luLbTows6cAW1z6M
B5FRatqFnZe/M5WKFM13UaUEjoQCnjlS8Q2ue5ymNQC1QZFOwDuahvG5+MDM8ASibq0TlYZgTpmf
gzKHS+pIYkBFkmpt5ViLOBvmuVfHjaGMEkJP1SxTLhGDDPjOwoCg5R7SxNoCiniHP7bq2teBXHyQ
CfxboUnSLE4hKkAA7RtIbpBI0xsKCiF7z1107Y/3WQVkYCWhXsykpqib8/vG9igPd/pIitqnlcoI
Ox4Q3V8DqJGFO+EKJZQlUb1o+3ZlEW+U0McAUwx5SYL9XpfvE5dH+Uqch6erOAxNHJxadAneWWL/
tLl8zPGE+G7xbAeNnxVbHU4hUUNPSIWUF2IE4MmHdZE2WZw5Z4FTiRnJVo65vUa8uKdaEr1MHSoo
Fij/unKI5uDKPwj9coRW8bzg7Ywok7lCMmOqz4AhLNJZ7rU4U5YNB3NcG3sPZ/WhaBQm/XjEcF5S
qFtp9fENKORZTW7TKGt9BOv+0E3rofT3ExhIJV+xYq99P/C0j9KKdN0MtStpyRAHpoYtfo9pWMbm
UCtcQP9sMdhbtLqCQX7Rto+MgGd7HVcCLRo0pilU05MZrW852upXtOIUwStCaOXpfGOjpODMBQdw
dFXND6zQEHvULFmtMj97eEFt1Zqupld1Le5ao5pOD/P1yx0rwUzyniSqLaXFkVUTKk+AweJ4JRFe
TNopuejtOSCnoLIwuuIQnp0lFUr2IxjBd2oLip3lrQRd/izmeuKRA5Sfa96ze/Gy41wQKfFLxf1u
aO24lLwERhkWeSfy9a4SojhvH6aSMWc1GYwuCC3fLrz1nVDDsZGV31Pq5YYZllVzVW3VgOwWfC6f
o0YbyxN9E0pBoMaCBPLgyfRRzJEBON7Kps3vR0slwsui9Br33KnkNEXtCGgheBzIZ6I2QzwjnNI1
+ulCU3oY3o1Uw88QyZ4657QjxBXY/T6i5nFDdHs2XxG523YpurgKpYWEVFLcBdNIS0P21d7Yy2e5
EK7BzJPW93Wqxph0vy1IuGtJVA5OYZf+KEQyYPNxw53emuMfaESMAOBXIAcjohTTJgmNZ/fgwWLK
CbERFxU2TX0J1y9os/CXBJI8p1MVuPA3YhjKFikz/2vElm1hSAI8/qCLOLqI9BQjrRlLXynVFNpR
GHCqs7XMrEnSn6H489j8/B1ivu8w+F+1zRjI5N+F8jcpRnLhrTnx+yB/oXdbwST7fyMC00/XUzew
r/eRrtmnDzG+m03NO9EX6eDduIxvpSbUvbadahjof8N9hQ90t+8j+UnY+ekVh1eg4UBhYOoLMb0K
3J1MBNFq6fslNoR9mrkmL7OL+dDz0Xix2dVXayjuKYYBx9ei1ba348PWLM/hpYyR8TO3PHaSLZf9
450JJrtSOfiA7KFzviiwU3Bm9bc/6AHAIc/E4u+INSdzXICwn357M6Sjq2bxudXuX3Wr1+39R3RR
hOUZffjNhDRdI5HTNsCcY/GWpBgvDiRD3s2g/L+M0OIKixD4O0KIDsbhR7a3UX8ehKFd0xjRYy9K
bKYtQ6w4hdxoI9GLKz9c1+xtoJ+ajIu3VrkfdNurHj+YJMNuZe7PCbaXICjBprxAlQ7KETEG75WO
dqYpBqb0ebhHcZe6AOD83ojlbTzvrXFfPwHR1CB4k9vLTLAd9yxw+fA71ogrV4z2mdHON+uOJ5DS
F2VIVXfpVZW6YsPAbqoChrr/Jy60Esdon80SD0bVpZezNDJZpemdmpiGuQKBxB4N/Z0JILSeh5N1
FEsxQmqBR4pK4jQehmmCzLoP/GQIIwGybRFBqE7xsfB3oiOA8cHvse4eTYEfCgSh9bKitjxhsOS+
MjVxes/ggug4Tk3ubMRPVkc2ijENPVmtTe2pZYVe3NjJyHIZX3bIy/apEs+ckL2mH6dmoNdyNodm
PKRpUjs2yN3Rm+xCocz0gUXI0ymEFBs1fgPz/tD9479yf4BqMcGdxMC/KFdF3PDJbcPynRHpC26A
MUr6yB8OigYmH8W0zrgp2WH8S4ml+Xei16d+a2EJFCUnG2IOrKeVGgSiVQfUV/Y21obVOMguj8yh
YQVVkJKgZd7iVGQOS0KMreZEcxwuHZxkNzEHM++qc56yFbbDzHGM/Uhdf0p5ZOs0JqCniRDprQQM
vj6FKpJ5KovJNmw+Xlea1mrlC0eihEvwg0JIikrXUMveqABrfhINxTtkRnquxHWLQKta9/l2mFOV
pY8TYoxm9j7GNv1LWhvVRLpe31OpV4bAUNyP5dsX7rDu6dfIlo5ZJVUKpzsccF6TXTZM7BcPZzDv
+wIcGv5OWQyuEB4EwXqIXIpKs8fMogz2oCj4ReM2P4y6vkYHEMXml6+0vr6YbtYCmqXikJduO17y
p1IVS8rCoHBvN8HKJILEVm3NB93wpyRHiTJ1e8/u3NYZLf39MbU387m8z13kE41IbqRFJ394Sssi
8s9psNtkheG9Oqzv3jCkg9KpEx25D7dn99qhkWtN1dPk64fkrOmBdqPtSAPk/E6sXLD4RKxxJ1qU
1GRa9wdwObFZNB68tpSi8zvG47s0eG8kfNetgNgZRLR2pIfTLZGJiaYmsFApViFzBzXLhbO8OKbd
ufZVEeHF5gntw3qcUoz6nKEXIRB50+HFFqsJgpoeJrSoaZrrD9M5dT+cm4qTD/G8AtBswIaMg6lY
W88FMBVvHCRDyJWpb51O82Y9G4CtWyBAgmEkjCmOEl7RHlJVguVYsrP7nyzsRSHHLkpiDFCYhDRi
sglm5zb6+I4+CpzYTag1XhGtdj7/2kqq6CxEYdv5U8W9QT/FJRspGiPVQPZfyv51CB874oxu/M5G
mXPEMPBF20z14iieKRIEc6UCkvPSFIg1zFe2+dW+4J075Yn2t1kSV7vgWm6xqHVfy7cu3EpZ5jV3
SiLuZ1NaEdB66uOsPUMzdDieycKAAAIYn/GWLacP6F4pAIsbSu1DauEyNvqa3koY3pgR2wckdJHF
F3zhHnN7YAHYaq7IEwHxzdLv//WYLVKo2CUPSLOF5knbc6HVAZnP/LjcHeaVPguxnzHL26+HfEj+
DJqaETY9GVr9sj4xPh2CCMtyrNq6nT6147X02J6CshnSomqdU2BNWaM45LONGwggtAk0J2gGoXo1
vZZWNUOERFkbY+mfIGjVLUqHOoyoRIkWTvvUV5QxOKLH6HepoN3e7+ls4upfT8hojfOasIFNV4vb
eSqg/HHN6cZEihUNeH63gJCj4G0lM4qau+RVt0+eX3/ODRQk7MmAxgmU21TDfw/DsQio/kFHxS5k
ewvM50ovz0Hrttco1ny2VTNdYlSw1zXv9g6F6qs7v9v36xAZDWHJd3NP9umAuMdNKn09WLtCc/ix
cyBKc6ZWh0G/kV76cqxWVVW5gbUVJ+N5eE10QCsMpRs34KpI+wpHKZPlHH6xl5+F1VOMsmmtaE+5
h7xr6VkSWIZYKgkThNDT1neaN5M6hzayJudAM+uJESBb0lLi1+WobnAp7V/JXH1ConSLW55boOso
umY17YOu3TfLmQk50WO/NjRgfvucBtO1UuDhsk69k7b/4G5g+ezHIPEsccQ/JFH7SW/Oz6rQ//qQ
vpIwtkXzo2K9QMhAzD97IAr8OGP3tQWpgEthuXRatE3Xly6dUREtp7ysHQEwvju1aZBY37Y+u1Mc
3BTkjYCAoqZcQMAnlCeEH1pCbuY+0qqWlpCtuiY71POYkvDEwkNFg0hHCEvMr0Ff87bwN/+OgVBP
IfZAGLadC/gbA5iKO9AGKXDMAMFCyrWSNoyU+mE04MzV30i24fbmXhBy820A6AQGkwmtbM8bLgMt
Uwgi4m6uWip9DPO/YMmgfRxRYA/mCelkZLEL2XW5aiPIaH4oNdcBzojUmG4h2bAF/uOxHqmL/2A5
f5gRyCDprpGKsKpEH/L8+Gemuew8DfG+M9pz5c1HzvSlx1MjLk0W0AxseBLKWGOjk8A1D5qqmi8c
Byc3/z0a15s0suOVIIpAA+Pa778y6mD5KvGVTcz9vc3VQT6XhIaFLNpbxRKFksdoX3oKEBmzE95Z
Rfxc7XFPr7r+goKoFYglizBahbZUfxNY0gr4e9gk+kXLCcV7Dbarf1U90P4PdSUqznM5wvHjQuCG
PVoxy6QrSEWu3zhlRRiNy6EAMOHFiZAexpJr2bTvPOjsm9xSIamj0q9Yg7kBbX3lhaNWPKmwvGqf
h8YnezAslPMueGQ2kyCaM7QBJXK2Au11PO/y57vwRey3Vx7vqQxzF8WCKDWt4EWbeVKfxch5TjaP
DzZ7EJsBcJG/cYhGIuJmSqA1bfjk7HkYNmPVS4/jp4jJkTH/OMnYOh0bGKKPHzGz6b6C2G7KRtpK
MpBQA6IRCp3kYwNJtrBq2/6sU/gBVxBuySASBYz17qP9nopOJJVWhF/CBoWAW7A/ULd1Mz4DWoRl
GioUd/fsMWszFC+a+ENq8SeRePLHvP6LomEWhgiROdMvlvloZ885O8ImzT5NjsgtvsXBduufeJjb
jrNrgTxSzU928GRdI7wVQXdepoVcjMalUTiZ8FScvSfg1rvL8AqA6f+zpkDyU8Fj/cuXWmUN/Ou7
VQtzCs4T3w5iyqx8/p84nS5kzJ+b0vspR9X2r6Wz9ouYv+Dn+Qo3tTOdWU4oK0nR9sP34ulwYDm1
mnu3Uet1tPrmycYKXMZ1xmiG6jKBXquJuFZoKDpKTUFMZ5lOnwYGdtGcofOuB5ZGuiD66HNY2Ih6
Fy32YMu/RKIa0Cqbw0IJw0YRDGBigQk39+wmZVcst9eoXnyaE7x0s/zyYHtR42KhoxS0WgDMNZLc
xnoTh4G/KvjsrYqEBLiaaFLqBpmbHCslYta8NlHApZhC/ptjp6bgkwFNz6iXJuKuGMH6v65hvoKf
tOtUgGRAmg30paTaJrjFjng7Vcj/tdNT3Y9fpj0KWBcVbRcXclEFx387fiJGOyCsf1Y64tK0xVeL
qLTRQ8bbehlzCwXwKZ808LTxo2D3nq2cCMYU5ZJMtCJRCWx8u7q684CDfVtbkV434aVLZNCq44IV
2IcaYLbEuOSd6oBEI/ejJ/G8F/Zom4seHk9Oap/jscECjfwFU7eBZFqdOEr+epi8/bSmLQr7TkX+
UlQ8ZSJQAgsHMNdL8CtikiC5pRRMTxF8MrGEEE0b570N0JlutLTAdGbmpHkLwyucJ67X0buf5ZlK
a3NJkuw9zXL1YBYNQfZwAggCgJbuANsGm7L9HKfpCXJwD3//+1AEInjzWmbwZIaNbgWexWBtF0sI
bEF1aJ5CMABGxlFgxDg4Vz9qTCQnBjLMJZB7ffdcRDMWM5kzsn7CS0/L1ibJThHvBKWw54eH4QnJ
tB/3tQTPriStAHrg4YwwbLtgRLtLitdLTrLaNFnmIfW/Tnm1uDAEMFOFFXNQRYtwwkCqajsCsIP2
RlzNzNzw/0V20hFfuRMEemhrHRcX84mXxdBo/hNyfHvr/5td5gSHu8ajBwiau5kX8odNuAhV7rpk
nWUHVsmHQjunhs7jQr+8GWMnwm7r4ERs3syxCXTPvF6PPuijGMfHtdvQnzypOzweog4Tsb3k+qtn
VtQKO0pMG9knar0lEgfEH9O04/3+etsh7oieeBS73ZPIRov2T1jyX01wU6yuzR42Fr+hcWHiwi9E
/tZa1ksVhi7+Wr+1qwwE6hzWmlgm3zhRj0XbxxtrdJbu8/aDn7eDP20G23KTmNVGvczfeLviITfQ
oN7c07ikiRSGk2sNqQ3LGK1uLlk6l2obj5JT34q7lKLp3ywRlSHAjnjx/5NamQydviMopPN5pDse
Y63eJmHS55Jkkb3p/6Usal35B9p7IZYQOet805QT4xHS4V3gGvycJC1d2f8bKJ56MfhsCiflvNIj
N8FH3+/IBiXSqL/EiCK5CWpeTcrgbT3R/tV4hLoIqlVyRyLmpxcwLeoKJdHFpQIRR8g2J3kb465Z
d5wmaeVINuJlCJSTxlQoCOIHVipNdjYLPzp4IyM9bVhT/eIipZxNfbNznXMD6xMTQF8mM8LV5UhC
ttbQuuDoYtgTLeVno+UCZcOKR1ZsIn9jwX1zWSY71h0YO/ssaCFQdn0fD4kXTmK0DNGLnf5ZXETl
MgORMXjYzGPCSFNhNvn5+oKczbtuLrIvu9qXS/mqR97t5Zo1bO72CGOZxsRuTRoiOCSWuhq81oDo
C7+dKbWGm987PlSbnJgTV//hBGcklgVgDJQdcIIXWZb39YsPCoKK4UVLmq6t1z8byuBS3bO9Hz8E
TXfRA/QG7sROzsWko2BtLRtUtgdS8WWIDFlOjX09oApKoFEnIuAUJxP0nRV5uYmTpaGhJAFnk9oG
b91OGC1mzaB+GvVj5Od2vESArhMHOwh/8FVW6auo6I1Muz5Qd6MylX2YHLJkjam84a17BfiofpKx
TStqzB8V36DXo86XcfQy02XiBzYLjm9YTXeS6vCX1F7xgEjUgKQnPFc2+qTcp0R/6XEq2yHJ+mfc
CwMrgzN775NvIbq6QfOIq64Xq6UoMBppKRyae4mFRGaQhnvZ2aFxJEugF152nKUkYzXlqfFAy5CH
cuxSATOpFnOOHC/MQvNZjbje1Auq300RxKXUm1d9iTs6Cv5XVZgEWFL+IfkJZ0rPekPY9IW3/zK3
bBChQSz7mJuyksKKkFzN50E+TxQCmW8BPsu+aOM/0ZhL1lFWx+v9w/ACVhnwHUpclBEBepg6U7QA
2QGmXm79mZleA5R4m32fchalAHUekptfhOX8YheTqn+k65IP5dxDjEfNqCzE5CvqIhdHqDfCuiaY
WdlcgME3U/eJGAvF2cdOOJk5UKLCYzne4w6pRL1NLpsiwEMGWJkNg2cuPYiuXiBcxihsB0eAtmQE
jGStt2vWR/Bt6C9mtOogQm+4tnp/ZQeBRNNdsjQLs7mfavp5tZwvPmi6sOGdhfQuYMvsfF8QtHG9
EYPqSxE2rMxwejvGyak3KXAcqWRuSEbl02UlzimB2/5gi/jp6iiJYIYv2KHNNiaZ4fFnMWPhoEFS
hpHkUlB0x2I3K8S9E5KnmNo8lIVm+WPxI7WMBK/lW14X61kxOgahsdo6pbt30kQgsqzPq6yIgH3a
kIM9wymeSagv/WfExKW2MvW0nYTgWV+aTzfBtqCDzLQMagp7EtLcRDgzBp1VIpbD07FShV9owP/h
gB7DAn+7sHwVoz783IPkozaaMOMGMdfprlyvOWZQrY2IfufKeHYnsa1bHBbG3aeTKxRiV8cOrWxE
YfcghEDNjLquvl98nwEeODch+GKoyzox6MntTeHHZO4x8zeeME+dCpMPa8GYkiLZV7CTqgwvEmSC
pgo8w5mtrbh85YgX3/CwnRZJJtGi4m7qOzzhhGmf+Rv6/Q+VUl38/dV/yR25nZV2F6vXCd7xatUW
NOl5P9fa+X9djSWW7cTaDo3eie/5nvRMBbpQc/8pBYCxSC7FIx3JT5cb29KDm5yMHrZdLrD6d+0a
pjjiqPbPhKQ83lAFT9iDThQXQ4/R1AiVuufMSc2X6lnffbDbgbQYEU6FFLWkjH69YPjHIpEtOZzv
wejglzWvXL3IBGBMk8o+/n/u8UO5Jv+Lqz8jcQQyWVDKfW0CUZDhiv1gS+dOFhW/ECpWz1iyoBAd
zwmppkmHg4LXsgIWreZ9na8IXP9k+lNgwpsYn1K7lJKe89hgVXWzsW+3JXseusJZxtaghNkjnc1y
PrNysm9SX/LUQSVGepWUqmGYjNfuR+VHR1gSmHUPbB2B6k2VXNLDxfGKWmSkJ7Auf+s6Luw95pNa
h3J9yxj3Lqn0AC31J9ZTUE8vRwxJoD/jjASBFFFJ6SFIO9mzayCwhYBuURcJLRtcZaqkeCp3D7qz
F979ioqhOv59oUOBw532Kt4KRkDcE23unByqmuFsZAXr2AMEOXqoH2M9XPOZN4q/MNva/PyQHF9O
80+qHmkHL6SP82ExieEgXnbZYt2OXn5aEtPHHj4eenAdIYpcKeTL7yNZQqSvsraEQJqAweSaGBDK
vAPbYyddXFx+nVh5G4ISjPNrVtOQXTkxtOS8nCB1xhuiCnfUM/vrrajjnV7u0vxaTwSEmJkndilk
UVBDsbrbo17k4I8Mim+/mVQ1MhkJlyeaNcQS+RNG9ahD4g/7kLHh/GjZW+cuHqbrDh0gjn07W88Z
I1ewRbmxUirl+9mm60cD4Og9TIXPsjsU2i16pLKjSb5Upd+Jo2BNsTl16q9Qz/wOvyodNKyDcwLZ
TIsAggB2gvkutIBlARwAMFsYPwhQv15tkkLzR6cDUL/6Qh6TP1wfoZ5MI3DyFd6YNTxZIiaRFwH6
x7wTM0ELtvL36gAtS8qPOpmaVOvZPLgepjRhf9sdQzXwkGPAZxxvzaXwtStqAoz1PWKcHbKzwCWn
Mh2+tvZyhy1dLHvTr7NEXBavmUJcCNpeVg57YM31l/3gRrCfdDkxb8voyRcOHEhBkVUkR2zLLVDT
NUddytnRgGJsSN3sxJ44cuxSktUenq5JFScAPKZVFYqgMXdmRPQyaQKc1rIddGTmLqDLrGqr2Ymm
wwXGjgurDLSbjFMUUjtL9LFeypATh0JC01xO1/qz1voWiagGqJPLnAxtMu6VMye2eoBv6r+YlhZL
/x86KCHbJ71Fx2rtolCPcitB0glWyTckcm89dTiUGpm18wEbKdl52prlWbi6dKABW197rGPHEweP
wqv9vAE7vtD0O6cwFXW41Z7qOll3/YFUG97l5uk+0ccusmKCFTYCk1Q0sW6hT1bPZEtTCa15J8B5
lr8+up2oRjDNFufmbicnFdVeKKzPgX9kVWg9cRn6XtUy4N25AjOU9/4qTMLScgncQDBn5V1Rubd1
JtDJQwDk5yISn4Vzr2a5JYVD+7uM7jN2FHdThsiT0TxZ2kdy0iyGHen3E8MVd5oRVZ2uUk1ZqIf4
nLzTaX4maXNsPwF+Wvj1T2eUNdlHkthu5rekZQSykCRv4SuFhbhFX/1QhVmyDB8SdVrWzZ40UUxR
NOSNABcHX6/Ir4dOa1KpEXNlxsYEb2+92yd6NGyPtQnrRMtJTV0MbR/kwAAiUD/VWZ5S1Vh37UfO
JuoSYtpK+ADhrY5QwHmeibbB5zvwPQuhVkHD203JGR4lMRv8hR6V/uxYpsauer8pRCSPhi9EdesK
uioEgaivmuwCQsPceEVIKtcTVbsPHw42jygnVk60EnlhF3BTSKJFmvwx04qla/uRodSD+Z3+dl/R
8NWojrA+afTV/2p7Ww/Zk3nv1r6gtXCYzKXOW5XSTycRWYcTMYg0vod/UKpwQ9QNH2uUMTl6UADh
NCkvJPTivK4XYYZ37tuDo2nz7oCb680UkKyNbzP91ukXGOWKMiO3lesZl9BtWW2aDGxbx0Kyd8Qe
AMVLf1SWoFfujiiAdsXHTUr5Hqkep6aTx9/3ht7l8fdwQT8oBbNojycHS3S0JtJzpjC68uQP4KwA
UAap5UpEsZNIXMZ1EBdflSSuil/R1OgxA/469NtBk5yAGOpZIQ35CcvqTbZvZT3iDz3ksjaTU8Ha
biig9Ev0KUkXpCJPBGTDd1x4inf95RbQUdjmfELo6gyB2KRiNXJLqSrsbSDRNks5WJiUk2TXoZut
u1nxJpQlXevSurozWl1wHxwQ3S1QeaJXR7U1obmpRH1acsbgazfbrKAmZtEAftIrlmvPDMLU/f1u
BGdZLr5uNILYa3L3wRoiGUZr73cA5lbNHrEsF7cjrIAEv4UZ2xRWsI9GebSYCUcnWGcZe8gd3EFU
Rd9YyH262a4aucbGDIdVZCOJCt/Z1I2zhSpaByjW4FlSy6qvC/bI2i7pBsencYBqdoqVXOopZ03r
W/rYqY6XDhRjy0UTO0cxr1x6Q1fHreWweOkXzSIlVm7scgfk5oyNHLCLgR1uuPxPGvOec8MW1e7Z
5mNLl0lwkZ85b6VFaxtriXlro3gh9srEjHQJoT+1orNT6JKD7ETB3yUqJJwo0MKiPv2MosTE+LUH
8oVABguOF7Xcy91mOiEE0peg/8sFe9NTKgEKsWfrzXD6RX1UvNXTNtcJh9zC3BJ+S72KYB1TszEd
zphruIvjUp+fU+zpV1tHGsLHZNAMgV4ojsYyXj1hbwquMM21gmJIJHJb1jjlHHmaa39RlyHsOpH2
Vu2uzipBVG8ymf0QxWz5NFGg2lksD/6BdLZOrnELiC8d5z/iBxedBr8+e01tp71WFXGq4b3XXKkL
jtGYBlPZBhKMXDKVkaMKa19BQidgcBNLiX9DIXqknMWTqN+kFaFNROOY25IvteC7F758fnTjSorh
jXssyQmnLKQ9A5GCvmyKMXbZsCpMrtEb4CxRcNl0O5fo2BQuAj7w18uZRH0naTdy3Sm3aKB4d0F/
bu4QdrBjRsbDx8FpTA3727cokKQq48ug/vqfeXntXpx9qgiaSKNrghmHAXeoaQb7vPMMPO50dhoy
99rfDG0807Toozg3Loa5bb9t/K/SgxN4fspSjAlcEkLu1Jvro+i23jhJOBgcFqBbQati96XvT2V+
iycNAC1PywBN4TLW08kbjZa/CxfjLQ55Zonf5JGh1dZCOuDfMHD81hmN370jNBX1v11uk+e8ndxj
Cbofghc9I8apjZIDN09MOHguqg313YFM45QM9ZGrt1ndaTFw04wyZ+TWMoSb7udO9JRq9HZs7KCH
oz84tsCkt+sHoJXJ48rXLWdv7ztvab3uldZoZuwvhnSu2foa1pULT2/tQi8OatU92oeBSD9Uzg/Y
gLGx77VS5Y4HIettu9tmPXTXuiZIi6yQykda8sjhPJp27HeZYQiP7XUTZbM4R/SmJjYi0sh9d5/w
toHzgTuCRRl51WLmXfeHhjCgRKrizUd11+i0NadO1SJwVFgmypeLCc+8UiA5IgE8vDSVVztQ67/G
RwZFZTy1mDjwdReVE+97zm/QfHHOmzZ8A+GSIGrR2smz69MuvD/K7doOkLqZPqljK6LObBoFfFLC
OMWoXt1XDk0tIBi/v3hItJEu0CPxQ1BSsac1HzQpQkqKacDsbyzup4e/VmPKNBheYntsUflpMpno
fBnj1Au0vUYfE7fAJavjc8DJ44TzVnX8NX53yo3bBNGRrNOyOhN8js7DJAc4V9BPZFaUQtKfl9MA
+31N7hHCSoAeNCNhLMkaBNekQa6P/YANgV7tRooof5lB+K1VL00ZaI2w6Pbw1h8loaxjMAVdvZ/w
l6tG/7mQv7juhbAFYuuHMx/8RRYUqiqZQT1f7eGH++6X9aEJQHzwNKGyzbvJ8ltYJi02YEZKlNIN
B/FNUFlD0tatFT9oVgb1+8rKNCvbIj7R3Hd8fFaHjv3GTnlbNIqOOn7oMZ0q4h1iO6sYdRV4LH8v
J7kx4Riv8t7j9h8ghzN/B0GD1K9kbZPuNzvazPB4mP6ljIDKOk/EW0Aduy5A0fK7eWWrGaRvBqLw
MM2Ndi84Clokh0bsVkZYPEq3vildtbooahK+XpKvi7naFfI0Dyh4RR4FUADYsj9C+XwbQgb7J+JX
oYq19o1btX0ABWqm1B8c22VVQDEMJUKkAaOBqRWS1gcoQ8c3bKV2cJbWDmgVjDkRjPRk3JkzirwK
ngX/K9SjBEMFTLeoIddgLDaNLzaiKMZuhjx9fyDAeFrRbNOnGQb0SOG4wMlbPNqChCf+Qk9ZN4j9
qYI4lNoCdfjkY4k8YHZ5rhSI32+Up6j3UQN20OmfT+s6uS7Jf5tgfIQd+dcAs54Xh4U/lAu2pZ/Y
E6gPv40X54kfwjDvHFoh2LOwQmRN7WMGBRbehLSPTX7/v/slBnBZGyfdVo0MbRCwRQziM4CdjsLs
Gs6jb9ZTQ9n2hWsVBFNveXsYk1d6BlJfz7PMsFZwxWC7RhGm0I2ENKUuZFRxs+pSLAHyM1C2xSNB
5wGzkPdTDf7RnGYo1Z5rdbw2OeXKOObxQ5UYp1+59wY7hpbboYE6MmRjuJhZ0v7J4r1Kr2DekenX
JgHeT2TFqMzVDhbyfN3akTzgvs8YJ9WEAGEl2F3cu/ruez8AJZkSnzNFwrmPfRFXAPYCymtbAVQs
1dMF2i1ZwibFzFxsEYCod/NKuvbfUfjVJu+v2QmhVuhP5NKADUHwmHa5cnhhzZ+Li1DEGpOhLkGC
TjA31eWkpk8Z5at4fzQcajHSm6yUPNDsGjA/VDU19iAuuo9IqpsGpiQGZn93CSotAZBGJmMMN/+7
JYLxh71x6OnFBaqdlypmcMxE2JWIqWk9KgT1ItHGc9SIYn21ZuCKDEbtIWSJxttUuDIb56adDzsN
1hJvM8XBB88f7vkh11G7Z/O2HEuel47FrqF5vnTxVdCJxGL+KgkWb4UJYNDAgp0tsHZepOXYWdry
TsWNHi5nKWc7SYmT41g0k2P+SbNDRaEtdy9QIQUEO/VbeOYH40STbEwylT5P2em1vXwalCQhnCBe
2+rRwf1mKeAnTRZaqdJNMBIyjuotiG0Q0wThTBRSQf+VkOzla/gImnR/mk1tY+UljVeCkzIpW4CY
8Z2ZIvte1F3s5d/aPCGa410kKEJ6uHAQpnmjQTvwKNd4WnfruIB9SLygMvTGYSPL68l/F9jWEIzy
z8TVPV5fYjjdQ7VnJLIPyQXG+c0tM42kwpqDN2yVmu2+LECDbO22ardLUN/N3xut+cJN25thOgKH
+7tTV3LqQsD6+LR17sQx+YKGe3XfVw6HxkjtTR5qK18h0EgDXDCo600bSEBAyxW7gWwypbhWhNQu
sXUgblnaQZiqObykoVpg3OVw7kp5IzsgOWLhX/YURudc0hCas0bOSoT9yP5kDBwolY7dRntxHIY8
2pxXvAUlHkODnAnrUgPbZBdBr/tDXkEM1F34vELDNqModJH3YEzaZilMwzmSKZRZcOuYVOPRWK7/
EW5ibqrQf1GoJ68mmOcIOrjYqOcD4f/Y2La8jNjljqCJkO1e7LRmylxlXcrBsjAts5QEy/gxHZsD
ictuchDmhXHSmm+lz5KcIBlr2CrceAKxFI4RpJutVgztGPRAubG0xugDN5YmSLaSJLCYMLUF6DyB
xpDcQWhIGASh6Ctlk26EQd+m0xcFfxf10oayRnspfNbz6RANKW1ZNGq5+Sxo21l+xcSNP0drIvyo
Qto7C41MExRGtaxObSDzos5UB6Cngt6O0mS0BkL0w72Yy0YwhmRI+me1TAalaD+8yOUbKnnCvx7T
5u8qNk4zdMYao4NIYpaz6ohsRHJc0tiMe8zkjSxEwWQi6rewk1MggsXs8W7k7h7E4z4A77KnRyW6
3Bq0tRFzRDB0BdCFyBx8tS4aBXholE6mZAuPGh/6H6QOkpXnLPJUp6apVlo+8heq9P9xkGUELlLL
rcX1bGUaumJOZYPcoP8kerpzmnWvrlqMgZoxUNsukwRbLeYQRcUrypUXxTtHSADMwYr5fdyE1wQg
VDtFyc/6ueuvQuSNi25jL69VsOaPUuTDvG5res+/G5gsyxhsfJdJv6biTukZc2hRaTgQ2jQ41JXK
qoKWYBPuRpEbLjIvZi4HFpJtXfERhydImTMaUxTiw87MyltPohwnDLNSWcFl7EQlAAMEZlvDYVZ4
oymUrPv5NNks1EC5y06BNRa/0aYJ/AE+FA9VNEcQzsHB15nD+5CX9Tv+HauFmRNSwUCEtxcUvU6n
Ko1w6G61MOJzv38reBF6kyC4ynxtNg2kBzxWC97LoWLr/vNMTgwMxMUg8CGJJPT4oQnMpoJT1A6A
+ccQ6KgYcEdKbtvT5vgcBjbR30BGm8KuiilbfxRlUPCfZAzIsXDQpObsCxZUjadwjxCCHNb+YeB/
MRBEpaHllSOARbihbWCRVBkdHQ6e3ExWdVJUyT5kmhHAHVfdsm29D7R0g/y0zNPnMpLcghvf2jGR
Ah30OZLQ0wXfPqOo9/ud9Q7ZyMIaux2gDBpH8DMUJU87Mf8q8HHdTZIW3RskdHr2ZFR+4DNLxOCf
1sMgCFnXjaGL0u2y0O8U+T17jA98BXUubEqyZnZOOrl/oWrZ0AJ7IlnrSgbLmmtkL4tfl2kZdQhm
T7yEA3X3KBvG3BfWAdrS39pyKYSBhTsLgGby55rzxnXIhwlUp/8ozey7koAQVhXMfMQXloY+RbHP
JsWK2TSDv0XNeFgNyzvp0ysGG3S1kLgyt1Z9f+RIUqDHW/AJbPLO0o7dpxiYWUMDBCerOnxQM80T
4lRsZ2uchbfQVPjZNkoDwfVjza+8U7BNGl22tgZHAUd1mJFSOu15rGUcqXA+93DywhtHwPXoUd2b
e9q+HlTlGeIxw8yjC+mWfW64a4lp6C9IHtOYMBxbyQbEHmWNJrYdlq2P0PwNip90mRJm7l8V8f0n
XcZyx8a2rCS8qZDVNJNA6YNizkiLvtIqKIpdgHk8padEFRTScL31jWUE5N7I0Etp4bkP5n7N112E
IX1q3Kjh6RulgdH3hWt8m3aCXRI0TtUeIalCU8qPagw1jZcV9GzseWa5DhTxBN/DZgTKWnLf1tO+
f5ZodCVUQ09pu5LT3v4a6A2WXhV9ZA7pJn18PLGx6JTlszVAOQDb+aU6p03gH1MVIwM+7Eg9tLEI
VzRi9oQIGF+Wk4owUyRSi1m4imvaAyqlOuOaDhMVZR4Hl7xVhAsmnrfwjMKsWRxXhaCxXEwK2Q6/
C1sPock15Ig9R2+sTGIQ/sEuh2vvpah7PsjiGDT6pXMwbU0t59FtivbTJB3yTEveQWVftnwBP10C
dSk9iHMRgzPclcEOFcNT/vOL4jQjfdbADKmIKv1egprVJkU6j5VjMBfzCXLTJ/ozEw1gGqIMFYA5
DlG2Cv8YiaDfpV9KGOplMmImeZ3hAPav1QXMKTR0yGaALL6wFvKRwZ2kneaws6IMayiWjrXV7jxi
UW5g+UZxkH2XY+1w+g2Gnf5OLfmgmQoNbnk565w5Tfxu2I5gBBYGMEoEt70ZTtws9+MaaOP+r7Pq
Bmor4hZLyRdpmOv9ZxHRgkw/xv9OOBo1i5BAUQN2uP7TKXNuhUWwKI8OAB1kISUhr6Y2BL+7I07o
DwJLoNzG2xf9C2tkVeynuXbhgGLoeYZLdaDnqKKkU6ruhX+QJr/GR0KkWFUC9fSdB7Aq2cYX3n1I
ILfiKiu1y9hWXyOT3sdKZ6hLNbNja+wrDTXLYfzL5qixkB7SWjYwRa3EoZXPYhdb8u/SxAtDgGEN
yWon4tC8GQWxKfZ7DfqUXJ6mgz6Z7xrNZQODXxcEzKjNqE1f03/PCqYVGl9YwY2R6yz1ov9YXTUX
VmZ/7EXKW8UhWI2ei1AMCNRa+g48lU4KsF1T8XtnmnAy9hDu1eZkq/mrpy0sXNk+B+BoLwdPVWqj
qtC81pqXn4QW07rrEz5BQmyU16pZRPzlZTAvCnD7WiqimDbJgMTPAnqYNUdjFUPj8uN/XzQw44W7
Om3UyuhyGYbHmNpsFHYj17WrngT/rwg3lc9HR9vXwd9Kx2qWeL73OxzgVK0JKVZI2FLLS8Z43+qa
NQcTFXuRiT0Rlb7IrPgL+sA1jh7WnIQaVh/xlq6WQGVdIVgJ3yiYHtrZPMy4rBOPTzI3rSioUWqI
VTvDU29UBZ05NGOqgDvqpCL+4j9Jtheu3/UKJGjEBUPP8TmsE8BjseHpuJOrkv4LHaS024WQh9g2
PobulNfAhPd7lwgcRXtSPbcj1f0uYW6fq4j4A9RjYBRWycyyNoTOGjdnSbiIskPEHutGRIpMeJkc
/5N8KfmaXoAUGXJt61KE6WEmGR/a7B7KrV6iuPvjoDApq98/osC7KuAfB6HEylofxvB0xxwgtIWr
orHsg+wGx0MzqCfUzme2NOMV+Fw7iLOeWG7lAPJOtbYr+61ehsuUI1bvZQ4RhbX53MuRAU9jg1DU
3LGu35qlpijOrwjKov914XkSjzBTk1uA4+0qrirCQSd+jWAGAEF/j+Uq5PmV3KG+Ua8K8BZRKNh5
nBise1nHeOZexJSapQ9RduO+3FMG7nV+xi2RRSJUnyZ+a+7bT/qv8BPGlL+Kj8WwOWB7wVBQmC/0
rMfEpb5s06QSHTG6PtIzRzUKvJ+Ev6a218tAPGqpIIPGgffa0msJ2p0bULwVamGfwt9eSgjiJr6y
lCXxRyd0guhMbZ3GhBCMvzElIDoqBbIk3Pz/3I0A7LLMMDeeFRZEXfTBM9T5zVjunUcrrMvsYBou
tXi/CT9SSoAYPCAlar6l9Yw54O9vn1qkQQ9tfJBpieHWEXHPcEOJcrVfeZENbftuBT/3jSFPt06b
n5Giqjh/gaD1PoM7Cpe8h2AezDkpKLcRb+W5XZ5mOSDI47Bkmxk253xk4lBdvCjenJ/FFHf0C/rn
4dSbj5XZEpk+dB+r2XnGYMm6wxQpXTP/DapYbFccF6qeOqn726ZqqAwUsdKhi7fF0n7xUdS4R4Ht
Fq6FgmPgA4Gk4NllkvVT5Nf5cRx02EF9poZDThwd5v5w6MmiyKnCHH3R4lzbiDhVJL5oybuQaj3s
CTcBGGasv3N4ICMM2YHQmRsQylLz5v9sKewMx9SNAZuV8ScrTC+z7EjhtYfJKj6f6WoYdI3HKYWX
EX9l93zU1lndsZmK63rcq4h1LwBAFbW6hZCFW19cDQBkteKuQ4z1E/66UPp950GIT0etUKvNtG/P
MeiWNH/mSfSnJIndigwsjAni3eq11y47U3KcTUhoUKvnP20PR/nwRgJj80AFa8pWs/AIWY6ZlDMO
H3Nri0mNdsPH6J9kNFrUdCJMsWU4d5WU6b5c7PKAbATPaJ5L7vZ0zztKgAeNJqh5+W3Qe3GqkIeL
pmRNypEIyklaw3tk16urV4VbhhArz0eGRqYOtT9u8UWOAYE2i9DPDeUU4MsbAeZnelMYn3CnMOii
e00IyFA6eKf5ei/KD/v5J60NU0ofsfnO6+rsd3AjXmPPahzW4/CQu7blC4cSIikLDA1i/O5fbw8V
LkyqOaop2dPeg72REDyYgbT83MHFOYFxBFfA3PgDoIV6JKT50TmlQPez3+RpWjchWgqoieck8/ET
yCgRM6CZPFDAS9+nuvie7OAwcS2Jagzl7K8TzrqF25ki8Ljg5xi1l+ruCOsBj9o2wOWLIDzW7V60
H2zAKoPMcuXlroyEvZws/Afr81y1nuvEuCoIgFGWtQg57ewHldS3eqw6NQdYgCv2i+I+3/tlykdQ
cg2V4A6oxdJc0cADNtQYcpxVct3xk1BmaJLyPnMpnzwqFNi54UCbNc0FMev48ChhZpG8xe8EbW2w
tNWUYM6ZOTkp3MCeJxyyjs3VNitLuTAn7BlNizRGju/i5h5X6riXtJL7SN1v5fFzZvMAE5aJdO2F
IYSVYCVcjve5NW6mZtFKWkOkBCuZz2hl8d2lxhFu52rCTqYIBKIfbveUe8o65UkMXsLenvjT34LC
aOv1Y4rBFa86EawsaSi7F1upBcSkGrdl01uQb31VIx/DwDvf1FTAOz/XFDun2GeldTXhcm9nHm9S
qwVj+FEmGyyln5GFt1sOZjeQNjbKmIa6ov1lHgTeEiHL4yLGqf84djTjqlk4vV4jYikVz/2Ci11P
mKfArZAQO7QKLVuD2sJiqTY0o/iTs+xlBkcahI4iRy8TXKhzQWE74iv3A8Nr2bRCKsFkxMW4GRLy
OUBqdBqMilH1jm00keoLBbmzCCuJAkA5h4aL5KxAgT6LdGdj0/FB8Wo6rwz8nTr1obNuof3NG3Q1
rulLjmOpolL6lvzAs1DVBT2FPc+1LrT73v9fiNMEl5CeoelNNVh6OJ2Z9Ml1wfznmjSHwTBylHz/
QV6qQD1aGbh0uSnR4bfEnPTSHBOnQtlWJwZ4gpap7qbwzvE3t80++E90o0814aEKCwJmmyOLXDVl
09ZUTJg80l6g4hlUHQgRF4JF0f2PEaCQFdNQbCdEhsrArtD7TP7nJtOLb6TIkF78xTxCGS0Kjn11
oHyzm8+Hhu1rJe455oXLWunzOeI92hPjPN4XqMvJ1mXIQgVRbCHqGB1VlUwm01Cawv4wAYVaepxc
QSPFg9K6UtmpZa/zBbz/zXGKjSV6xnPLXAtCSVknPMfo7ad8y2v3IAusUytM48qGUAGuf9NM48CC
v4VI4H+7URAmU5oiiVmJdQ3OBaVv/UMAiPQE5S8LkIKRsVjox60cLPD7eSsYQX8fcKnpPlV8DtgH
rzGRVCUP8rX7MvQhN9kXdBaI0ocCiFmZuhLpOIfYJfy0rEbk+BpyAoqu1DMUwlvsqV3eoaeW/vLF
Z2SgTDap5tPauhTlfto/9PkWX41ZmJ2e3/5MFYK0wsdIuEL41sVUEF0PawXUxIDpkDXSC0HtRPiz
Siplbnxp0F+l5+RtqXFO7K6tyfpgQnOJIDLk0E4Fzgv62LKjmxqSg/mwgX99cSANgLLKVPA7dne0
kcs9ydYspzrTIGJJVJhAUSrNed3IWe4Fnvq6oFSJxADBQ4XxcokowgfNeg+3sIOPa1+Z5jTbW2xy
wH1DNseY8FS1+PXVH50MJzdpCSIB5o2LKQ0EhT9OOMLP2BUbBjoGIGGq8SKi0+71FmiTRThZPUVR
aRtc4g5L3t51CjcoC6sUG1aG8711g2a2kNs68mI94iyELo9ALePJLVeqydX3zZBCtM+rn2trj+Y7
HCjCWzMHwi//5liD4eASywWR6sK0lYlDymKfR5HIqOUquo43wzuAS5F8QxRNJysI64N4dzG96q1d
N9wsOW7l7z6bSWLtnGVz2Qv0GzSwLaeysx5kiu/sdkiGJfST7kV6G5V1btbzFMoPZq/rmFZTo3hg
YZoYJQwMC5eIqK/naiWfBdla97vFq3Di67J2C/f14fdNgdhvkirWBFI5fXgdP5C6EV/kKrM0g50W
Uy5jSX6sxst7kUnUV7/J7rfjCVi3fcPJVUPSAik1AoFl2mZywoK3OBMG5KmLrycbvm31tUpXlmHR
LVvoxuhITB5jXGRYILR6srArYfl4BbY1FsDZpdEK1/zpMvCt0Zt4zqX08MNKZ0Sj2dKdS618fxCN
/xcDEnZ82X3R3kqRRB2EmhqKlWB9q4Pf5KV2JnDANbsHUIFwQjSPz6bsAhLkvXk8t+TUfsRD0i99
DIUrnV8hjwU0LmQJlI+9x3iQtisziL/U3xxAMNrlAUhQZH7kzGKbFa2e8GonNGCgz4bCNSwZshnY
INtmvIUDmtoldg1x6jA/WBJ4Q0KdOj6Yxcy9eSnf46ailSxd5YmYly3IYjg22Mxc9lNULapWgxxz
rvifFgM1O+3POV1cvYWvnEhzK0IhU2XPr6K2c1KGswSkHNsQ5SHdhINNzTrNs2TM+DImhPn72d4a
E4H3FzmmbHQA541T9pVkKcyb7GS9dMLfGy0ZhVMbMKHlV28rBt034ILcwnplzIJaDWdCPSWNThA3
4bvr89BR7Wiy9KnyB6erlYfwKVYXQOIcEAZ4uB/Zu1/ve1sfiVax93Id06pz+rUN8Z3fvpLrgOn4
hE8rWpijARZ/aboGX9JbK73uTPmYUuxO/gL//ByomAlOvlkWr/ZDqcgy64tGLAY0qu4IfMYX8ip6
1JcN5kPHF4WkZ68+qoVUg9rmMnaRNjHtJA0lMYyztgbM75M0g3Znba7QhE/GXbJ+/GrrQ4yA+Y/J
V7Ys5SnPC3TLfTz3XXzrtFunmjnZbxpEg40/otH8wWsQ7ImU3sm21YgjDlyxd5uWdHP4K19OOoVu
nMIr5Coqt4eS+dPzZT+zW9FCqkBRBzCGmEgSXZ7m73YPB8G6dUUd0nJ5zlFny9RHhXaxJ/mnUIvu
J2zX+nH5GYfjqnN6qmSQDui0FZXX7OmTQv4w01ipe9BPvOK179qwL9QYTPpyWXkFrrFw6y1MIwlJ
Hxts5cpgMrbLt2rUOT3GQe2YACD5iK8raEnqErHhkhCZhaWodgr22MU3di96qBuiu6oJMNgKSNrz
tCwawspL5unyBWJHD35M9mXFcWUzaukCX1MQ5UyKjmi5lTzB+CSYkSDXA35EUD6cOzSu+1p4GTaN
Jarnr/xZiWXEo7DF4nL20rL0CrNG8107aoEfp3C2ickzbP6+ZqdwfKU2P1goGQTZrbU2XyYv0BeH
5OoTE5yLSBLPe/9q2NaEwwM47yD5+oEIGXy25vuqaWZRhtUmAo0hzniz1Lc8u09SxU/5bdueMT00
wnvqYWHMlpRt4wdmMOAx3v7P/RpSlgTCq/mf8xzl1+FIk7Fa0kSJwD1lWiIyBrM5GVvE8fQVY3dX
dCtxpZrrBPMVIA+ghjgOyzgjbHqd5Jz8rNiTvoekbFWnsxVmJ9RTeXyLoaHso49dYBIb8PuHuPRP
OcgVZbkX1MK4UchRAN8xq45rsidprnOuvHCJI+b4aKdFBh7rTqTZc0833fMS8j5wAYmbKU/uhNU0
bostqIodSIrKFl2zpqFpmsFQyvwH5ADyVW8Gqhq4TI4r8UCK7Y9S19Yi8A4OtpMru6vFKWhfoRcn
QdFAIDWROZtMu/kdmYTKgmsyMOM21GAvRzQ0Y4zMnaQNNWyWrS6XWhSLX18mVknVl4Bw2vqslqQf
FxiM7Tc2wi95wgfAUePiVOgbFwr49gXWO6SIAY3GDyjN530666bZRhJ/m+/TwKIrU0+9YGdweEMF
qiN0bJ+YDDOMls6R4NP6CFKnR6Q7pO392nXlS4w/ofbKjqHclifLAAPUtGGdsxgr7VyRP2uZPdOs
xpuPfB7DPdl/csI4YLpcxl8U94tHQ/FG95W/Uv5Z+PfL4CWlAo4CgE8WAJWN0Fy9Q0+qQnvq54A7
zhGOp9h3RSvW4vCYvCzuhkODACDxJUCmMs2RMHeQyM+V1orG73B739OqY0BStH22oAXt/s8ddH8N
DLjyphFp+Xn5eXvC+u8bGQJm8lrHJkBate2iSsLZD77HOUcRxIToxtvUwCPbufvr71OwJQAl2Clg
XiXiw5SUrs51dGChuPMuzQbPVt+nQLMLCS3moctoVrbtZ7MTclPBZmQadjF8LqLRMYhsEOLFpuV2
evQcFKzhGQmXkzRA1JmHjAsyT6mxQ89DpgaVcbCJS2+o/cW2F7uWHmoNEs+y+NCxXTS2qaZ0ikY/
NLH1gAHEFo353sDRC3autrQ36lw8aXh+QJbc+5QaSTzTEFOKVdWg13e08xd51/RSa59q5jgBtJ2/
ZJBpno7QuUsGgHfxbq4bE1kuBPO17fFYxtwvqJY2NWTKpOMuGYc7cxc2Hh4SulOSciMRF2tl2GVN
DokUyCS611cw2oMIU+skx8sDmYIy0QOQCLjaXXRFEhH/Ce9iZVVzdNEo57WYDBarqShlWGfJvRsV
qA+A56hq0iu9hw+iSBw/XlAfmajSfueNn2Da1LGfe8IhnXjzvKKhNLUTUetDP118txyUM37IlrVr
Qr1CA8xg2uIP2ukmbHBF+c0xZQKtp6wmsU61CXDhqY1j+xD6tc9n2aeBBV//fY6M5UIJkauICZ84
USJKBReSOR5vWBnGaM0y/Lz6t+GbDfvcBFwgEG47cwXSbboWK9LocxLnlFssYnBPk9LvLWMM9+1n
n/GkfmZs0Dt/fyGqMfYnm2WCiqJxaT/sfv0A2yTPrOVVxJO34DnvmDawAqzDzJBrmepChnLRAmtp
xBGVQpII3fzQpikzc1v2hQ/7F8qvzuhjbzeblw0ETXx18qKTC3gltg0rBgk2iw9cx9j00toMWIp6
yaX5XvNdrKIlISpi9f6bqe6b1yvrG3y44uV54Y83AyImJfhJZc75CUZyoyKIjOo5YW1fqV7w5Kay
t0OQK/BrhWMn4fPbIhoGkMvodMOp0PYJYvv9j/lgUcKg8Qm+iZCZOOkkPDahvSvMh81me1k/IGjM
QfXxuVBodchAfmbl0yISmAbFhigHu0givcJllMgUHeKluh1kFe474IJGrYMlYpfu8vRHcah9h8k1
n292c2AUTavQSJ+vYnf/5cucFXNGB6ZY3KGKrlPx7lIGgQ4yyALWjJxyXfDYgAT677oCRYqS9oin
5ViSUr/uLltrMHscwuBYLswpKdFXdwLm8h6fmCl+BNYFNIAkItmIpf8NLVQczIbTgI139FWuiqCD
qVLOHrxIe5SQ/uA+cqG4VDVu36mkWxs84D0XZZdQdzUO+yEUCxoq6qDFIHUBddG+8cqPcSnzjaCa
j+CX769CCNNHmSYdEhrUkwwC9WnAqXnL0kGm9kwUoluBRO/6gl8dG4VMZAN5Igy4Ki/oRbKQi1IX
IZVUEBOh5OqxJBdTIHi9BLUQfbZ7vFR9QBrZThOCDT3CdsGDLHiyWh9i5Y+8SNzISDufibvImcMr
WgiKT7ym3oTHTvsPxG/OPz1NbIE1XFBasfJ1Ys+ffrukBchuCy1uhK9I+66LUzEV7zYSkayhro7r
DxwBGSZc3y8TMt3gdp/bN9wbl4IKKKvSMkFfa8pPKxrpWvMm13dawgmxY8Z8t6FZAIdr/h3NB32q
DII/jjKvn1Fw9OhcajTiAvCc4wtmCdMLQVM9CJ2TJ1EckMkTwMZdA/n3lWnRmAVIQpZ37PxyVUCG
QUKoXBiI9GupmpYY+lCR8ZIVbMnywVFRA+jFMK5mSHoRhaigwfbqOrIKRZEWq+MKxLWUMn6jJBue
vVOcJfnVV7gpzoIJxELsRM48e01gn/VuvtINB2wn40BGOiOuZAeB/Q4kYl4PuCT2nGdEtSOuwJth
ALczPnI0UDpzjwLdPAWHjs3PRVeqabZHUMh+IDe+vqJBy8awWd+a9gFVlt4g7GZbFKKrRDeIMOkn
3HTZUkqcJtgMqKS8VAeWtcCEWVxZAwAAyjyhhju0L3BlvIcipOqtMeRikLiJBO+WUDShbiXkBYiu
L01DSwsEHLnMQ/1zTc+AoLaIy7umN9EpbraEbOaghG8seoZgFM2VjpbwVrI4dtq/jiOBqSNoL9lu
DrWyCupXdZuVcj59gFr3sojqRsFc1Wtq1+2YFWQh9PZ7FotefUIIvHhbA+EEbtPE+/01qx683KBp
Ofjvym3lVJEBRZfBHWh02WwUxG78/8eEbCt3cRTNmBeTGYl6J9rSi5fvk+A2/HAQnd90DougrlyM
OKI5doSm8inqtvfCk+hW4bASD2zhYxBWITTMCnTCdzjtfgx6NXQibfwK6opMlvXkp0TkgzuUZhea
jHH4HuMJMGRYZcjiMpUCFN4IF7EwhOtNR1lRGRz6JLPBCiU4Korq1ggnYlBecASUhw4vnQe0eOms
Qs7K0aMTedTJe4njuT+xGJLBnmWHpiDDQrc566a+3NFYAtBDkUCgvrxCg/0QX4ISEoSg6G/Sv/iQ
imojFWuMoOAyyXTNPJPjY6atbZGRp8U0olXvZ90s6zJeo6nZtg4DelBpIAumey6hv9bl9rytCr2g
fPjM4UKK2/WdJnnPV3ovGbaf2qmsdtY60wQSNucmVwlRxusxiMR0tHkHEkXeAol31Ac6xkHdpinP
jTFRkObTO7DUHbnRZTPC5K0gyIioIQ9jVszcIdkOV+7EotYrj5DRzZ2vZsOlKMq7KG0fbZl9FnP3
VQW0oTtL1BPn5yUfMAmc5Y9xZWhCl5u0gZ38veqwEPgdtImpdrxSR0omp7Jta6YqvxSPDwTKYGS2
qwTcJNtATT9OwXd56IPdlNBSok+3yYjX7gowejiF8UVlD8bXJ7DvnF8xay/jBaaT8RLVrpNIXwMk
HwvViu1MCs0OKkT/VKMrberPzBZdTJEwCUonvEyeX8xyCbGespx1fEWMb0Tea0rlX/db1wYutQhE
ADWsQyaecVQIdi9ESS5QJwzc7SJA75D6L37X0o9CD7L3xqDEUb7TeX5W63qCiD9I2tCiyaRBRYys
ruFrIVNy4G7jII7MJtV14p6GvrLqAqjDNna6vaRvXOX5fSXevNv1ZbKG19f+CZBU074YEQxvxnoP
rtU8YMOUfBP/BKYTRuIsDF6bn2lsRpw45tHrtkIkQISNtHqoAnOu6yd7eRVH0r6YOa5xEeFx52LS
srTrSzyipITMcIiyi7B3s3YE3luRAHBq00i1PsAwIqHoxRuFt5JblcXRqzI6Hws6wIaYos7kudym
irpja82KTCGGISkwsJZUN+Z+Wqg6h2FoBHnb5K/kp+mC1725NWKXFfriUijITsviPjAaXdRgIOpH
pCwsWXF2TIfYMREbMFVgA+ORG5UGbtWFnlWJdqrWnrftjCaZ0VWstCuYSj3AE9k2UB3FN/KFN/ND
Sqs7n0bPuk+EG8rvw3EIBC0OebTMMHWe8/5lIqjmdum7gdfLFeGWws4uTbr7oMYufEnj3lZ7i+Gn
qPKNjYhgnKhM8WgzoOCVCQCqsuqC4mENEo3gr34AVQn2Sr2z0340XbhDwqHOPFY2xBGB6rvRDr6c
n4XYF7PQKXO7gdiFMj+zmynjWQphCMYiRA0wuS/azOBUSiM0lixUamevA3iBTRVEhn6v3oPlG+jW
qdtxg66egN4XmEZQvHtfyV01lYTpuYl5VA1tuooG3eqoBBUxq6fUw5UlcJDEUjM/DquH1oxRAGZZ
PUsyuRixAXsy9JAbgHPWW0LYr3mwV/aJSM2D714+DzAybB5T9JTcJ9GQ81AWZzbu5QGNBSIivifC
wspy2BwBKcgarVCteSssTcQyRwcm+Jr9kJEE44gzn78h9fJnM1B0mvZrne+xT3jZRpYLO8uVKYf7
Ipa8lt//Dv6NHZAQs3oEHDtXcw6zfEMSKChhxg7lh31zAidxL2GI5tzaUvaCe0OSZatD+5c7/8Y7
zFu2Il9bhAgGd4OyiGA6Dou8uiu6jYjqVFTqJhRBhaYuPL8g3fk1LaT/J5q5lPPM25ep89ev1NJg
OZZyiaP6vBt1qPCUIiswzlnetqt/EFvMdd8K8kse852qYYY6wIhONBjmwSwmeGOI6jkKnM/w9Kkt
LvH2SBBCxNtj/kHaZDrq7PhU5tLRiTwPA2xAV+ooDBPAVr6L5D0w3t9PwO/Y3jFtUfa1IdpT0UP2
bZjSoRqr66FFQ5RtuxCZhZ5KAYhc5Mqa3+L+0fVidj09f9keIENoMoBvUUMuSJQZtSRjKoys8kVx
eMlwt0hJ6GY0QD8MuHRA8tEKfmIOJXj+yqt5uE49JsSgwaRd8PMg8IQTqTLfhIpMqKopAhFIkb+p
HWQtxyT0w97nTIv9ZO9sO/73Ebvy7dUmsu+RqtulT25sz+pwoUY96dVCfNWe55KCVB4MXEnP2Bro
XpdFedHeLzP3kBacfSmva26Njs7yyEu5eP9f9iAngDx/dD11ih0bZiX6YUg2cD7ELrfi5OCGNk2p
MTcl1702YPTMRyAFT8rqA4XSTJrlv8+Hq3S8L82LA0njseJyg2iMC+4VuccdS4Wyv0SAVCvtVeEk
JU6ZO8a0H9J9Rv1ZcgSgMdBXydOVBaNpEZ5Ysh6+WYcNH6bUxFKfuonIxd1zYjIKB3yCkuwt+ycH
37VnNGbnAANJr/cwBaQbzjTTwGSPu1ktnaBq7tGbN40F1gT0ZEEEbiyRGvqeLbzT7qukdO0OC7W/
JKa/VftRzp8NGJTQpSmlbi8yA3MwLZOIK/TIbMwzEsZunnqIjZq1buLoUwI3BtJqi8VL/EfO0qrq
q7MTHPDZ6Wtk5H80iixemsQoqqMFGDBJzdQepkqKtEWdMU/CYtlFqBwxwxBWbTQP2pNY6QZmvPGx
kU7mZzTNUYmpfKX91NFOza0y9WI8IE6HeKmE179v69zl2KT7dmU0axNcl1U7YSNE91B5krCNutvD
BAPjCdxoWYq2Q2FiTDXuBrAEZCFhGg8wkQ+VT6YQIobKUcr6eHf0RInLpZMKbS0lGP5YOfgEaSK2
g2cMLS0A30zZ2VI/pH1H5zMmh4WyITKuSTj5mqYEw/bWdmJCxQ4uQ1tdLBP49LJjtBJm9AWbdGsC
28yrzMs7aiu/xuh2UCy5Q+6oWBCfbRZGowijtia6GUf7TdH5NOdUH3A2UY2qIJuPz32+rh/jS0zQ
QmlOKKvHJkYlgAM88TTSUmdFu4Q8tkE50moypUmwB3BIhDDYfpzggOFaWoRKbgtIEaaD6QnlcWy1
A6c4ZZ4QyKM01V89LZe1vDkZJLzz3gcb/6VCWZaMe1y5vqQQDDcWk6bQPJQYJEoVbGKZB32kDzgG
XDe6HeCJ8fWYnwCkqFh+7/MaFfvgrsrVMg9u8Kq5cHhbr/S+KcOtCGqojqv5tGcwZpQVWUaxqLEg
0aV0Vm4Wa6MfuABosIvmHMVw4yO8dm8nzIee+7lgZQk824UvL54iYS1wJl6V9Zzb+7BW+8WeIP1+
U6YLj7AlIuH+IHqX4fAGpmZfJQTOWvM5UmZ5wLuqL+2CsuxzZ0rVJ3HXcbU5kBqD7i9E1ucoXqkI
YF3G/VZX8PCr9nXzYd2i3yog4CYzXNLqN0q2pGjo0/P1kaLX0PD32XMJj4wOTlgTtfP+GSWmSQb0
C3bATX51UBYL9TiF/khMg8k0SHygpVo2q8Zw7TxLrbAMCv5JbGS+WYrm2u+KGBblq150KVUAtMzd
oNmAdZUvX3T4bYt45bx6Ufzy8vJrv9uyTtk2k5zV4415L8oqo2TDQ/hdrUO13en+JIoiAgSCqaVQ
+mlrKyY7qY2Y0bRanalky/1ezLa5glyJj2XibQ1km0S8qE/fs/eBJoqGN49zU6FG9P0q3yxVXU9d
kaW1SdHOhrlvKqmnj1MChhhpRri1qhptCzJtwb6MKUwtYfs+kygpeDRvN5d/ympSLY8YnXlixNvK
c7xOArVgvD+xuMHdH4gegfupMEOmQmhr7JPKFXutXExZ9/R80Qy6E7u8oD6UfVjYSRFcsZahw/Zt
aBH71JD6a7JhXhn5ftXLB6b9CC3CKgH2sux206lxogNTg80uowpH0gaGWO6NaTGeHqHRU1xst/qU
WtLGs7mI6+j/X1EK7pytBEzHrYBuTO0PvjVzzt/DMNq/aI5zWjjeUvY5b/NYc7ePrSFDis80ek7W
+u/30cYsbG4QO5NYryvkj0FApFAwJZkfvWLJ4nT4AbRSWqwGK6HYAEJMdztHPDhTdf0aXRc63pvy
Q0MjwhBAQd3qd6dfrRA87ZQWjZYPzk5quoMZ4jy/ChGFmE59Bu0eTy+EUJx8BJXvZFeqnDu5DGR9
4j0E0fdLnXfBss1EOer/8o439mWxSwFEvP86azJHzLZQcM7cHqCjg0Pi4WOPXEiQHljjfScO95zC
LBoQezmE2GCUCf+02X+1kX4DqfnHJkCL4ukohs5qrmoO9sQjXq5hk5X62WKKu5AZ0dJqK1/2hV4i
dM+3yVLOqDT3EzgmygfixLNcqgoOoD96Tg6AMvNQv5QzJwfMYxGVLXE9U0T7V2swkGM2a60EmERx
5s1ZWGEx17kzolQMzuiHUwSZNIoTjz9VbsAkCO901FnV+PTz4+RbhcKj6pL9Tf3Mt3usiApIXdbc
mmE6wW/he6uHyPdHrguVFdiVoIdUYNbkvzBpyoJDy9j4DM17GRJQsYyF/ILUCT2kEVHokVxR405F
76ZuKxoXxxtnyL37BL9ogizhPFKCGIVPhuGll+VQ6T+izbUVdc1/dAbx6HinZojAhpfwA5mTQ1e5
5TY1f7ICsY0Kfj62HguQl6/NICEHs7QngvH4n33XP74Id8XdjXBduSuevTpo9ilwfzYY72Ccsk2v
NiWqCkL0440qYoTdONlAxXbLU3Dilpzv3rVC14YH+5UxbZ/D/NA0BBah+hygx9ofAnL9NOmdGrs4
1a7LzCnJ3/+giKI+iU8vmofj1BhCx6E/fsDvqPY1einE+mg+R6hL1Y53lmQo2SR1bwipdNGEtwh3
7YnO115U4lGhuHwj/RnWwoVXfnyvDcZvTPK8tKDhUPDc/2ZNkR2wUaiM6gLejgBnOizS5DiiLY6o
QzFIBC2jY8/dKrnzxmsH8Tdwdz6ewhGflvnGth2r6IS+6HA7yy/ZyF5qAh+GPM0o9+1XZT34flxa
T7YOjIyo9G5szDmGzDn1DWsM9O3vuyyG4kmJWMjyHn4jwQ2wxCOMqXCRXr9oeRDlJ2Egn2L8mcXp
JrHhBkc9jN4zQIfyG6LoClbCM8UmRL0PKZ+J0qu0kvrFZ1Hw1fu2gZNXC3uKhtz/PD19JY6fiOhq
NtxCMIC2a19n1Xm0PHEz1JpTc/j3xCO2lmag4CleQs8iiZ98ITFh1kK1ccnr/acM0S1OxHMa4Fog
kTuZF9tlBzK1jVrC5yh3/mLfRmdJ1aBfXF54tLQU4AhY2n0OiqdBHPdB2fVk6X/ISiAWUZQniQ47
vr0/HivOvauvfeo7jIiaHpyKU4gvZQf1epm2MCNGgTVcc6zYFndK6mYUqoqFOi3wgZk7IGAb/7Dl
TKn06/S4lPLJs+b+1KeaqNcAkEZXshDXxA/pyHnBtQ7b8nJlCDXwH5G4Fq4+uTefl2EVrnhpX1cQ
CnsgA2NmWp877drLs70mlBuJgahwJF76QD9h0CH7ncTCtLoQKP6cVQ0cNMVxvccc1+obR7OO86NE
0u/J6F6B829Lqj/pfLUSZSnTDa/gjYt40z+JDchaXCwNqdj6i5AsBVGo5kegjLzYWV/+3k35rNZ4
dgXbeWLqLklycTQ3/cSNQuWTKGpSQWg16kunGux7FebRFds3pYQMvcNVcukJMH9bUJZQRmiywfzC
up4mGsrSprxKFgRUzK7zzCYhKW4hgFyZOgUeOmgbDjEbOVJ0BGlAgrMijfDtpV1hoZB4HAnqM5R5
OJRIynE17kEABqzutqG0QrXAxsBvVTeXVRmBm0Wj/xzcscwfDSM7snOR/Dxi0L+ULUcFvDHUIpwh
Y7mailGN10L7esrO0MR5DzJSKqKAasVeFkVp/Rvrc3ueDkXoq+MUMIsm0ub1DMrTe6EPQcQOxT6L
NdxYJE/0ncaw6TIzUr162qsHiheKLA0SHsFL+CfmabpOtbDQP5wZKGVRG1KlBYATqVurhqxXENJx
wvW9NsR/gSGfBABOg1o7HwypHUVZwJU8vR1qI1vG0aHMnxUoffhLF7UnkQuA8rmmRCipaW1MysNN
fILa1KN6f6OiFuyNx7Hpoz9nqWG0GVx4CWzhcqwAI47lQeDZ0muf66mQcYUTl0elZjTVNHQdg27Y
d9U0/1qVHAliXAltdy1jboG2bw5Gb3BM4RmcMuNCgA07K7+oHMDB/wq3SSzFxgy2I2Rbevy8IH16
BWEFrU1LY7vlEZAJqKECmbf2+JFh6N/V2hoREdTYmB0mTqKfxggBEd7mecrG4TM2+ZEJNhUX+Siq
z0s90qOZW/Xefd8WlRUxL+PfP2pFc1snP79Bu104B9d49ADzWMGeP1Km9P11mDn2K73Lz9JjzaD3
NcyP8ZcHAuTvslZPvHHQ8pZufLcH7FFZqBnVSkt+7zRxnRuVXIRrdyvtNldnKRpRI60IOWfPR9nA
9DMn39blyHlq7bMCrI3d24Cz0dDcfZ/sdwB1aCkdWYXhfU/NFiMMcYURa9CTkCD7g+2dh0gF6TGZ
8WMCIiwTfpt8gW+TFULiU5+V7qJTvaF9gv9O6wGtz2O92INDMzPR5RT05X0HsWMf1j4Ms0PaFMhe
6WMTxqK2XwfU/0iBdcVQCl3QdcHfhSgIDcQ6MCtU8iJx9/3KzOrQwK1a3wac+lmqX2SVglyvxbxH
tojgvf6AfSeaLinNrmL9AqVFTFlV6BHMZzhOGKqfKTWbABaDuG/zpBoorxoyFV82lZd/PhA73m6R
TR5+JvjwDv359y05f+ADILoCPobbAHD2sbuobKQQgETAm66UIXMVEeFQox5I0T7nGHN1jKvO6zN1
bcKIPJugHnvRgk/b6znJxF+PvRMmp1XsBQUbcS7GYl6q/o/4mxlr2s7ApSI6BUotxtnLILxbhNk4
tlXH1Br4X/5J4eEdWkZIzTGO3NEbyTffgQVcNazlupe0Sy1/4K2dVpxb7Z3HzdUCoQUB/TtYzSN4
DKzDAGx2azhJHCC4Djml8d5M4zkyNeq3R+s1OSaw4nBu+DhD91Z0NiDFX/ucCvEdOW64kkr1t1GM
V+Lv4KceSPBjAIn+IYCC/OlnaUUc5XXDIrYmRgRhECD20yalCeIilVshzfw+RdKklmC/tpko18Yg
G38RyToHFb0qVcg2Oh9gaVoSwYZyloNxy9UBPjSH6fc9rBIDMcc0B3EAuFjbyobt2tvNklWC/zWb
RVvgAyf1vkvivSFID2O0grNwXvCpedfbJfiAZyo1HQpNhJuHpo8b8Tm++xmXCPvDQjO+Nov66/Bk
2rQ3A+hj/JCKcEo/Qx4smzIevGUMyzVD+smYGmGJluV7vr0TTiXR1siHlYONhAdJTFD9msgLSSqG
KF7EGTNG2DtiDH3SodU9HZjwgca+rRnTDfRVYnbioQVUFz2I0NoBoRtj8dhW2AGtVCZIQL8Ph1fd
RfAcE2Sk0350EP/Xc0INQfDoB2wnFk8tbnT+FdjSwARql05IE+0uFHxn5cKhh1GWJIbYSGn6Xj8G
YcVms7izM7eX6+dV6FgN5bZrEAvNo0LAZsCiU+6kBCWn/XcjoONwVOhfjvmpdnhDIUPPd1606t3W
AtAR+gRDBi1ocrsMgA63aCX9Y9XezP0oeiDDIzKNWkbVg23t48ZIOnJ9d3RfSZnE2MBbhCwZgn8l
vNEf0aqdN6/omULDIjcrjt+Jz5Kx1JQiepMyStu19MpW9J6Fg8JgpjRxOA1JUhW2aB4YreUnRqvX
388Fifmi/Bhkg5xt/V+VmwvO9AHZ/cZyE+4X6xZMjL909yq2w2+OoKQukETOXKXFL8tC4AAkZRXZ
ZGWQs6whElxXaDBGslAnwsAuPPbTduM6EnVZ8DH5/fgHglTRPY5lDbUJ4wqQfhmzt5xVbpK1vhqu
6h/pV/oEbrSKYRM8WsPAFV4v2Hg3E/IO6RKym5d81eu1BiiXn+uQuLjRNRmUXFaPpfYtRkbmqx+F
CfFkpTbleej7PqJQYMcpffSYxl5sTIK0XTrTM9zrBMDxLE6X/sGs6aoajKCCSf0YvlvsIiZ6/NQc
Ol4b1JYHz+v6lvgVB0wtQyICszUxO8xK5Vvy0Rmg8TRhpzOfuGvPsem7tGWWsj1lQ67ns4SkGe2/
zl3X9nEfRTfkkxcHfQJWbEf8Yaxnk5mWrMFXjBHs1DU2XOTbGEqTGKE/gZung87iy4FMOnHC0bN7
EjZ2jxjO1Jr6MjNAQYT67r0+E09p+lNmo0NuniTt5h15DOG6ulSTfncTZ5sjHym/xopPkKNOk8H9
u+IVymmk6K8fcqf5NnpIIMHhwfwdluj/CO8fROsRhzeNyTYvGljkfyQYw48Yiq9yJJdzvZ6i/A4r
mg4zMddxzujcH+EwBkCnIBmB0OJCsjZw4MGEeKriMPSWZnOhGggqn3MblFJLo20qVvSCKIZtM+KI
JISylIAKfMjCBW/ZwspjIsvrufsJe4jtY0AsR4Rl6EeTvFLFHs20i0Fkx0RUMClH28Z48Ko0do6/
nGpcvekaMYhp0msADMOJKXFQ7oVjqetBqbMRxc5R5FrxYyuNfNug9d7fq9N0grV3OsoqzXVqg+NG
1NLB9JsIWYSBZtso0vB5zhPl98WatZNBiybaPoeV3BBNaFQUAe/zdozYZxGoEo77sKgjr2BhGfEG
1a3lb993BBhKBssSwc5q3YnHJ41inAq+3Arq5VfLKYRLEWCTCWHvuPzlQRsapZKvzvKrkkJCjhSk
N6z1z7yo1ybtad3actLyjUoe9r+9m1q1wyFFo9CQU8UzluyglHbQ6OpeGDNusmovCURYb4Zz4zTM
6KU74DYYA2h9rYiJH1R/6A2RlRIsLE1quIN+R5ruRdKfvSwagwTMGl+fHUUGfeDb9zuROckMdGlC
OY4xMfqMYFKuXo11deWyhWjsKohOCyiU1qLb7zXg97Yby3zuQhUuNjF6rxbvjli+zi1svl/eKVW3
sYGxul/7FaJqaZXixFRzudS7Yudur+CEqKxZI6SKA7dYNpMxHmRG6M//13q4ek6GKVXT+2faz3nx
r11XJVkgjPrsY9IugqnTLNfFlFGOe8QkhRkXP+mSKcaiBwR257/pumU2WlTe1sdtA9QXe+mfZOSz
C+PgfDPCQEq4CQgWfv9l55aYIS0EE3Z00N+8d36pwHHek/mvphAhgfxn392zzzfHhodnMW3WrfyQ
xDX3/2EGqsjVF0GUY8AUtHjaD8wFCt8qoBiy/SnYZ8ZHY60xc4z8/TL5/eU8IRRDobXOn8HxjAfa
zrOUzz5TNdkjzu79ryFgG5p7bwlFwnI+NVjdzZCdyKYqY9MecfUvwgJ0jL8PDHXD3QjsCqyx3rx2
jq7CAx+h2HPYBqv9eq3iNtblbNOZl00Dszaqika3fFs9Q0llIVnFZ9E6gqhW5IHmZCBNJag+ReMO
iBFQIz1d7ZmUOavcE2qreE+tERc61u56Zb8nlCSK7cQ8dvian5bHq+BmAG20zHN7hrPoOwxSbNK1
Jg635pGTlb7D1i7NhKSWXKrR+i8vwR2Ktggi84cSja2dzn99dBMTTo8LZiT6jSNiXtme8hu/KTvY
ZwAErwlD7yVfpQdgngDxfMcwwlLaO2m9vAJV0wc9czy7BCSQI0l5hLkOOSW1/FALJGuJvxjNpxkH
AOQNA/JySq4/CiNOyz1gkEMBt79eSS0ItEunao3LHQzOxJnSTjuntFg7RUYuExIIGNLw44nIokDy
iL/0GEUWPOU8QAVZlNa1R64icACH4D24bYYNRTpAoNXUOf/z0CtG3p0T4ZPBAb7cU2R6AbXCg3fo
ZLUvsiDaA6P9kJr2zkGEthLoYF0g2vJ3i5HudDepZ8M0RNaR9LIFgmdIjW6xU8YNQJf/FQC58R+R
MW1C5SaVF5BpFYIiRZ63aXzQ0s3kPHCBtEmOGilPTaYXj8DuK3HS6lOdYMe+jkgXihcwujrh4HRH
jvsGIs/SKiID+yOmd3dZsYpCgPMLbGWtFYXooMOXzOcWqEcytKsl63Mjx8JRG2j/Y8P2jLrwb4cG
bMciGmzj6DaBw/d7GXj0QFgnbgpbNoiQ5yphqyrvkE1WbZYmQ0NA1t0gMr2DaFgYVIFT93ETay7l
h3iy8hHBK/vuQERQ/XGEYcrvy0QLDyR8EWipwpL1fVKJmP8l5U+RehsRc4sPQmqkn488Cs+P3fHs
8/yuD71WyIic08443ggwjOCnYG+7IqN0yBc2X7l2YpffJcaYnIPTdurnDZPvQm4Ph9u7q/LxLX7b
F4Yf41v4090xKQA90BmYJZ0ugtKqO5fUb5+Ayhd2VxSfIgLnW1boDdrxr6sg0Q57RoH+iSlyDHNC
nZw2KCG6qK/SXlZzlvSbsCg20FrGoDbmWR4SOCOpn9ZqEypjW1LCLPL4dEMo+EVtcIOJZvy4PSwy
St5Cvu8glHcdPH9gAKWiO3xildnlTBSuxnrZOd9ga5LxfvxfwDRcNJtENzamedoCLVN7OGkqzQe/
7RPRNenTLxqke2cAWHNhJ1eQSaNQPBrR/OzH71+AjR47gDeJCD5FbeRPdr58OTFN5yafuFGEFdKd
MqggGMD72/puXEuOJCf5TZPOuGK/zFWql2H4kGxUga09116gDPUch5c/zXIQX/sE/L91rioWCU6e
z++72kHhEW4ZXPYs6qTcQMl6roe9eOTlMoB71xsKoOyRE/G3TM+wlkXeLlhPSe1xx0zTB5ZkTc2s
IWeZsLyg3se7juANO/Vj0KE0iO05hvvZfXXNlJ5cqshDytJYjB8ac9ZbDTy3ydqN28CWmhAxc0p4
DJXWbO16d5A3r2tLdGvjAjF7/K5RgEry5DRFwgX4y3eJ0N4Mm3sPzMozf0J00nh1Rk6naXk49nEQ
8nS98OEKoHmF5AftUbavOgCx1SfkiMLynGAkz7SS8VuLvYiAVn0xP83MRyRBW46EUwIPsebDRqMZ
auo5LXUijNmWI/MkGLhj2PTfngj5WZlcwHqHh/ywNz9yR+zSqN0cR8t2U27l1ZuvxORECCbrOubR
14hkzVWwawR8uMA9Ny6yIGA36bXzZUF0G9QWnSDFkv8Ij1tLbDzsHfOYhKOWphtg30MmaLetNUvw
+/H7G2/zkxKEGpXxIkQ0Un1B6rGuKdvwqknnplScXVdokg+4oxzYLigqlfZUaERmr2RWZNAnyWfl
UtMIWsPMlWZuxjXtz7NnFsGA/bJYTqrehI57KJJkGa0HnRQ7T0kf+qxBd7X2ryKa5GwLiNgqRieW
CZD8ckt3UUqueeB/k608s+slAGwTBs8in66QBM1o3drd1Pdabpb3G1YTobH/0b7Xtxkbn2icrhIi
9cbOSuuKfFDwKO2p3rIWQA3MTkbq80A9LBDpaUOfQLmlQAe7GnZYrKxGMEPGapb1NGqif+F6L3Nr
8VVom0MoouNJZZJGAwRKa82r1k/5tyA7tbFu+eKyZObFkBqJ+HOKLTPAcDidF+/53BGs4Sm/OZWB
x8rnu/4b5g0EruPLfRcN+QHuIZQAcA2Ty64D24BgpcGiBxfqfLyxUb32vtbNTqYmwkmU0+4IWGUm
QeXccLTAJ1u2TqO955PVpanMsZFdDjjjkcxWAd86ONnlQmiKjNi+deuNXDZYGZjKrVSKe/8yYDj4
X1d8Q/diENTEV4TkA+WoWXxSWJjy7Yk1VaYDV/fmDRjaktqDq4HQnbnwkQmUeQHDKRGU6Ki1aY4G
oYurfUH1gfRUACCa1YXog3W4bCjQeyVfci7jlu9PjcPSl7EwJmDgeosdPMvk+fmWOhu+klHvzcZn
oRRJ231VJj0z5ld7slJXjibatP/aWIYRK7GKzUwNnhNZAL+X4Et8N6ShBIrOgjzH4NX1Epir5Nsr
NwuX+OZ2PcnRSyyloW27E40rkPQHYXlqi3rTK3jx+O/Rbxmq4TisiVmkHYxeBgut+xvzNJ2q1s8p
KfDKejzpWh18N6/tQ4LQh89d3qqDoGgxOT+AfAp4THM8SJL5bQpn26SKOpT9qSiV2rfKut0DeSfb
W50+QfrZz1xR1+VXnz0pxS2DbJQQJjZ8R4I9ZX9bwkgoqMqPzfM+4Cqxyph9pigw8Hm8EhXCMpbg
nyN5MiL3UhEwHP8r4Ecf4VvNNHp9gRxsSffKEOPOXCxaKpkssL+4YZc782IXhQRHu1WrfM4XrnXF
4ma3ZWcPWN58ryTRIbqCosWw7mtNxgNVSyo62PIpPnrIrGWt4LcRJal2f0VYuG6VsenRU0NE0q/Q
RvFvq3cEsk4X5Cny+RR/HbLa2g0T0kwNPZm2Ps8fWlWuo5e6nYu3gOWb4NrT5VUK/GZGvUv+n+ZU
djDrSH+DN+Mls2z2XhYIdDpaeHIQ8COGAZNrwfQDa4OQJBa03UDtjdGo3DVNy9gD3/ArG8qag+GG
DSnkHP/GcmneziDZwX8i6UZdJlZgeZUjimHdpcgRMrK4bgzS/GaLyCBVBuVVrLO5LefPfn15WaBK
7a7AfnSCdITOFs0z+v3Se6MqoDsKDKHOI9jY0S3svhTwxphsZ/mi//hE95CpcDSPvda2EguvM3z2
laJ3wMgZi3sntSitl+fR5fBR8XQirwq2ruQ0T8bqf6h/VHVnWc8lQ6EIeqjQ0/EY2vaew4LKrC9K
1+mbmyReAkKGubybGVA2ZizxCrRBZygH/r3XRt7RmluyyNhI+KEXs5e1/tngeqMaS2Im73IxK2JF
JxFTgWXZojiVZRSLFhnhXa8v5PNn2Qy3YdPAClvcebbh8GNrr7XxWQxA4SjIyeNXjG7UOnvwZz7y
4++QPUCeNnncnyE3HMnUmu8M1WyYiuBn8F7InF0LZL/M7AisN8aHiDpP4FAGBGoZ7i/V4NpI7o9M
Slp8CzMO3oNwjUvXu+ru4vdJaF0yVJ8BJ7zPLo88XkK1B9FKFTeb7IevnBWwdLJ/g1wOVCN3x8vM
yXgsU9PGjq9UcuWarY9zAr9yY8I6rq5FMQE0JLesTa4cXKxWeeelXwl08wfeO97TKKotL59udER7
+56/yI95xn9zqeX6YEUhxrKm1af6og9/8ja7yTZwtkVuLbpgs7aKFFRQhQW/T+W5pMdXx16Rp6Uw
CfgPnBlj2qqGy/Q9tDbSG+vXeGMlbv8wUl/4VVfgcvn7BczMKzG83MwDLHwDouxo8BjQaJUwN7Ec
MmpJcbn92nPZKoE0SDDZZbU7ujpJxTal88GsE2YSMZmdqViNdBGMoGQ8ElJKBSW0kPWtBSyf6Lcr
2fqyak6mWremrfFi5u+1+Ck5b3qitELwU2RnQu9NlA6Brzuf2nbdhdW7tm4i3dMJxq2Jk2nUxb7R
qacgD3wUHd4CJoRGxClOAlD7K2/ZGLdQkWLW+A0/B/d1gc/PXlOVcigtvehc2WTvdDv3RKzxbGup
yp8HnZGSl4BbPa75us0P5tLdcN3LRM1AT5otaEUWdHxDziYIYQxbvEoOslGNIXfmI6MM/wjq3YR1
OGlrMgGoYFJwtHA8kqSM5rWdi2Nc9T3zoqZlHLX6PQXAihJXNqSyqfT1oehOh+w4Kxk1a5OQnn1l
1Z27SvTwrFu1Wu6kowfpy1fLF3ACZy5CkM4PUIYGzB9xrkyCaHIWo8VWwzQH22YbUDY59PmDl3vQ
2Q3qABYKpIlblxHNxEnNjp18V9KxlZcYKeFJDkjGx7LF2oy8p0tvR+tPj+neiSKJpvq0+WjHfodR
83HLbIAtGj/+RSPXRS3077l1bynh5CuRiUaH9lsKEJiZ8fVx9SUbDlkHIcOvWepJUo/ckABqBDzT
HQfJvbU1lDP+KgUgMw0Go4/6HTfpTeLOT154UyBbpWk830EVaSGTXBLXCDy4yZdUELIQvm1U5SSd
am9J/w6pWU8jgAmZLvG1AttnSfBJfrAUy58LT/loR19hCvi+qIy1cV3Xjxuy5Tn6Tof54ECMFhpb
l/AqsjRNRTFKTWD7I5cqwdHxqQ83QRbU6F5ZrfJcjzObM/KifjBuImtiVQxJDEAjmcGaWPQ5aNHT
r6wG/vNPu28im5oWnju93IRdvMLaZmiTM8YRXN47xdEj5/fJpILyL0OCaDMAnZ1xcL+q7Dljjj9F
/n1xQ8ONdR9YUqnztNv3Sfv2afpzPticx50bskC9CWZGg/bN3ObP3hdvkyffoTnUcHFKPMKuBdbT
JqBA1xbigxsRgr5Uz4+iywf3bDFRkcnfoZsSoHDBeboL3TNOe6DVeJvNKSgJU1amwe/q2djajjxi
G9xLEer37t1TfyFkz3F/K8MMj2+gLMms6IiAnBiqYLCbauDXI1M+T8CkGEDWLSB4K6KYBS2jjO7G
0i0m5HdqjvzhYdodvAuCFfAMPlJO62hwjmEielwsSHnU0ijNCHNbY4TbvotWoCSvcVWk3joEJy0n
Spg3rfqJKxQnKn63mmL5PP+NdA4ZqXwou+m8j60tf2RfO9a3ie6y/jK8XmXQiVaM6qZP1dV9qhSm
MerEsoBpC3UyAobAiLCLWFCsVvUxVS0d83Sw2LN8Z728svBoPnLv5qPFrYkAhi4hjMvYzMIant78
oVA4szMsOxX6xS6g/youn1xhsYETHBMDZbjbZ4N+0+B7Z96mBnMisxM/CIFd3v9M/xRPvsNhv8Qc
rIM4BuPiU4XAC8HHG/KmhHDVmbuQsZQ6LRwChLhZAK6al4PvRZDR4Yaax1otoVJ305gur5NoRe2s
SC4JzSkwJNNX/cIVvu6MH7mWh3/UyYPaJw+ySkq2I/8gd6fUK03h/4xR8DoMBY9526C+YabAIYjY
2pCIwLkW+mc9cw8KwLbYD4J7Wbgw9clCQ6unFdF9jghu6Foy0A/+3TkDpb2360eFseI2iLVppU21
exJD/p5amh75uHNQiJZH54OcC1CRLikEvD+sM90RoKJH6wVMnul4/9ItdyfbgdG2ERR3VF9RI+Fn
pj/VGX7dB4UA2Y58N7FAF5UtbUFAGPackQaprpG/NNYgdTUsyCUjiOzZDMOw3RjPmRG736W6B6lg
RvTQhq7NGXmuEx9zSLEThbGkgWgJMekY2+ChWXbJisAbSAI/xOtAYHdUcH/z/05Z+WE+NMaOWn8U
IPu+brGbzAP1HRmpQrCGeBvVgUsm0X1EHnVI+YMtHuH1asLAqpNkhb8r6Z3upf6cENErKxO+PAtI
HfjFwl1epHsi9nJ4HY5W0lVg6V74eiFXgz9/4Y8S3LHWudrh2yudy0DbLA9uXT8wxXodQyKkc3yq
/+/9/UrM13qm0OP9u8X8t7ZU1dySP64YYCioif+psWSqfhm3TZp6fPxMeQCONzpsddOa1v1pknVS
RQCr3MgaWd4x8y5Q9pbXg93WcvLPIGUeWLgzBCYQTKnVYgTqvJX6U/B22o9XktbW9WIs2pQ1cyfE
VNHjEbReJm5RJo/MGZinMdVO6BnZj54A/pN51adV8A1xT8Wuj1nc+UJWHyO4DApmzb0BGMWDdXZz
RtEvbpSV8/plz6U8SrfZFCrD5AK0qUO8by+K6n4Emt8jXcumzKidoRTCPsmcVBoUUxPEmaR65i4Z
xWSgwzjZqy8NGyS7+/Ms+KFtCg/mREUeagae9jpDUvXmR6UVvN5COh0SWI2id19ARLmOLrer02rg
CcHj8EVlk50RYlQslzYxBYgQQ+zeRzSJGYlwTvVt5EWcEymfYTJplf6HKmaBR9nqrHP3t4hOHO6/
aizftki0NjyAG024zjJU0uAiiWwziDeE9Cuz5lGKrDrHS2ftaEKnzjUFf5radjzvCmUDAxRZWP/z
VljGahlE0VT1KiLOhi+FCBAHbLyNOH66VNnXUVxA9Hu5Ni94yWr4OvUp+xQZGu1GbYDv86L5Yhvu
p9pq5zXuX9yizZmoCipjbm1K1jDSpV3+iEz/hSijGHyEfNwqnlM66l/GEd/EXgrI8ZtWmE36PDFY
p2OxK/JOLz/5HVqLEqf1KxSCdgGRJM9o14VrzFjU+wGvUklV5Ij2lBYacsMvoUj460SDgbLRRo+B
BQvgrUWSUf/blAPZShdlc/aPVnRwtFSyVv5G3U6NIX5dSt+Ku35+7bimNgD4EIZ5zIlBATiUNsCN
Nr0dlNEiiy1O8ja6i+rcGsUXK53gkYE4l0MNxh5uuSd78U6cK/EQYtRNGitD1Rcx9OxphiyZOjKL
XDvTeX3pVhQQSXhJCDkQDJ7uNpr7mz6zrk0B0ywNg9Wd2g9g1FMdVcpK81l7XOKbxxlrucxpecrk
p8VWMLlVGNvsT0HuVq5rMfYHhQ1PQBBmDNYFHQzZrICgUcxi5liHEkzlyWtT7Ds0WS3fZChhoT2R
/JC3mhEEjBsP4z61F9ggdJJAk4e30RxvxKDZVTTszPcnek8VsW5YjlOfWQGM0S39D88PfEOQW9J0
Wg4ZKWheB/D3bhP08Xb76SJ3Su8xFvyFqoRAyNHwGrrnwAPFX+JgkYVJjg1hcH/UKBT9yopuzbc2
X8ONU5hOvCfb1SjOCXO+JNaiVmGM7xmQQa4f0Jb4X1ZmXnJ3l/Nu14/yvqUELVQwo133ZBs4xXtu
j+BVQ1A7claOpTcfdO8UNxjnBHw6XPpO0iWhk3U/3vr9MC/8nSvcyRaCPcdIN21QCfqM+OI7GLXS
X8j3kgZMCAp6DiN/69RLYRm5EZDeUgFrgZkXUA7ZmmZ+ezwU+KVFVAgt0wlr4MJTm1JPqyHO3uLB
w8fRPwYj50jYhgXw7F3R3J3qesn6ujAxuoE5TAEDzUdXywmbCm4A5V5qV+HlRlGCpRJsDGi2P0u6
ETyGFbDEgjPvfVLdLZ1Sod4bUnfHpv2rYLuuUC9kWZbAHBIEj6jeNFYh8K3CJbiSRUPGbUIENlLp
HuN3+m4FPkNT/W+qYgrq1PkKXHJVyIPdOau1qcwn6PPJAAa4dySp90LraqqrjBH7yolOctXzQCNZ
qLmPEvAhpAClaCEcufc6W969eylFOmhyGnCLE8ff1NEjWQ99WiBmhyEg++xblTjNLgQMY++P7VJS
GL9UEDz8sxGJxQx82qNznXh9Y6ApTSGHiCRMbVWXkwovxxS687By3gYuJHLZZKB4YiStyRws9PIq
9HsZ6QZT6fUkCjdA8+qm7DrjWoZPUUx5aaAcVfj1fmekrAi8SzanGzDI6IBrFgSBhocqlIJh9ABM
Xt95hlg7u29jBLaKI4JURVCexl2ueUP3sj3m4KvmVeKdIj0/kh/fvp2N5hszotGY1f/zOxQwvn/z
B431ggkdlGLI9mAbjUT+7H594BZJhA73eZTSzyrNQSBhs+H9buGHvmYbxoLG0Y2T0uEKE8DPCGxy
u0SG2F10a0NXTnAlP98nYSrXx6gX81VwZVWcPhUFThWxJZmm3S518IYp0lMCsIazmNfbcTBz58YV
/6BDEarRoaD/nyopfqFN2V8Z47AvXpPW5J738dVCQD/SthmTKL2FzuVtrg43LIcVOKkdY7tK/kJf
PXu/ND+z2dqUQx99TRvHxJxIQo1P8qEPw+277sEBxPJisiI+94zm5LYe+m0n/JzH5yvGOKfLxoli
EcmwUYIZbc0ot0GQ9MdltaFoy1muSEzvwsko5DZ0yk6vROyn2WoU/5L0ApRyWQ99mbve9o5wKUad
B2oNKj3lFTZRJikF98+qlNun8Agin4jPTAouMYmVt72mT+EnrDg75cLjZghlN3AsGoZXUYG/kUeU
QQe69vSL9QDPgMKJt9PDh1uMmJoyHomJ1B4PN/OyIr/ei/8oxaGbk4M5ubgZnD62KSxRFonrxFNB
+dkhj7Hzw1Ekz835iuUN8a3ajNnsa98l2gzlSKPyEkiJn8IUEny7ZAZCF2u2eW1ALu+6cv9qvhib
WMz5qkhijjpsakbyW+hIfagZw6hLDeVlPDiqD61Nfqt/bmtB1b/KnsPfjs4sJrO9I+YkwiaGSmko
WwHNYwdFY0Lju8sQwTa+OsyZTZgYpI90hCCY4/Jofd1WgLO4PI50OkPPK8YCb9RgshZvt0iBlxJm
vLahgb//exU6ApE1MtTr/Ee7Bwhj0zSTERPWei5kDl3qh7CtEJqqtMO815mu3wGgaxqmjAstvH6h
YKYH9j/IpCFTRoyBhkRB4m7jRrLVbhzqbTM5iQyqCWFZ02HkFmZ1iA+kCVTbVnXi802Ic2K+uEb4
PwDKdgkw/Tw/IjWsoZiYzgb9UwsV0dwaAfTfuRaWkzB2zeCpCUsU8YV5WhPC8ErcD5GXclCQ5LZF
88OO4KIZ41BXuN7tzSen5Zsf66fDg5EM+Hr/cEW2zfSEvwHwBOthWycet9FXTC9qz9OZ3ONIhOrh
yP2AJEqwKcEGCuwy18lXoP9aMey1XB7gKMAOVWvevRD+C1SQxzCaSly66L6QmMQHjawSaPlNLqaE
5zPwusMnTKjK6EZ7o6bnQ6EgBG4wnomajeYBFOyg5pUQEL/PWQ2QrAvuGokd8+gxzSjvVoE9Qbx/
uZo89ifKetPClpWh0LNa7mNYLy5YlKa73fHMJ2pqQaK0RxxITYN9TCbRHnwKGXuEmyHckXIsD4Ah
0BHPfTVb1hNjQn1Il2hoMk3NV+Hrz1RbgByS3QAVv5m7acyUedQI8I+39DDp9xJsdWsv1rB8Q2ju
TnNdhigSrHeVdLoNwSEdD1nBupOtllgDRy5LVnzLc6hzPOKY7Wc4FbiW956QtjbOp39MVy/i1K7j
n/s5pNKsv67h7cCUFYM0N0fGnhcAfRh/g646tqShFkEArSNSXTMLO43rKkPIohgbiitsFzIl/1MF
5I1bdBhwANNqwkgZyOqOMpAktZCABV6yc+dxAiagydRlx+a4kDWZ51sJT5xnQaDvQgDLMDECdZhQ
KNJv3xyJmsFAFFESfpbl15zRunAdZ0GFhNkHIWoGlnbFbXvD5BTVL4JRIZ5cHz0t3Az483PzPI3q
CGwQv2pk2m1vRhJVn+9/8jHX3huWpMu2uggwSV/cqjHy5gj6EuSS+AC2l7Pl8+/u6WTqEDeQrtLo
vrT3UkjlhQT+4WtSpjo4XSgzvubha0pv2qoDpGLwsQ+PayW8/ztrbs8K5xVe79ljeWhFd2esGGXc
9L7AE8Awm+GhMgk/jARUwM3az0Q3q0FgwWqxNYxYURp3ZMQ26eSAT3OFBrtgoJTZEO5FkSHOZcgN
EVwXHg0K2btT4qJPq1xmyMzZAO881wDewbjDbb71UkRwJoPzqyTqc/Y/CNK9SJMcEfjaC2eQ48mT
YUQy6qwVMZeEErZUAVs67WEKIOJDEkHcYlK25oEr/Gl8Zi6Dm4GeHsklwC/kBp4NVhsAiv/xK9q5
6SWv4xLvQtVWS1q9M+plOvn6JyJhgrYtTBaUmXFPIRc1NcrgbRETAVvidkIVyJBx+PPEKqaVAY9x
vrw2+HpR3JdLbMMERbFERPfTOU+AUrCc6oSAjJ1NP3zcmTS6scwSbAS3Y9pylmLdpZFdaP1Oix//
sJX0WVKkwt4aaZjxIWSSs4trLWs6v0Z9HfCBXwc/UjsjB3taJJ6seMO9p5eYj92ssOP4OzHaYaNm
iYCHajW1K9R8bKa72qTckJ+x0ZBRP/OREczenzof+0nkuLE9iepK7zPriBCqlka3Fbf0z3BOos78
YfMzEWZRhFrDlX2TFnz5AdYV+r5+/CA+Y82v0xukbij+rH/Do0D5Ze6mhxYxB7QIadrgzozQMQUT
vWtRAJB4VB9tsxfyOnBva2YJpZKSALWuUYYQwzKmuLYmU3da5PcZDzk1uKDEWrGbM3bMjfiv8EQe
ml1pYqwMwDjrVl49UbH22L+fARN9Ud+v/iv0cQunirxBlhFQ4qbLhmaR2Iu+Xwg/9DVp3Z0pK/mg
ENnj31JS0ePz756dGktyGzUMcCfpPcVk/bffAXo9AuGFnwmIDkFxw4jR6S2JSTIBcf91Gz0yXZFV
1MLLjtfps5Dw+EgETaLTY0gB7VXtJdr/vF9bzk56e098Hj0qaP+6pqRmleUEEYs3s2RUMDhY0yNo
qcKvbk1yVD+xTpyjBMAkMjYgt+bpiLmmyc//0t2jLuYHh02GIM5dmduFbd3bXEGb44kRoyGjXFDT
FJKCuCJc4B4bNSUtFpba8FNsZfunHL3Dq9wyXujavLdiC241KygohUxV/hmeYGfH7+7j7fxvtAVI
2OqXHl7E+O9YJ4sizDpdFsmmSDzUvdLDIqjik9gYlHEruOQKcvgp4j4G+wP0QLpxVmQove6gEwYW
CWehV8+q37ztKVm6icjej8xbEHx3YhMBF+3jIlF6VP1DAm5OG2P+1AUIu+GleiPh7NjGFlmRBUya
nT4xSdtbbgENQUkIbmqLg5B6Is7NmKNQ0xLSZdiIKTx7F8IyqW9Jy0oKhffpFj6nEq9VrKYiJqUU
fks81W6y6CjE14FQojBmT7c+KpN3Fb9lCsy6lWWwgXxYWF0nRqTq9tRVTAeV54X/H9eoESbffQcm
8iqB7ocMoc5sD1AVWQ18NnX+n4CjCZsVlKjkC4bdg0u7Dn0J/zofrIndXi0NIdhfe3pwazmJ3dpT
pUDIIeUs7wryFyBxU37aWZ2rf191d9dEtpjxfQevSr7bIwU63n1Kfj+uD6n4VTbiFszS+KT8PKqB
EpCInI8JQR40l+eMz2z83T8ihrsfQHA77xg2yetY9hlm4bzU9wrUNEf8rzuN57oQXofLgvTsV7Kf
Hjdms51lj1zJE3Zw56eCnP6HQtN37zGsCc84xihjplepgZC5oZWGZQqfyvXMXPxEbfzwXkIrzvk7
oUnLaxy/Nt2NDmmHLSUhuDJUUNH9ajTwGLJcssrR7j5ITqzbka8ZlT49kjyu6dQe/s7xqzzZ2bJ2
u+j23TFdZy6j8CVRbUb9XQjSQEYRI+RP5pEaMtPscw6iM46PKUCl+dOmP4bY/vjWoxyOcd3h6cQd
uH1oHjG47Gng7bZVO0Z+rl99bha+ph2PyQl1YsicdvatY1dWzTiaMTvnKCP+P+P+mFtgSmGW0ABO
dQk+GyoEuh58orZcQMRws1CrzTAz2DwgDKvq5DsgOmX82j3g0Q7lgYQblRt1GBuq9Qqn50nfOwKT
tVi6GgZUgd302a7uB7JuvM85AexOuKU56zpGbCJTbwl1b6GzkaK2VirKwLIn6qeDxqg9uKsdnUgH
lMXEKGLwXyNOonHZr22jIyfa88RmbSAD97L5yKmriVWCO5+SuKTclebqWBvu+HuTz2pVafgqJYsk
e9fWH/P6oQGZD5oFEK0cEP7QSId30xgkHF1q8IRdnkxv8VwsfMYjwYUwTsZB2t/AYfZpi2mYfEOm
R2/rGLoMhQctbz9ftvrkeSMuCyVuskkBI43VBxGXZCzhZ+5JQ4GIFL7i/4fTv4CrBvO6bjTj0CTj
J9NeDWuhUKlpT/SiWMXRucYDf4lbosmKX34/+jdDs3TjJ/tI56hZkNwUFqhNLwBjv/Ll58fVzBYE
NWIg4siZBmBUffr2mkUwEsOF89ZEtPxaSEGEsZw0nYXfR+bT8cZtsMBsg5teYSmYLmqoZ6bgJNAl
5QS9owtI6B5STWNGGbtUB/vvpsyECAVrIa+co2NP5dMVsFGYszmn/rK8tWRlmK9IxYTE6pORTHOW
G0kk+BOEEuDf7NqnRvtja1Kzxt+ooVWh7UY7oRzAaPkIPaJ6eZXnUwRTISg40LxCUinq42yb9MSY
MDpr8ErrpbC26pr0156+LP2iJV2QKFdiBFRmwB0ToAzZ1uYr5JkGtkDyJzjN6jB/JYk0eJFeDpg/
922dGfwtz0gqopZdTGpVdyXqY+63cZOJOLdr6U8GYqFftM53YlZ7VrmTW3/nJf9qCbI47tEpveDa
zqpRF6npwncW22Q2R6tod+9kptmEcJfjZSCVFg1V/jYFqX+7MLhuYPTwOFU8cSWjU4oUCvF8xLE9
ilkl7NXoTOhSdGyTDrEaMiD8unc/ykSmvKoQJRT4BFUBBau2pod8mulp59xG23YRu97vb3bjhfna
zZ4dRq0pLw2sX1nBVpYrNfsxsjjbWHoa+4AZsx1bKxudUsG3k5dEL7AUyR4o+1YPqtFow3/3QQst
dHODQfz2URbzTPTHocx7/8wLyB8AHjHokzKA26YTs+yfp8ih8mHGxrEb2fNMeGbLpwuZjz1qz0Au
Ox61qJtNMiQxPSkjLvqeOhwkHGuzHsKNPyN9F15YUjPsWw0Bn2vQI8/zoAhA/+8BUR60KeMc6wzA
amzk9jImI61x3kEjwFiUS5T7qc8lvW4hZzcpVuCv+M5ulAsK1IGYUMwnabPwy7lX3SBfFcrw4Bzl
CJ6Qqzt+6dM5nLfQjoI1Ay/3aSijq0HqUYzRMS6LxHKERcBuys2SWr73UAFs6akm4Ou+zRxMjIgL
EtxAy6zcS6w40lihH0+izKpOoIguoVgktmDk4OEEbo/OGh1Gk4optqnyi7MJ15FaIiA+6oDARs4s
lRCP0EqGBqWQKZd9Ri/x9RdwUsWk/GxPq1VaohWTJ0FJsHTZyZvm+d/q14I6wYEphafSb6zZsOYM
71UsFnIMQ4aNoTN6KiTcXT/T4yNBRf31/sdO9TqdLKPW6ZA7mo/0n1tSHe7T44jxbsruMBRHDE61
VJouADLpxDS27qu8Mh6QZ/2M/pb2qkbBn7UNyNIoiJMs7nqk0ofGeVR7fbwCRkrtW32I9kzpYttp
/SuEjm45s5H8OLwbR5c4ps6zxKVGttd2IiMqyp6JoYOvysA/kHPG+3IOa7PsOo+01YlvPEllYBeQ
LHU78xeWF719Hwo1A6WPDXokriYa4W2XtfYybpq4L1vbLWj5xITsP739NL+iwYiwTqgxx7Hp66i/
kVLN3HrivIEhSVBp8pQGVXgAK/uJnQGa57phwhU5mO2qoXEDw1Z37pG+28SgwjNz6Zh/K0ISrMHE
psEb5pPnHNz/rOYYPKGYidKfDu4GX0GWu29PEIxN3DeagbBtvKxMWAecLTk7Ln0CKCLdA44Lkzgx
PzHMP4hFLFCkJp4oef4hz0GWbzRwlAltBq6iXLxlUPX6pmyFXlbzEmIFQZaxPM2QCurcaZgFdUO0
Pw549n5sM2/ztvXr4nyRrdX0k+TIHsM6RHHRHT9Cx0ci+S8TMwJoiZQanxpmpUDv2hlRUiQsxZeQ
LUP4ASFjPz0qpSRoUeFYQqireCjrVcfAEKY8eyUmbkCyW6dS/ATFD0hwu/cXdBgn8uDMAWZVtwgN
U6as2LycSYU4eghbw6qeiP+lBn5HdxYTp2eS6huTSaRbrk6qUDQAllr36Uy50VW1YSD4iXfJ7rF4
xr2LEXsHEy2YjO13ZjVV3BQmBEJWQRQqsZE/GYml/UR0OYocc+gBzz2/imdt8n+0tc7nYolOBfTi
GChPOIn0O4XQ6vSPIs3nH6GxK5FqA32eojOLr2Txolp63ErOxYh8kdoxN6OGS+f+T2O7rmvNp6Oe
vkKAZRnLyQ7HKUFXUgiEmJO1qdQC/nXR5BV0glzNRGJoPzpRZx7axCDHy56QLL8/GMYhlZbLrnJi
1wmRygjsyB4tvSYDdbWEGG0oJ8PdBbTo9z0cp9CQekMHAeH5/z/kjEuE03BUTt3JA742a4UzooWp
CaKTfG5nE32dE/uSwv+2Dak2ngvUd+MOBxh1Iug+0Jbq2h87Y0zD3vuQFPU/RjdL1zeXgRA5gcco
/RhkzUy6Y76faBCNpQXFE1F34Xnnhq+rtB1s4jLP+D+NS0chjBcnM+VHhM8KvoRl0Iqa2Ilwc04e
7RyMtI8eI8Dmuns3SD9uOT2kZoRuxJAr0wTXpxnm0wIBrp4XJ20p5I1JheWn6HMiamykWL1OxwQp
vfBK3c6bwoia628YEmcHjCTjftYcTVrwwbuN7uQ/P8BUAxYKUmgA3YEqazOi9n7+6G/mZryWx32P
6lVQHA54L4Swf4EQuolBx3MFQYC5SiQBwMp2t4WHNeAgqPalDX68XgkXGam3ui77t14Qeu+2eQuF
LeoKZBKHOR4aYW8k/gAbxy6rHVB/07Nd2ehmH3zVSaOEPmELR8t63ZNknOQNEIezMETJo0aBxutd
o6d3B6qRMOiur5IhHljSiIbIbCJixm7u9wQtiXLmym68PvZt/GQY6oMzUr4A6kZiu+KAnw58TT5y
bknZwaqL2vq4pT8NnV9ceH4AVeMkdJqAj0i8NctK6AvYhT14zA/jZUKkhi/sfoyor+v4qZY3Ua8B
lBCwSyizk08wxa0U30f2reDPWCh+QZKaJktHNbyJnz0LIGBXOFPnrqIUE0SUSCPaAf9H1MFwYjk8
9jKMFbEYvtmhhmfXWan5YliQHwYpU2PyhhWgqyXyGFvnrECe9CfQjdwHAKZkgdN+72jOjuLb+Eh/
kjZg31Y0sYUCSwwsIQXukRZYCZVMBFFleQONJXTRk7GrVllK1c7ppIQPgifvUp6PxFT4F7+LSKmg
RgHijqNwqbBPnBpzLhsy+KljOZJrmNBbu9yBOlkNIYdksoecLzdOf8MlvIWWBOkHUKZ/U+P8AXy9
5tFuj6vqP3pzOJSMe36eSpxNjBbl/efDkXEznmZJ8CrwaflyztbpyhTf7Iid/ZuUC5kFUPhL5Fa7
nrblu3DdmJgUrRieYfW47Y7T85Pez4a0KYu8S9/OkxtRxCiU2hWeLpE/v49aAXEFogrM4EbMM7IZ
JRkbu6S+5d+vniN2w0mBL6lhl5y/jNvm4CQ+z/9IXo/TH1X9M/uFPdqV5mKy4hmJWKc6baXYnu1j
fEVob43f5Y/YXXTgNON0Km5tLFsru+MyJM6YWYi70AES9gGyUke3c4ey27HNI2qAGm6zsSKaBu4l
W8GMTZdhjHXD4ZqXsl7TQ+26XhFl9OsQCA3ewf+1Y0YRXh6yPXOn6nGEqZqruMU40KN4FQ+rh1Gx
Qc0GlGLRY2ZLbIC2iiEVAD6FI6FqsE+FDqoOtov+1U04sHCncFnTGtsutT0x5auMrM0NDb9p6V1b
We62ERYfYreKtRmbGIBCtnzZ/9nTheZ/8/xYuM8Mak7AeZatNVYI/pmya3J7HVAQVl6/YfpK3yH9
pSyC7MMrQZZDWDvXwkt48Y1Z3Z4UWfOptv9fy4Pv5HbqujYgeTzhw0CXYP3GkwqfxLbQzKHzzSGT
eHm3nhT9zM3nQbZkDPYoRv9hKCNSqKjXe8+vLZ9qhIOTUnpHt0nU2lShS2VHb1X7MybMl1LYv4En
y7KVeS/nYJdTCJq6e3WPMzI9feLTGu+nyTlY+b7+0A7gPs2mvPVdfiveBHa2iWk7xyE/r6XSvKvh
VhBUxz45k37JdotcnoSTotpxca8CNUjLffQMP7dPwalIU7F33WwU4uK0iwiFrpVL1/mOZ7FH0PCx
ZszqaZX1z6S2/d4N5dxoo2bdalnp5VaEAaT82LkWwt7cuKQQFNzL+R2Wr8L+dcJonE8Ypl2mahT+
1NdCOmBW0h70w23Hp5yAuTYoZdC/sTzlg5kRBhX2BEPMYbj+O8UOEIfKwJItoroeMtAI9LaF6yIj
zGhC4hIc4x3YPaZAwqQaKtfydm4Q9lmTWbD99uPVrwRDo/qtYyImzqMwkSNesidihE1Oq2SscNE5
whsoGyd/TgRsvIRLFGDnyjW2z6nU6+lsXOoiLbtZuaWUGP2xGxsIV6L95qXvGpIiTbLrtDsMEeCh
0ZP2npvXDZZyjBXqpso8gISQx+Gx7H2TcUYqcpJwNBQ+sFBXb34J6+4/DYk6UF20oQYPmM+Oj44B
ljh8h8Xet6v/bG14wJHBjg1o4IrbCUR3l03hf3W9XFucmBlBKzRi+19093gkZfD44QmslPzp9mpg
8O1fMrH/B6xsyq+Scu3Py+aN13dKA0uNO3hS1sM98cFQzUVCcbtiMwVacy5YdcGZntXah46MagXV
SfqxXYaOL8ySBO37jXNN4nHqEmbUjQumKsDAgWzenkXwB5TxbPkngxXl0ftIUveHgHiXWyMStqaG
riKEBolklzBYot8d1+sK3jLQPCI72wdqUnT3JLujlUd4oO8DaI4xMag6lAr0elei00YMwmkiK0mB
SQ5ybAPikd4ECfXMrvK80wYOEwlwqtghbls8wA4t/ocpYs7zZ6Mx3nGv1WlMkxQHUkAWvcp9yCEL
3NKQqhDp+Oe3SAh5h60sZ6AGfuDR6+72EOFw3XfzaMRhrG8SR3d5FJ8JSEyYgkCnHdYzcEIy2LuS
rYO2mEvZ0EZxjOxxmmhZLqRg3m3QcbVNjv1wBa2wnWaJl24m1NQq2gsU9TTFRbzxlgxbT3GxiscM
sBWkSji17zXecah0Nk2FmkV3/8xXfCxejpHLIsgin5mdQNFaXXN4R2ykbyClsu1TPuN63Hb49D6Z
2bY9KB/Ao/PTehNYWcOwd9OMNQoLfoNgqIxtb2Fe4WFblOf86Iyj2ZezRQ0thS2o+sQI9Cid2Bfo
kHg6M5b3VbuP8K7V2uVxi10ti+pBieSpzZsRmF5AQzwU0fEQde59iaPyQQknCmdpny9xEoLJxwBa
3VZ8LLYT5fTNSinkevTXFFFWVYyWvT0sPZFyIoARfkuEHn0nes50e6Ev/zP7Lv4OQdpqEe2z9P5x
9kNV4ylOBPPj6fygztMCab0PfTb+JokSvitexbtAkborlqfGx2WXxis0d5TpmjvBU93KaAhLBj2G
0dt2kfHZZgKZtQHGExHeuS3oi/0DpbHbRZZU8N3LjPRuDZytScSS1THlxwJEfUM0g5oj4OhxHeHy
TaHPgV1JxweAS2UJG9LXgBPz2lUF9Lnip7rn4CorvIXP5ovak7soI62s/XEK44AYAtdZuYkVwVeV
u5SJgx45XsiTErbFJUIcrDcER77JSVv6jZqQBQczqOu45xT7lpAZvDvMII2/CR40AcFm3EFuf8+H
mCcSs0DnEglBd7lz43atuIrKhpOH3Ca4cIm7dyyg09GSz+MVvbD6+qjYodx1Qb59KVI9PCAstGQj
vWn96X0NVHZYS0SmqB0FXTUhqOuBKcZd4Ijzr9o5XDsFTphTyaJlqCEsAgEmiZH2leijAqRRcRqw
d4IPi0/tHGNMZ91DeZhRrvOqGs6lbQ3YB4+m1jdaSeH/WP3bFyMBAZ9GSfz/yb/bChajUIV4xkD0
wqDTOl/+vYYQOmVzU03HBUUtek5pLaeOdViDr+hZsQIeGBnzpHJjHJtM4abMzHMMrAFnUqctXJLB
mPH17iVdS1eGxX15O9hHUG0uuuQFyy6nGbEC/Vn/Jm6rCugugVW3/KZRC4VwZzZpW8pTOMbUu6eP
85BQ1EJBDiaWLfLjbPLkpXmIclm5/hjy3oCLkGKU8OtCAQx/tnvz1Zk74JrnD6HugD6cmHhqO2IO
9KT3cBUDV0LZ71i0MYuWoLFRbFimlarWLoyfXS1xBTBe/fND4YVw1gGDZCtbkqbTDTwbXWxQzTk6
Sq6vW9NN14yuS+p1YpLlbousFnTvJY1KLBtznOOteeroslylv4VnfKX6pLysLDRsCFNRjEe1oyQg
ZFb3v8cDj/H0lDG6vFkTpUTxB75X+jxtwDtveITnS5D1aQdihU9/WK1rE9TLF3gjavzhZf4InEyO
85tu79HSrecPhL6zw/Q1vwCHyPN47hUGvblUv8U7wt5v1i/hQNwr+FFoeNDD/J68Bz5rQT7xiFqN
x64T4ST/L6m9qgYtLZbu9uLTxm1+5EW4ebkdUnv0RkJSwvSvzV1Vj/3fHiQQsMWae0ygzrwOIgbJ
HMahuNGyMrHA0SKDIPBYstBbTGdQcG1CVYJMLLZYiLMEBR7II4r+x1ahkO5MvmESeGjoh4R3km63
WkGH/Nz5HJLShprSvzouEUo5Q08h28gVIRX8N3Y1mwi0h+OGeffeXzGUCI0kKNkc1tFnGSSxfPEV
C8kVVEVvoaWptAjiflsIBMbHsUl4QSerCiEs3Fml4aheQ8FpR/uLvz3I1dvIWssQd5uCBivPqDAS
dJokKJEv0TnyKjcMbFomDVl9v7fjmMb4BezyxyBsviAHd7P5cz3ciNQO56yfMzj1dT8vmeWV1zWj
cDR5MEVVn2kEKR8EqbY0ZPYcUjdiABfH5pFmL95I9Sov34r6z0+z7O/tNa1t2BJp0G8AeXPdefLK
zZbH2W4/lhfZuG1QHqQZHq8Kdw+IMSJVoExyW2HZWL2dhCg9efFfn/QTxd58do0OCGnEiSjDWHVh
dfmyzjfVw6PsEirkWD4tXXzlbKAHIRJZ7H1ELzyONaaR/fYHoCTH/i0BH1j6s4YagLwJXZAoqZar
PcTQwxPh7aC0QB6MtAdWx/aZDdSbS6W7F9sZxITmuXVOpfDwbZSq0DxGV969NK8QRofhowrPyRXX
gdUpMZ0f2dUJt0/0SPUiEbUBGpC4m3JP4mllehiB7VKcHxqLdbj5tLkTOzDkUjMpaznMWeE37Qmm
ANM19DqlqgNQuFifWt+nU04iNxszljfpLhUcC8zpw1qruqqrJ2nG6L1PYbHPSj1xzP3tKRGSFHoG
/KFt2P2dQmHweirVnVNQaunXLzheLsI76Dqr/XV4wjkwzlL9dgaVkgaQcpZBGHIPgWSen3LVMzAU
6PPGXWBpRkrMxDpdlnyyL8T9UcN0BMA7JR7JhiQGCXL2SbaS6X/iPw+NrsXbOJubmWwwfm9pmbxb
FctFHV/RBoLkpw2FH/slO4MSuuZdP356nvT/krhmmEFkg5owXx1yMB3VVlMO4ihu6qPiebIqo5Cd
4D4KMf/KmHQyPwWaPAjfJeb2SWVequB9G41qzqD18QWZBaDs9kjH3oHMDcF0MSeu6AUMmrsMzaoC
sOVXN0jqLHHANV9hXre82fg0pwn50v/prQH1IjIezlQda+YzminVX562LnIpRYKzkafam5mfMRxg
+on/NTarf4rVgLjeVFQxpMD8iBfj3L02PEVfqdIBgrr+i/pYGzHjFEWNrHsdN1B/GUcdEAJ8Tl+s
VWdUkmGRai0hry7d2TA15JGIsOvO0E3QwCv2+dCqTt9EcjFFe1N+gxKVTRKA7L26eUUh11EYglFX
UrKjiU0cvUYIwE6KRSeKi+dukTVT/4yR5+n6CNYPZpdNFWMGXW+V0/RZH5XjC2bmFFKeFfILQ5eo
5swn/IisTo3mMcGJUh9gOQDaMMj9d1I549wTIur5Aek7uScMDfKuN/Li71daizsXclLc622s+cDT
GdTOSmJdikTxiPm7DmmCtEYoIMfUIOLNAaGJ57Ed9IYx+w00vuZ2NUhL0aUbuq1GBftAWade5y9m
3mA1A5Upq5GOttDkyh1ENgwR9g1oM2o4YnCBmSqP3MlmwOS6II4TV0R2OX0XiNGxWtOSoBFhYLxA
ji84XLHf2ZoTx+sAPbcn4mBMWLyfy6lLTmEFcvtfRuXYEciDvy1uGCoZNLSZJhF5ikB4vnv83IOK
+N/gssTsiNvTpeYjaEUuTApDF0I7lcM4qnnNfuVG7CUfJrMSvZYvQ0FP7y8oyEawj+YkJjjGlhAn
4zHV7dR9Iv+9tXdcKrfd9oujYECDjBp+vHma7Vzi7/JaCrWUwint0EEJR2+JHJ652upjBABQaQE2
wuXMCqALkd6To3PgmJcMOKIC72BQNwOOicGePw50Nz4HwhzfJqCPprg/D2PWAJzjimqLDpcwAR1W
1FTBT+Qi8+LQjj3rAhR1U4kszTOsxRvTfcEEgPSF5TH59WaG8DQ0/8kxi983Ff9K5rGsA5d7v5qr
QE9shhZSRcuC9ImHBIKfI16PeMu1C+eUUBSFOfpdsAEMt+RlaWwqEz1ac1vlPlIor/M25DJQyWPy
z3NZEGWTGQQa81Kv6qWiqS6PIAzRVmYWinlw4w87IoKaew+36ZxKfRzhBp7tc7YYEa79FFWFjhZn
6hlRz1eC+7DUTOYygMfpqU+OACA/3xmvV5Bj9ItO5x96TVWiIAzANsqJh6xE7HkKIIwyFZ2VgDZ4
0ys5/izfwXygO0fFeBfXtD0s0nop51ttVJcEpb79vTcm6Oz2sYdhEteoY4I0chzLrgQUqcgLIhFb
eleY5KIvPShXfxAiQmZVTXb5z1IHDBRhgt4PLJK5KIK0w4uN5iXZ78vCp5gADj/2MSN2GE8XEQNo
uWuv2MZSeFNLPA4/9LN3k8cZCX7qtObhkagzpDNoNNx+QFd058DuiRJarpmdWwDtakRAvd0sryVC
WM23H8H6RIU8FahqK7ZZ/wfVLQAUoUo9RUjD4t4YSfsZQaD1DTxOA08b7e0324VnAUHudicoUKCB
JBr0KR27wo/xBE+k2wwJDxtl4+ybFSVrhLAlB2IM8IeALmhDXvqcDbrxbbZoKJiNudnbKYxgZtVP
+Zlw1l0I2K/TsDn6Urb2pPafepaL7Q0V+064G/6PgQ6O9sEAwncmEs3IzoMLZOL4W9z0RI9AFftV
9cslIyPEvbyEr+kLmxD12hwmwL7IxQKsSo9wpKL6cNqCN8pcMD3+2gnKPCYG4eGKmDGHGfcuYGwS
xXbXyvfsVDS1j5IRWK7X/Dne6qWWDNE2YCYG6AzzPNgrC0Yi9UBCYZRgorZepdoOQlpZxCRTxfdk
g40IYkodsoEZXY0VN82vj/RDpvotk5k59E3ii0IniGY8QXPPNMPrSvdUTTUltkxzzj5DT66zms8/
B0Kpalv9jbhyJpHgQMudQm4yNGgJ5PbMjJd4A0aogb+e/GFRQ3OH+j9hu7F/voMpWd51MlLKdsjw
0bBTpvV+gNS1/TbTDsBY6ZnB19TQlWpT0TY2oiwt3OwRZlzh2n/hkUc4MmBghr+LMoEmhX+EtqRm
3e3YJNg38NPXHWo1If80SbY2NNl668/tlXC8esjCr9ZS9RbpTfWm3+3oryvXV/DUvj2DE5ZNE/Jb
LroQLlS7u62TTIj7AVM/ZrCwD5xgRB0MP9mcRZpwaK4DPwrYrQAYeQ7dGPxPHjV2JA6K0mhZT672
YObnGbkCj29l5BEc2ee0gKIS33RGAWFSyIsr745cVKNKuCcO49/qoD+KKacmobDlC2frZCqlFDgs
C6JjqxmlhksuI73YrWJ6zP/ojtQyHeWbqlP6PmYsu3wq5QjNXiNuaeyXr5CjklXxI0uGVy5nQ6rf
ElX8aVwQgtx6HSUEn5Ks3IpfqMUCUOvDEgf/YIRaAyMrcq11J+vFfsGAu+aIZgrq1EamBp49hLD/
oLwVy6CxA31m37Ay7FlQKRJOSD2o0u0p7kWfCZsvWTMjtodmvVUBmIaQmdJEwUajztC86Alz2nqN
yV5dBJD+v/arlX3FI2dEJyWPd16+SbxJvFfXjmpC/cCtgHjOEq+aBgJF+c+byTuQCs+Y2d6+OIRm
aj71W4g9QBgxSRFbkXaelgkcEdQWysfcJRy9+Q7lfjC5eB3pLbHBFMQwb6leuK1tecdhOBWBsDqA
PeJRI74lS2T7b7xC3Uax6hVxLXHl+0bUS/gTMBhO/RIRztZsxAM1VKWUslaFAY7I2/iyNc7/A/w9
hA4Fzb/gzwN2wQXv1E7eETP+VKPHvM1CuhCb5Y22fFbB9YDk04eBwQ9tQvi3jxyZKN1ZK4dAYS6R
nX9/br8ze596KljmF3iuBoym8Va3XSVQ5qFirmabC9s1YOv5D9ufKinBaY/E9utIRxnPvhpV2C34
4P8GFQW9tlHEiHrZ9D9qZo4lWORXkD6gNciHYwg9do/ThRz9PtKywI2hIX+lzA+q68wP6yDUyO/w
Fl+T5ZHOlqHVz9wLaY+Ihovi2DkXI/1otEBB2PiKMNDHNRe4inEqXpcvVJCwzPhvkrhH33EM4nDK
mwU16isnHWT2zklesw5x5cqGNsL115/eszTvLB2tQfB4ZwahyK4oGO8wf4OVD9ezfTEEeDcIa6NK
m+IIGQMzRMJjxz+ph3+fprH8ril01GWWr151W/ngmzIR9Nks0JDNH2bOz6loh5XiKmDrS2+6E59K
xq4xYYDL1HsiMSrJ2VeGz8SEEajRG1ry/OmP3MxG0QEuMfbK7GZZ3eHoQLjQN8bNJaZRUHvaBQj/
Lk8vuZJe4G9jsg4ExkX8jF2YtHJEkkpCU7Dii2RrwM/0odGJpFQioUHm5LxQuZUJ3QnSF5Wv/9iS
D29/ZWDfyOZOKEcrNbRHH+WX80HZdQ324AoPJcVieAiizJ8hy+hqdhVdChcNNng34orW5rr01cjc
/VR2T0XOWZhB8cxEpc1991m4EPDCj3nFPwLdvWjKORvXXeQ/DTZAVPs0zwS7YZWLYT0KMchp3AuU
v/TZMafg0hxuxNnB2VV7y7c9iHthMbPD00WCgq0C5EPTAlWx+E4IOez48XLkORfa+RdKvuajoH58
ozmWga0mJfOyijrYIe4af0dsPLohqsiqfLZVm2FKVDjRwT7Px6skNRLoNNV4Azxz2umY1OjCPwLJ
fGzbtcavjLjcBts4hMa16sg28bTHWsMxs6R2CcV6CdHjtDZqYE6nXDlfWgVNOyP3C1QU81LbHUvM
OZjhjmwZWupR2x1fXTRugG4C27QZxByqrme7uEG1jYDdZg2rcpzB47gGJ4z5gQj9dGLPuB3XdsGq
gWEj0uvVHIdcslugFTght3BInIksroeC+N9bTqwtLV4dcDM4/bCRfK6IQt9EA01VJMbg2iI8pUAL
BiTxRkhi7PE4Mm5FeB1MxvBOnrBJ/nzymElEp1mkEk+9advZbZVoWoD9UFMjiFBADHVj9C26Km/m
+26ICcjfgurcIxRcQPtpxRBKZRAwun1C9yLUEpc2O8uHWM1SNINmDyOrRkbSQQxnsj+BEDS9ZARu
2aSEDFvHuJiy9xYxAVOoAYgRD57MtF78cxLsLx8p5JnFa7Cb6hJmgJXavXUg8Xh2CQdVYnJF+9M4
k62VaKJncwZwtkdd/2t3omI7AT8sulnB/dKdbmxbIE9gvM2uglSNTZCooS82d3Ub44+eUDAnheGS
b+aD/10etNRY95SWmLnbmT1FjSgnkC8eoay7n9Y/EBiWScPAK1+plabfgZfTkTDe2fACU2dxxEBv
03gK9173CbPwPOlvuHdjCfQY44jdNRmeSlraInE69qsLQleab3XQbNe+ZYHhkRc6A/t6p3rZlA5M
hbHxycDSGQtmuRDRpwiM48jiY2nC6vVgfjLgp+NWRjzWGKowvttKoDS0J4jO1rGcxZlELZvI+4k9
g09+3w2dxbqgYjEEmelUrNrMCrIqUS4MuAQ1ZkGqkOW+zFL302YXJgxbNZaelupDAAMWt9xfHXW9
+phexaimN/EiWogQT4kwnSey06Hflmstg2FsQEjV76+Ghy8AoYuKxZCCfqo+lzY4I6wlTzTvlTwD
Hqy7kbP+DO9G7WOoN7V2zKCWarql1TGDCJZerv/eOrKu0nWvpzzjWsVzf6gvs9Qm1WJwN6TCXnAB
2eHWDKySeADF6DXrCrgnPtv/S3W8emmN7nV5nsRTp+Tl1AAs37E46Z4s3lWBPbJsZb90LaEMyg0t
3LQ6mDIr2zBccYESd20nLuIYwG8IWMnAypc0MyogrWg9qfIYrGevXVxmmW2R0tixtYG/NIFMMtgH
bRJgsCrxu6OmHuUjOr7G9WeneMg/QEFX9K+7kW0XqilmvsMI93QY4mLcD4Lq19EQhqZYqkcQ0sEx
Uqp0tTdZE8Pyq5vzJ7v2CSbNPsFgC4f1apY8fQ+atUVcIU28M9rvE3esxYHttpEo3qN+qqRW1pVX
J49D0qgAUyClIW6yVNL9f0H6qHh9bsuS/xcfUiX8sUxTHAov0GBOFPyRxvU/YGe567TjbToLU+az
r8LtrvaJEF5gD0wGlO1ob1jzDJLZ0/3jpQYtzxEmlTOTPUUuIpv/kvDFXWxnHeJ6oiW3bCzRPX1p
UkLRYGoogX0CDQUG3kp3nMauEYKNiL7a5JIdvpuWW5Sm6WQjKnQFj9hKizzLLJXQJa5702+mDxgb
nhtEN9MpP9iIQzGNRU4s6Cp8l+KpCBolqZuhrd+3QnAC57PUeHgbcKC9kO/xmblWiJiBB9iHKPKY
kqa6d1F/sSSG7+eoOt2HzZKzdRpqVyeO3Y6xZjaQLenTRItyX0FKwbyD2AqFtbDxmYOM2Lw1MK+F
zHYaXI5C7SwYmiyr5x9gKNbKfwP6UtVLflpW6Zxa0w5qQtujNWeD7BxpMVv7J7oYgnyJ6VmDqiVI
xeWowMRyiYYgLbdXXYFXJNpcFCmaMfsm13k16ILr6+YBxb6aohQRTgPubK6n5tmb/b46MH/Kk6vP
dMlaj3FPzl7rVqiw1d+5UgPzl+FO/4yZNh9B4ccvvxojs5jhM6SfQtT7VdzyMrH+0fBrY2LE8G5a
2ECqe4dpe5igBvLyqjYqwd1iIAzXjXLmv8J6+r1jzUNwtBzfKffIBevwO/bK+kupPq78bworNc2n
H7P6V6Wi2nrpvMkNjPdRAl+aip8dfEgqmDKyH0bxxwaOIqLAue7hBsm6fQixAwpKxS4sKxSMF/Ql
3lR10c2qae1X7Njb3p3xICC1QR1SAWgJ3j3V1FN71LMYixrNJgTlCd5D9IkAQVfBvopnVl57z6wP
3SEn8aGMNKnLnUbpxV/2AD4q8st3k/S8ToFDoM8CYAAMg7yO3fLUatdNYQW3GSEplnnhKt3hnGpG
l/Qzb4ibq079kWL3Lx8mu1iSBO6RblKsgeTsbwP5ucI9Ce3P79DTh+UMsvEaCB7//7rtRKPg2WPU
Nth2slPzitmk9UpZ6Dg/5cQ3jVmjm1aXQ8d/KNNnFVippFrRH+oWbOZUkKaPQeeOqZMpWCZFnJIN
R+7Rn2OTOdLaJB/N+2Ysz6mTretzsrYTqGUKirlzaeSradVQx9jIxWzkS7LW84wgy98W3syD3edv
LYh5Dl/tPlR7CCeCm3TFq8bcWMzWcXLRWyTiohkEYOwfRXXr+9JnYnxQ7QNt2f3iMnIdjbhv+TYm
8F3PZaTdtnHXDfoMnuKFOAKWPBR9Tqss8LRkYrudNUyoSTEXz9yYw37QoTUDwAUcfB3/9M2kAw6c
a/C2cCI7y29TllkhKWBaoE4ECWalaYe8/rfWHKZGmHg9b9kHK40nmfQyfJkIG39TEP7D83C1a4A1
XhCIEygQhNyzxBkLjymjUBhmTTq5vbhVh8oSW+Q8eHKfKE+BmyuRdtPGx0tftkmVfvdOWpa+TSv7
dmomvB1JLNy0v0M/YsWnk1a0Of47F4lS5v0R3aRoce3p7QUL1wWH8Jp+CkQBGBBwYzKwz+b24q7W
xugSibXdG9+zDy7gPtBRiqNuTOAvV9KMZuzA3UblVVWQ6jNG1opq8VVTFPNTkfKir3i1uNqnEMF4
qMtOrhfNlsc+u93kjC+n5g653sSqjBWLtbiY51ODBlTb48AHSUiGbq+hWyZtbjBIiD0d4RsqkTqs
8EkrTd479NnkjglW3bdhEiP7RjbsaFi3/q+AQQBFjvTTrpTKLeE1if9mfO7Ac3bNIezu/ZukjFro
wSCqCnrQrG7p/M+dWy+J5D5IAkXA29M9etfHk/qGE3t4EkArH4zNsciI5UzrtZXuDr1HdRDLT0LS
ehEu5Y/hePNfSg84xKJCTZi6LzqD2PhCGXLtzsijRA9IvgwraMdtTCZ72/P3SSX12OSpmpoSQFRm
2SqR4h4rL7pxOowyFiICc1nydVUDi4Jx7jIyYnWVjzkXp47JMDKv2IRB1SZjHSsWTt7Plx5l4rUv
Uy08ievdjuPdH0bCxn4OKz8MVPCv8nLFbH4KnWP5MbwC0jVu+/STIf+RWMv92xhT1fz/OR6bHqGL
8Zxe7jQOqAQDivpwaNWbfVkmR5/5awaFPIIJb7bSgl/F58Myt7PvFAiRscS+rjIto0RtndMKfWjB
oZ1ovPyuk/UFxwx76cBJUWYIMj1UApNIkbSzi5jyHJMzWRXVEvn/C/zV1I+odVAqE0L/i9Ru1Inu
E8sjvphKeH4faWIG6EEtFixKm+0FHFj5Y3hQ/SiFMmzygKfZmYoMKOzpqLs7bT171MsPGr0ABqKo
b9XJMT1AdS9KPNIS0HGi9rgL05LgpHgcT2j55RGVcuvs9luANOl66nxW42JlDO7Ye8Y9r4KGD9xx
0AT/pKzQ+SeTACZ7uHmky/Cf1w5Er8d0NWIye96dMEu+Q880lTqb7M9Iq20XGt+4xEaD/JFukA4r
yCb4ya9hRYCsSJ+s8nGQOYbiNFnorGnvwFFdO0sOncIyQwVVouJhQTyo3XeHjWKdJG+jtB2pfDgw
MP4klGz7IhHNtMnqBzCjtrJBQyl/xjaEOHPVUNi5xzH+6aGW19mqfWEwM99hONAUdx8jQlSNR+Gu
PHlzjJtTyzJ0HmGFE2Z5oPTuvMA2ndwvHLbDMX7sfAkF14p1o6KYeNYMKaEdfsJVbkf3KdfVtudh
uuN4Oga9M3z0AfkaGhKEpSc7adP1ZxbvS31qH0JW/DjM/UoId+57RilQHAzZFACamePCHLYyPl4K
xcXIpGiJvqAPFDsCXO8c3eZ11rIVwCO6VdR0Htxlj0qtBWvu5ECMRUso42JypYjJUvh+ozQDGZxK
epb9hZtwypzc2AOgo+MOvMLx8I6i8Ql2khChkL+Fwut5C6vKPvkdBu8QLPLzvB5r7FFU/Ca76jn/
iSzH3QN4XUebJqHefH07F4+KDwyY57mmSeljd0nKyqEXTRpcIvem/syg6QKfvWZWX69wBUtdtFPX
mX4ei3f/VL2SGLQYX62vnH8MDpOgw6LhtnjrgW20KjY15f+kL5BRP5+hYklkW8aZmrCFClM2lnto
G4AQOIc/TkGGZobTn9Cm8FEMEOaQydz1ZkOMMCCqsNnbUVHhCGQfBugiPwa1HY0pLr7ZRPY6ncHp
OE5AVPP90zQr92oQz8KfpoWk6D4kUcs8f43MWc1MYRCaQcIWlM9HDllqHhHSf2EpneXkm+51vzzz
RYWT4gYpJGq8mMrXQvbB+cehjmWDS/3fCtjmMgdQesDjya+BDhvbUcWMJqffmb6w6sQfGnCt07PF
VYqyvW3yJ2ju7+EK3N0t1S8QtvzEksO39h2KS8jzl+GvNPBGL1yxWOU+VygtVkAEJeCgTRyYTJNm
rmZqYkxkaLnUtvDR+d/1+hrWiSGeYth2uhlLOU8jVfJMhT0O9jWzt3ewQdP0VQVEmtP6zRQjimd+
5YhMf3g9oM9zcmCAQMt02RO4/uVp66mOzCPudzByCeMoFmLrHVDp8XDR/Vl0a5Vg+5/mdlMdSAiQ
QwmQbveQXdcKCMCNjJ4ese00P9OzfhRz6m/vG2mnuCJ+h1X9RUWc/SxMH7C0q/mKMUtZL/0c7UnE
eyrF2fpXpCtc729e90vmzKfxvLJVP8CQapRfoaYZAtdHYmqGEkSH2cWOfZ4yTMwjl6VGTqnqcwZB
MpKBKDU4tjjaMDKYogyEemI++wQEjdTphqfVrkbr/XWuzZv39CbBQd/VIKVtTZlCylgoMbZ3fAhD
g3TlRrw6nDDRdrNCkNHp4bGudpccwDYkgd5ZwgJ1cYGXjvBh2vDfolAJk5m/SWc9+tpJoR8RfP3N
ErN9NmlUNbfo8rSQo6iZy4AII0W+n7jD1TOk1nuLR+BznL4OtaJ/zGiATIIolcCQJ/yhbrv8kguC
yKGdRbd544aaQJdslVXvWxPbaLEwMW3i0ipqIOhAmj9Xy5zELzdpVrGbcx7lwprhddZiTFIrCvEf
vOEzAFf4OCWC1WZLuw/+a9tIXu3Ujm0kDt2R07/0qsNnDBpU89aKEslOZNa+Wn2UiG6RZVw4CX2O
w+uAV2nHTHAC6anC9YgEqieladQl/bJfiPz65XbgXl+1cJ8kX6nXG3iY+6gsVpl6ky/gn3Gr1jBX
JtqCWeH7PhwmINj6TUopx6+eV0w1cqf58VyzvM7nyqyeXA1ziPlR24ERWQcDpUyFZeZmlf1Yp1J8
ZkICUB4UIGfi6gKCbI1PgUPq8F4Vn1fk4gqwowYeZXKerDO0DiwWcHr0wjmCD9g3hvT5CAuom8ZG
9RMfxxpzftFiIJeh4G3PTORhudLADeotEyt0IQUcDjLQpsM7dNBBM6cvz+PXVyOqCWoavlXig4IU
2ipyL3AA4ToXSy/kioECKlI54pH4CisPmcS4sZSY1OtB5B7co0H709/wVeUy0jlXfKNfy2iNTe3M
o4i+DFvQBDTZjr0vNSi1YKayK2cEUVm1WFywixG0R9AgvB7xYepJaScdxsNa8eRiD35hkfylig56
SV++nlddNAcfs4YNxtVevPWUiIKkK8zt6682caTqdM7E4Ot0j+670c4NJi2Gk8roENhDWhII+gLq
HNHTFj/fFfJDUgCx7+FngPPeWJP5wIFMFK0dMON3x4zUreZkW+cB70ijVUQdaNgK5AXZvuBPkAL+
4FnD/hMcuynkEejJDc+YLgXUJKSc68jaS7qgAPJcajBkZNKQILXzunbO/MNu7Hf09LhtEVrWzQJc
s96dDppFaMapWJSpdZ8w8OFVa52mLKwity6qNdicoQV7QkTWy1LaVL1AGORRTgi/+fn4u9y9OlxA
36wzi9pIHaxocwYtLgMmGdVkjSSd/iMIFz8tP0+10LxnZhMcLPqFSoEzIwG1Pv2pX1wcriic6Ohm
GqiDFabJAe0bpE0bgTuXrEic+J40urGzPkfUl9m+VzFpSBLf30I1K6GjnkmQdo3viVzDQbQBGjGy
45olYdKkhDIl3HGE/L6wDDXK8+ZJB/K/+yJaB2qYPmI7cMA/knBlS9HaOImi7GMyfu/2GI27Tvo3
jA0yGgzExTAy2m8e18WKYtchgaS8fbvMtagEYHi3z04twIbATz2gbocg7aNR8d1NJWU5ZOWBHs8I
IkGWMoIw7ky/v7Poe1lXUlrOHQHJQCkxB3BPAFxAPRDCu7AkR6t6L7V6CmcI5ksVR8U+avgp6CBs
1GdA0KNxaaujeUJVxQZ+fUzUeurgSQdvDPCpLuon7GHB9zKwEjxTR00u6rbD09OS5BYkFliTy2Ho
PoHWXeMExuV0Kh0fBr5V3M3FmjGpaL//2OnbU8ELTQOnuTwvM6GvncJecyRiQig/Jh/+NaF5z6Nn
OCN18YTLUi7t8WKLvgFbN0svutZOwO/nNDur9Z3mLKtarhrmRPiiccePojH0gQD1+AKJNS5WQIpl
G2UPBG9ze4t1nLnpSXo11tp8a2rOUu9kAfVHMC6XhWk2v09DZbPvtgahsbE6408w/nW3dd99FeU/
pX1BLSWr6XdoK7Tt79P3SjeJrC/ScCk3baggSPWhtPNbQ3i1As6V3H9MDaoALyYICKU/ZSCGcw4X
BAlsRkKtVWq5of46wMU8weNbjJh/KKseLu3UYA0vkxWU6EaXda+hvyf5xshPhzdD9c/hYo5Z4kgQ
zd9j3dkQD18sUkl2RUrgus7Jpj0YhfVOuwLonV8tlezwp7rhn9qYkIemyRji1MHjnUrLQ2wISlN1
Rx4hGuPV/Yqe/oxcAqh92yv8Z/y1KS4IFsh631286IO0f1g+ge95mAeeBuff29gwwjzQEiFWjAkl
u5VcX+I0BjXkowWAcfZftSCm92qCIG+r26wNMnQAKE1/0bMgdO3DFBq5k8Ir0IykEqz0AL5OH6EP
QDS0UtCiUHghxpf7XUD1+zDEmPK0NgC2GKHgibyYXTuKAR628duo27eUaD8upJKS9H8vPOjseDxf
uTlCb8OGS2xXTuYemUKi0t/SzbJ9Plv0BGOO0eDt6mf/8/s/ZmvPhD5GgAdSxAUVGn0wD+uHF1SG
BT9mgbzJ2rQ5jeDVQFln2QD/lg+YI6JhBrpHZftbPxkZDQnsuX6wQI7LNDqb3hlc+ZZc1Q/L0PSM
/w8Fy0aV3fDKKGllVXa5MiSJeEj+0zDKZNg1JyHdGBjhI2WV4riPyH/zsEsQm7UW8uVt0AbidHNV
scAy7Nyv4TacpZmVqb88HyABpCwSqKtb+lpNB+jdmOK9qTsH+etkpodaUYyGr2PsAQigZLlZXklo
t/VljFiD8GEOG+CDJ/9oQib3PEz/P5O2ABHAegf0Dg8Bo9TBAcYms2zXpjgGERDgHy1dzunDdnXM
97ufqr7rjqVcEmQIC8rWl6CGjUgG3Owp9GbyCeRdbkVYgpnnGyzE67S7Q56YR3bf/wuARrXUg3wx
brsNs297dXfk9fFY38Eu+fF7JrZ5cqqlwd9khQrjWDH2pz/E1MlOo091GJtyhAky9I7wKPqXeq2G
p84toVzs00Y4hZoHSL9r0fCm2VbVU3UpRzT2L4mPX+TZ5VyUNSK/MBgS4fmvu3FLjh2bRJ6TztMJ
aS6fjUsgUpnqVUFsOm4b6j6ucXk5gZesutd2eUXpXwaLKkCby4MCl749F/IKHEf+gMpj2+e3lSsD
GYtm5fEnFksim9BR1yrZlnMv69tohEChPtcEB1RTqENesE9yAO8JGg3+a2q0WbluAULobFkZYfod
BsV7NcMJqMsDgj6ukq9/o8MkxVijGgX43UwwGJys65qfuotg7B0BY2OClpkWd4rz0Ve+dMBGZJ2T
h+Uniz/ZYfzJ6Pe7VdYsSGf6pq5mjAgVqErsjJ+bZiTmk4bI2px/tKnTz89FRAeK2zNdnZ/EUpDD
Vq+8a7hJtg6LHHsnKzjcd4y2FGS+ZHYkFEmNVsJG4OBhmiTDEXEje69PEpSzq0VIN1Q09OTfoVxV
sqRUVSCtrokVh5viPpnzEev/8gOiI5eH+GR5Kq6i16p1NtASovd5QFImswEFHUuNBqkwRiWE+fLM
FY94nigfckO7g7W76yIYzpkqJWPaVW1y2uLAe0BTcGuah3G/mEvdTJaYVr2wSixTjG6+Vwd+6uaG
ZV1A4YT0JZ05dzsgxh7ojWsxurbvCLv2clOhbO71NWxX2jglJFFTGGyd7a9TW9kc14o19SkPpMR+
g8R/eZKG0YnZLSGdpJ5iEhxbpljbcKIc98T6r08B9tNW9Oc3igg7GKPflyPlMJrk2WiJuQMGcn2J
C4FYT6G4qfCCU/VIRfrclFw7DxXoSlNVEe5iiQIhlasz1nweoAlPUSEXOjen8LyUZzN0VZ6YkxoU
fbdcWF8AcK1Nvuvynbu9UKzVFKHscQFY39WcMUxSIJHwC6YIIkV1cWyHbtdtaRxVp/e3oqQOUxCg
Npslojwz8HdTKv5JF8OObo+vI3BjCxfWctSzUle9F21TZUk8PCPtxGrIRXjW/c8iK54MY+4vXvmC
BQL7lKxp6YzYOzLrLqpu0qaOhC0p8dr5e3h4TCExBRyx3c2LwYlIZUFKkck9fj80SER3IqsZ86kg
fA9lREN1j5dXKgo2d2LVUExA2hajbbnngST2ysh9QWJARdgT1dNJLPvPso0NLlc4ndd6Tyx2r6Yq
lxy0JZB53nLeGpCfKAkE8nz9P+b69vm5603Nsr5nPRV9JMmMPCNJqnn3oFIFZmHenjeRjazdrRqp
e5czNvmcaCbD8MzsXeuM0fKJDpTTc2X9rU5z6negqi19k8pMuhGTI50+ZV0SZ+DhYvzWfJN4lCuw
upAA1/YVEueF/tcvS+8rwyX2dyPuhIshsgGnyrEr6rjQsmRMemiuYJF3OKf96krvTpwGs0vs7Oko
bkcb/OpVCyuL9w4rMRdTa+0wf+rHoa6FNENX4Wk7GO3LU0phASTDw1URElfHYtsD1QMfxIz8uB8k
tq575xuCf6v08UJXF2DEEdygj8HKU23xaHuI/AfGQVkV0Aor56Xuv0uSDnqqzxDd43KpVnhmEuaS
FGOGU/oNmPV8bGMlg8EB2q8FKLo0MuwqTNxC/METBHxcY5KKVuTQVdqZujomsed27jM/d7lka6Z2
+/ZhqL684AV2s+2qVEuxS5Yf+Ue17ORmcX6scoKpCdTsgzxLhTcn6CG5hVvTH9hSZEyVyT/GKuv1
Mcr+nIHcMAC21ct/imLCa8J1vYCq+CIzI0ZVAmJYhAbus2vysa9yUEhcQOGuC8z1g4/4SGTQjvW7
eB85O2n8Pd069sRtS1nV1B0wvdUZTfASCKcW4obbsSeAofkzmKtgWj7cYwbddwXGxG2zhf3BpoKJ
/M+c1/aJITSc7GsBWe/IWhXazLtzCDexSMFq8hGOAPUTGyB2Ua2w4H8DGKqX3TRxxCNRjsrDcVdb
Jouyuen6NF1HIxax//VPSi7zc5UlwbSYI9jl2G8N2pHDZdcTeBwtReO+oa96kXo7qTDuSAwl6+Pj
SewTGk6U5MQ/0VTRwq/tJ8lrY4GzsjSEytB4U1fd/v5EsypzlGJ7IXc/tdH7JY60RRzWZVAB9moj
4r2zBSdWSuvlghikNn8kP2t+YKJXChUvLQ/JpGK/lv1cXvnu8CgT2ktFtZbsLR7JGeN43Fk8Lw+o
RCsplQ3gHCeY/5RrtrAFjAunoJs0vilNVw1qCtny5ufS5VBAVBWNE4e1FZ5dGZubYlnPDIBjTBgK
26jWdTPCZxpUve1mpgFAFa8xc5T/Mf+A7236TvbtLOt3yDO2YXihi3tuag0lBPifoyTJp9WgAetF
jfwEyC4K4TDjqzDLh2eosGNsTpi8Rlf1GRJhXI79/rpmL+P9RNdhmSWKF4qZ+Ao6iqtQFvI1wEP5
kUk5LTZFVYOMIx0tGQmLVJvOdZUcvkC+qHQsMle6kZJU5NZrw8ufIwJ/Nc1S56W34HMPe70rTcME
HGwqvBgOf4TwOlqiqnIKrdpNHgrzNU743i9l76p14ig35+GCA0GZrhqs/qLjKp3PqD3+GeOnzcWP
++jLJ5LXcCT0vXXzicHSzQMsclmfGtGFIBxzEJQ6sGjLA2NnztNFuPcSEz13E+qVs9rxSon4rC0e
cdyl4Znys4hQWOBhhK+OteaSbf+MY8hVEMcq1XZgj0NkZHp3neh1HbSBj2y3h7yYGP25uZi60ymR
wtLcziqchsMUUW4UA6pkDhT3Qsa21mbZx8qWq8/y+jBs72Y6Rk8XL6fVC1qc/iEvb15xSETVO+1T
DAQebpNtcksY4ndOdAV+MQ65yOPoATuEH1DpVNhOResLonlOf0Vxsr47WtrYNgApmlPimKV7Rxot
Wv+Utbfu+LO6BPmxZStafeDAS4z5uNrSQPFccdi1xYiLoGmeqzjHwPn4fr4FoUwfdldbJyJqwJiP
2oPvxx1maRjWq6B45oQZSsIo26XJgK424M5LA9fkCsnqsDqH1MqTh9BJ/kAwqZubZbXyty0dCkL1
e86ULyjlgtnPkNXPqeYdqWmxb5Y/XNIgQzK7QC3l2qRI+zSmLplZpyMwgdsIjdwvNn4Nq68MSm5S
hF4uujnPK4pF4awzRh+2WtZF0OU7zN7MFhOJeniZ/ouxeBHbQik/CmEXv4K48S2Xao6Qsv91Clm1
MvnN86giF7WPKdiCCJaQpiUG+sYFl7FPzsmfFRDa/GxIwnJhl7pUZQcXfSwemgYIyzYmgacioaB0
zF3LD+aNuqToVKf7WDMn0o9W3uK+7kXNJ+R61IWGLbvbFTLpOJXvmxYgvnnGnpAGIrRGH4s4cQlT
ihG6NFbgTNyh4pPhAy37aBy2OgwEFz8aSLZtrGIaRfBxcZ1LTpziuHL1s6+serg43GaK/XvxxLBm
TlQPKPE0mk1S8ogZOp57eRZR+z00NEqbtLG5dtSGJOUVy1spCVeOYnuz4JIPZNFqxCPS9K0Aj0R8
ox732z1IeSI/5UjN/DrWonrO8zQhQelFpiLB9mzvsBGqB1DQiA+i2D0anQOzWit5cvRnqzhCbNEQ
UXp1GniuSAE5XCHhhcZAJoV7w+1dWsFbZnd7lpHCz/D5ypTFPX35t3BSUditf++JgnzDwu72lgPV
mquax60kfsKyVvLMIfm5A3xpejKFJo4D3JRck3VCEGGHIc17NmxJSXA4hq7+r9ITsIzPtnAbUdmv
i8rmNVrkZnT501XueXAepwjGFwKNI2jcyTXUiOmizm56otX8aL7lPj693QMelZSEBTnYEbMxUQAf
43mwrBoZTLq40H8JWZWoOQSz6eYo/OUNAGLZBM9y4JZWcTH/yRDdlPI/97tCzHJhmOp4CGOQ8wzm
pqOtkbS2Ts0gUuuVsR/zKf5BwoAQldSmO/mPbNRxPZK45RWpb8zLUM2V/dW20drFCz3frVZtKA7m
sth5arDJ6kCANdzv2sLHpM//eecGCAvbv4GPm286DHiCt4JxjGO0wOpWNqtnONCTcSXgwvc0ZPB/
vfJm+sxicyc6AgfV9VZf/g2SfjJc5HfM6/H+PpJfxvvbZbWy1SyLf++DvlZ5ByzZaER35UNJalmO
ATrQSfPo2Jf8ZEElACyYsmVjdfrh7kFvya2BOqE9z5MEB5/THyrBEw/qBztP2F6+AnL1Nzl+mZZB
fNOK4YHBW0CsSM3/VWkFqPF8qVBAwzzeny/88iaReFZqZ9Fs7XUk0RFQUJAckHWWYlQf23ewiRjC
HEqb3p+yM7s0NGPnsCgSVSopl/RWnmdOxy/VXq6jeh7tWMsSAiSNFhQoqIDMnz0zw0uZoqFPDxmB
SkluPO0cyelNiHaCg1iBvIc2hphpn8yVCUNhnamwH3YiOhcrrmv9iPN35NhY0miG1/enCSivb11O
jwfC83gynKsUxEBjlHS6kEyvUHmXs2H38kD6UK7Ici8CdoOtptvW+iSM5a5tqUFzGcEX3GUdQMTd
p1oCGQps3RLtASHOjIt6opp0Y1OcvwJkZRd4k495OUSz6JwVfD5s0dLi3LzPo5L8jQLxS9NTbRXf
FPU9DQ/C33Y7R8XTGCpLtkUwih+fQtPfwp01bwSqG5CaN2UpLvB8/3rfp4q0agj5c4oEnZ4KXJHC
ksYZ6u8h7Xobkze8a4hJaJz/RJfgbsgX+8L8o5Kb8rEsW6CpXNRXjHJxYnyhlVQSukKF592UVdjW
KPFN/PqptyTo8A7rjIAj7r/nsKzUJ7t9W5YCaAbnKDr4EbWnCZgples3z3kC+iMQp1teTQrwyn9K
Aq3PVmmyEvTQ6bys/jk7CWo/LzH86NJxJG7GCSXDB5m/vkkTgKx1wSvQXCMwV+JnGP5v9lsoGCi+
yvDWSjIEi4cKb9TK/so8D6O9Y64nVxqp4k3XBwFA4k3ifhXcEloh07fcFWcKjPE811BnCqvqnZ6e
6REfBScN++vJTx90urPsEoNJYNa8YOxwudgTDvdbW/5ViC0X+qgsqyKhmNWaK9s82VXcRNJrdA2m
dohu9cmPO55BzRCeF56tKl7fpZovEb/o8cGevMddKGeuqhlSYjvtob9onGf405TywweU9SMU2Wcj
CR7ptdsFysOhM0W5sYGeL9cthEmauXuEphtuBpaBFKvYKiQjEDuBMddFCM7DtuJWZrxXKt1vAsNS
mRfXyz+l76vVBaU4C9Th27UWktv4pFbtFlk+6QvzR+TnVo7dKS6Rz3z3wuzUrNVsu9f8Btalf0o+
kMbGqVmFvrzhGg557xxnmyO3wx5k3B3h2vYjmlCI6NOHX8KTmwfe8ZmVxii2iHgncHMz4lhkhjxD
EWjozLPLOw02hjc45wASdAV4HZfzPbW4bb3s8kx+bvL5t8qR4iOfYQuTV70N80fDnVTYEMd34NFF
zn3xfGa2Q/sFgPWphYhcBuzYRrkorNG484+OOQ0Zq1dWvyMypEdH6BGRGZHMpRNI5Z6D3ZZp0oBV
/p7+jBFn9E4IK9oB0RMV/4YiY2hcy6AwJvxnrPa+IOAjqWETckua04EGEaBekLw+SYyGK5q/oEza
zU72xSOQb1KcfFQ3v7wlnS/+yALcKNrEnokJTgflGel83kbXl7JBUPJ2H+HN0wpJr4lmD4LJra+G
WSlAIlG5nosYv8L8JGvOzAwEvFeUPSiw42EEb5Xd9UlQVbJVfqS6CUlvxzV6x68Ft9cbn0HqJqK1
IdlFhAotl9WMov/u4IkjzEm7u6WMMXRG/hD/klO7ZSLSytc126mf+59XIHRDHKGhUQnvnnYU81m9
zqUOk2rXxlZJZm64reaWs2tSlsSM9zhRBmlTwlH4iayb71/yjJBCTB/z+Bycp86WI/dNrmIm3nwF
YRPWnCXxIXaxyKcJtTBAXi7+jse5ZyVgNJthF4ZZx6HpjkFoaYaLWi0FFah/28i1raB30V7iZyku
76hdV+8X0BUH5ZMJJ8elbKXRH6KEhVAuGViibolo7Fq8FeFPI9y4RAOUC/cVfNzX8u+gbtZpO0YO
v5665+nxjbRJnaMcBPoHlu+QBbiMm17vQvChio1gxuUrrpPrHbgUnt6vZG6njS6xnjlGTsQTfd4f
N93fHRQOZWdZNlE7gb+tS/qp9zwZRiMoSjFkS2VPF3fXawjrUSDi7bPrwAU258Jms+iIivG4FKKp
804z48vWHc/xo6PDC64w6LqF5C1dAs25AH3MB1X49iMTTuxoFZLVoLeYjUuuVxtgHvPhn3IT63eD
DSnHnIxiOTZ7LXmfg5x/joXX+QTciqgjiJO2AQ2ZosjmeT7KNhdddFDsqjSKs7DPOtaV769gDm68
egCTrhqKHhuQrld0Yd0YpAAFnvcPo5Q9g/9OR94KJM5hI336NyVgTIaLXcpSr+ZGK9p4sDi/cxTf
3fCpde81kFPdu1c48G8gYkFOYv+SpXkEruFLl0tHPMBlWdSLCcw6i0KL6yLBlv4osptNr88JIh/7
E++UQetMkSsAj/ofxZjOuLHsN2noiEa0ToYH0hu2G2u0WdnCQ/OTgR1MbnUV8IqalPZpuzJODckx
NZ/PBC2Dek2qq6idZ6PrXmRpsFdrQB3YnLdusNBykLuZENCSM7iRwClduGhZmP1Uj5y5ra9SxEKQ
7KiiEhCvyC7MdElUgvjmFNckvm1OxMZ+28o+pLQiGmjnR6XWLVJuw96Qs9DMqVPz25fJJRtda1Yq
NG9K5OpUxCdy87G4EsdU6cgQUV9Q5kF7QzQ2qTgPnsFdtgZq9KGw8Ulz9fYOkBOeJ7zP00OLBYrS
q8hWkOy8+Hw+enCYf9O9yViWKDApwOZYqrPjx3wm9hsOiqFRqdM4a/FKuiNEeeKtY5tolF5Y5MoV
DKsPWWA3gp+zp3QS9ST0yixqIj/eRX5nfOskRdYF+14tvlFr2HOfPm1vr8ka7mpIxSp7/paxELhK
7uZRxie1+JTE2thp8TulSQcYipG2+42avHvCpPx0Sjiun9omi6w4KLbGqEnQbsaYW1P0LxwfYCsf
w9LeeEOSroIQSXCDw2T2grlxFUXrIxH1LOP5tUQXguFPrD+328QUpoRaOcLEQez7efDbkZIZugrr
iWgpXYI+bgivGRkzahljRjfuNFCwQz31kzawAsXKLJTsjIGSv5/BTDDWo0UqsdC684fL2zV83MPw
xamlp28DEIBNQzaW2/yJFGvaEUOWpDE2GLF5ALQlBDpOUqJ8d4Fi2cPFTMLM0hryxFMsgytf2qA1
og2js0H6gMz/3Dgg9CLkSxpaVb15jzB65aQ+x6w8AKLfAWh+TjPuQddM0IExIgIHAfjx0cTK82AO
nt+ZIecA2ijyqXtWJ3LzvVOctu9v7cqQnz4u0qTaEl7Xe2rDtO0GC6j5Qshd9PnhoTRj5y70h17U
cr0aDJZfvhhoqLwsnKa5icl0o0z9xOjL7lDSdy+d14v6MKvORY4ucuOnSRl/+VbDATuOh9ZI4YyP
1JodZUArynVkwzIfwqs7M5ttGHeW4yAPqdiwxugeWc1oPCZrPjH0SsmHzwtbNcfmobjbf9OemkCg
uMJsqTgbA3wGymvB/5HJP25csGfkqj6uMSNFynV9xy18sr9vf60/p1v/+glH7mgqyXLJ9bPpYFbJ
9D8UNdNYZ3CIEk+Uqx0ZjUEbuVvRPcmzUCl0sUyRkzVpNVvYEe2jeI5fM0lIjdR5mVwO9HTUYFRj
0mroCKmK4Pl+jIyWojGw/Bh+DZY8l/9pNhPdVZSa7GnvOurNXPnPLLDFcaZ8UmhSd0AO+Sv0TVEl
FWZ8pOy6lsEW43AoeBoM8u8XL7aHHrAt4Dd4dmKcSiitYFGmmISX3jaFdbPiDmDTePCXQEGKSLa5
6ewBA0YFr9gLCBbwf1wiGZoQZp1fqvdHekYJTQRzxiGOrMRdCpns8wafVDPD5Rp3BvFIoQDA8Pbt
d33raKu54YrQPblFRfXWp0MIRDm24Cy2nqTAursN94+OYikqGnQ+PBR43MZMhXjxnSyqdHZFFXkd
ZdVVJfIqbQxIBdrUNPVydinN79oNTquCzs6rVhbs6qoqJJ5W0VwYdWesTdkJIgl25rEHD/lwVDjF
K/IGS6+cmiemUZeyuN1PVK+u0mdWGx7w4Xzd534NpKYGtp3SQtcNClgNCGMjJVHhswgQ2NEpwR+S
9vaQdT8FELZ0kal05K1I5SWmi7bjd55JMcKcCl7rObhaXfFhIRpTGR2gSmSm3tlbhtAzkWNq0j7E
RLyaZK4Endz73drrZQnvJrs/YETShZrFssIrmxapS8EMJYatE3oC2FvzdOJIXK2lLD71f78BWSo6
tGh1LHeu9cHfYW6sK0dWsf075/Ta3GUqU9RhJnxYa9gSkhVoLK3QjxJbgBU4MiHpPE4bcLv3Hy86
0miV5WEDlLZ8rWmKDnxHwH9hYKVX4WxQNwyKmXI9rc0ARZM9qulo7lj5lVPcS/JX5oKWkrbt2Dfe
9KsFQNatqeTR7VORSEVm9WqvlTp5tm9E1/Gy0+rap5ML7P2rIVjifVxdBuKfG9LbTIYwiVSO76e0
RKVj6YpMucaE5R7WEKdstWiWYSNamG91nH4BymL+z11PEaMNZvNxsQAgp34yjIDQiFLJlrErhtEr
AcDeTlyVg1gjxrNh6YdKDZOuxk9Gg649G3itNYcdAoK4HbR9+NfHf7w7c9tIDVrE4ypyadUlHNNw
/SsgEjEK1OwNKZm7NqBQZaQS6bwNYrzPABgNMXWkMGyLd8vs5CbJdxQ3sqESGV62yJJxZSXKJmwL
rrYI+DbQy6krcljSZUYFKsCO2MPfk2pVdFY4lzxQrSw00uA8dEZMTi3j1a9E4c8nCDt5xCWZ7uH1
5ygJDjMqfadscbf9AyYPldgs2lLVSMr8sdhgEoq9NXVDR+H25tCDEte0+5wKx1AWxV7uy3ihrthE
kFakfg8ArNqtvM6ajRr6d5uriFKROoxmsncOBFfhmtPLAVkeR9rF0qxAE9RRWjLvBU57IPS+hGvr
D2Hmj/GmLWUXkkjFntvPQHamgY/8/xiyVmanxZYsoD7ckviLCcVBVUZeZQCyKxvKdJtEtYo1vABB
JZuGL5BEQ1QUTRAweMhctQp7dGSv7HcAsdXlExa6vAox0aTNWapN78r/1rv7Mm2otBb4iiZO9TDg
vSDD3IhTZnu1IJzF1eX/zLvqgrFbugWB+M0VMa3/Npnh3hoVklQfaUXJ7wYJ17FunSriUmHhumz3
uBZEyYB7b0eHFxTcedM4KzEZbJbFFOzUXjENwIrl9+7iYDeDsmJFnPaslabx+OmKp1xbrXP3YGqt
yEKG3tt+wjK9J4XoGSeag7sx/EbEaCi15eApbYaHnuF6jbnAXK0y2mwDncUBQ37z+G7jHhlEBi1L
mokNJ7QCbclbyJsmvrmkv1oymGW68YE1feDHwRx6497toHkkWzp7OFF+qtSADGVASN3JPJf3GLlr
Wi47H1+NXBiFePtMMTyr5A0Xe02CF669MZ+0SQ5Uwc1RlYUXkzqxUzM3wfpYquQ2Foj90YE7foAX
vq3f/I7l1jcpp4UD8bnrFG8H0lmzMSRoy6irphdLCcWwgvAReBXgb+tu+4IfauTxLmJavbzwhJDV
22kpcN1hEIX2xrPzauqst959nnpEacE1M1eXszc/eNgg62PG8ir0F/YzJRAQ1iDddlJJGWdLpFW/
z+LKhBeuhY+NqO+L2VasKLDRbq5xepMwONEx6OHQXfgDh9ZabPklmGEnd67QnIgOdtwzRCAhOyhx
LSbLLLSFBPODc3Cq+By/afFLWcO/KrDgIJOZK+6wr7bnNE74fYhKBK33TsSlqPI4uyHI4UGSMmto
+dhV8JoCFIq/uqsGrvfvynOoAUcjljtjDVWCSmj5Axi4+Jz78QaLY87PTTQOKqBJY0jgmK2Ylyuw
ogW3ILOihgfl8yHN6ZAyMrbFGJxgxNLbfsQvuef9MrQrUIeKWVJdz38PfUZGiUYwmBQGh3lyy+4R
7EOrr6tt/z7eRFD8AnFrEck+K4zUD0aSIEn2tJX+rZ3PgZ2/1pBwy2B+e/T6hFlsCw8jO6MMSFLx
dXlHOpA6EnEZsGidedY/m2+n4uQdIpRAVNPC6Aj9mppNt1zZAn8IHH3YfjbOtS35E81L4tP2Awpb
BS5UfnHC671OPbDPBqanICAo0Ka3nktPiwHqokgJnsUEAhXMR8EF5ObUMEAe9WpIrnUGT3LOSWFr
h74AK19bT4jirFZSzIRZ7zpdFvnt/3dNOZEGbUfiVOcpFkIJZe/HaKgCgiVoCLn4GO4J2bBgu7ez
v6PVuHVBDJ30hGeN9u5syeW9eSWN43wxLLi0HeaZkct/JktWcFdGqpED/siIEGn+q2GYtdtwItUb
cSXJxEt5hHuv2kTmHxqPCekftyUBEc5lZgLVAbH2nOC2rTRiBFGy+vr8Jzd0AXwM4szvNNUMHJvm
Bpoo9gBPag6Hr34/bLl3yni9xyaH5OIiRhzuVzp/3csRqtm3LZMKfdz2RUxA2L/ScxI6ZPTlSgFZ
lVTh2wLWnK5N/ihM85+Hr4CdDdumMOsDcwmzk0V8SwS3BPpryNfuDDy14xHsb5CdisEKUUzh5JMH
K2dRic3Crf66S7gjmSFXDGDvsGu+HXKrzZjndXS2ntbwFFFluCByJllOsK9YfRWwD3LRsURK6dcn
A85yXgVZdPtYc8GIavAt/USrf28/UnxLdjFwY96o98qcnrKF7oWGROqff1NWtAPt1iA3Temu9FVM
Hn5vqb5F0s0vhzms6l3qg1UYz5ih0VKaHT45KA0o6yU+GBpyAzahpwNjxjX9MVMMbN5dR59nYSVt
malbUq3hvv+Xauu5xffgwJoQcYIMs+Cj3hn9jHj8y9I/p7Tny7d+PSz69G+X8iSjIxv4MV1xPisO
OQHt/hQgJNwJWgdydO2XlW72NxRGzzJDbQ4W0cFHNOpOBP0YoK2PVDHQYZmCPxQwKVmg5GWJ8xd1
hmoGqsSwI5RzKGHYGAFUdHDG9jeZYqK4+FRUWEny+EXzDFcIoCeT1Nhn3TJHMp3xMoVLU83+mDpC
6Fpr0YWp0HDKwkSVgrKa/tJtzNFU5PxeCX80wVg59PxUGDko2HFU/sIPLNYnfSJChUauPXPNAoS2
GhdJPOX8hE1eHOunzaz4GxYuMJYKDC+rpGENhP0wNzm3Ri2Wsu3GxeXVozifOnDjENeZST2d44IS
2IydA6JiNuJpePB3ZwyR2OL6SCYQoRkIkM7VoiITArck0MNFXuiIJppSb9ZQLnJEXc93UBUc2jtm
1jJqyNWe2UV6fIC2xmRAJPLUMQqlV57Jhd6PTdJrErWQVLQb1c046kd/2mOBXHIW+envbee5o+yT
GYHs5UfQ+arHHu67NEj5NjsR8mwBXola6YccEKw4tll6VeDLg4hZ9H9wcjZe3kgKpj69epadQtGJ
7fcb3YaK+Dw38EVsWMlIoPDEKKP4n3G+jhbNlKVQcSIrW1IBRh2zy+MR57EWbT9ccIDHzVV4ce1J
T/bCFC/p87ygAaPzv6YteWCzsaZkZvm5ouktUaNsjVrnXTXiGFAdE+eUh5srnAb31p+eyjraApG5
FCuNF8W5eUlIzlBdyXzeokroInsqTOTlAVzJcKnUcgyTN6+bQIJibaE8LHDHPMr1fOd04nYjpAlU
YaNHEAsy8TXVq9SBKQY2I0dMzQj9guTXFyMsoWdw44wlzemv+I/Is2cSu8nZS6IxRA4+M0toUhI5
KtzLUjGdRAR6mkIyTNu0BITqTIKIP4RG41GdBVZ+mHfnYWpQAzxZBTo1ryv7yeARrf1gZ5qSl+Ma
yJdMiX9EKKDf4vrwQHY1UC46n2vPX1KedtZbmNAy+EzhDLA+YuLh6LWHEWlGHzcbof5jKTgoCwbM
ZWOvCZcKvzhuTjm41a0j/oYZz7szpZ/lBUiZcGFvdyBDKWnmmgKyTpgbESBFFH/6pqEULuOyCUZg
6/fL/b+Ne8gkVM4GiP77z+9+jr7JQrZIqrqTP54bqz8FshuPHDx/sHpecsNHm0M4kD11hlUbDVG1
YCi2cXirS4pme94wjuwa/DNbDLmY076w2n8PI3Ixs0VkuDnFS3BfploZ8S33DFEGrELjz9Xt/syP
NY7Zbu8mr9DFUb3W7x9kHHSYRQbq5z+jlDvRjuIcnMA/wE/6mBTovM2NLDXBbd0TqbUit55uc0oA
evy5WHHvQmK2/fIEVCDskVH7ZxSe5+S8WR1wEbr/cT8gdn3pafQ7zVt/4/zCmgjETmhDYBk0LGZZ
/7f9TY6GDndyNtfXyqjrZjouIkmC+gsTSKVWFB/dd9KKoboAjRHId8Bte4cMuJdyHCiFoHgpRsny
TBbInPV01O9wEsgnlIk2T9cqBwTQ0tNINNDecLHSM5pU/2/LQfgzRjAfiYYRk7nM0kBIM2dDC8ML
o7jxxRPYz4g3ZLumA9FqSb7nQ6Lb7FFmReEOTINmWMC/TpzNN5Ietr0lpa8mBPUU3UjljJmRNJH/
Et0KBiDJvMYN6abqLUk7rHWZGOMn4Cl8h13H/XUCAYKsmhs6SIe19YXoJxazn/pMHDTFb/is1pcq
3PHdcnSmqsd/KdAW/55vYySP9f81lsOLt50RI3j9zHlM9d/s2EqibDGtOC0g6+5vW5UJ2zLodLrH
Rvgk4j8il6FmU1FYejouGnPQzZQBXaAi9aidg/Aixbf/m4y37qew2yf2FSUn5c3XCfiSsZ99+KxS
QcPXRhZdzLpk0O/is2Clj3RtMrGrHUKByIj/KQT32dMdqDX2cvUmCU9PUpJ4zkv8FhSzK2NMO9Aq
UOgSjnO9ilhiKX9IeeMaWhTwWdv3JUzmBOqMNhUysnh3/guIf5T6RF/5VL8WcheCNmJHURnUuPa1
8jMpQYwTdlHw5zPoU/8uR3qstu3+eDcweLON17kwHMLqAtHz5hID4yHlvE16Su6pvOe4R/Ljexpx
a5G7xmOzfLVvcFfrDyUDvcVIMPjK6SPeDp/u6PB39juyb/81CcATe8+LlDoN9pjXHRZYdTntpykj
GOXkBiWdn6x1lIErRBUjq8AzfIho/c7le/JlSqTYBFJZZy4PJt9oKHxUCrwaiZFGBGhrPCT2Eo0H
vaIZoBUkO04r4v89NIP8ZzXTJoHr305tMT8pL+xiucSmOnlwrvxqELxlBsQaoFdZGaVV5Crsk2XQ
6aC+x1FBbccBNrGhhgtMEXqLf6VPFcIys3Wd99j0R6wopTC3kqnx4PVlDGLvR2iC25NZ1woQaAoM
imQ6xGTVLa+/kAtEXi9Fc/RHNFwnMhpHwvWD1kRJG1KVWM/HmfrWNy3fQ33bdv9+vbbPFgmmcTLW
wKDtSNlVXKCZZVXex3TZreDmzqfxDY1wksCcMzPw9E7QYTc/zY/WRFiW6rzytzoK7ognmfrWDqua
Oyw4opWN5OiVD/IjLoA7UKVcGo8usMvSV7QC7d1wtc+2aNOueFlzOEzbUtLjj+vIcvESkyAi02mt
JMmJjqXGENBpjU+DaRra3nwfcRQwd4RVd5ColVOsZQoeWUoMwLdhQFs3422KiQhqtZoxprv/EXJ9
vdQyLNpkc//IUedhGqBRH8gt6WEmLvG7gj7RDwjhEI8mFWPB7jh9+MhgcoH7iyAAHEiLkw/xmC65
9AgVyXh92ujzteHcwLrJERcr58AeAa9fonKxSqrsem/cklaYX9KDCzhO/hIIPOdJ1aFPXBIDAkcf
9qMYo3Ik0HOZHJTuDPogXbdfbeUB+vQT7GLqAsipTCx/CFOro9rW7OW8miIxSB8+fCI41WHtBXja
FL+oXTqyOFPZ3XTVeQ7drb0amtMpmM+DlCecyau/Y2wPzBQL0BLuo81FQdBQuBo8ggfZnPgLI0h7
QfMMOK+r5h95EdEquL27yzbuN5OSCkFNugj5Clyj0GyfnLsR9LzLX0eNts5ivQIvA1jpoKJEk1j4
RM+mCJmJfoKxnoU1j11lkEqwS6hEnIQLZXA8maUb0G54/xKixXXwwiLzvHJdcaACIeBqHjru9sCP
VBp3rxZARdq3+SirDHZmSA52goNW7aSclgELfstEgLTkj1H2aXrX3vL/jhvqs4ycMhxgX0EfH5n5
HwcNY9NoA42eLdRv4pQSAuzgKI0VboHZ4z8z2M75y0ChdetIvbPLDsOxrPnlwD/l6pIPijJbZfZt
0GmU2N+CNEvoszOE2E+f+2LQIgY0n7k3YmGP0vnOT/IhO2iLT+95T7o+1P2GzMesdua77AZDkP3g
8i9vFDT1DgBRp1z0MFN2QzHbw+10pErhgtZinnB5GNQ5BFO7FoKeuJzxa0BXH5zbLupQqOUxhu8A
TpHCbxqnJfoVtB3C66V2P3rXmZ3Was6CWOxQETLYZPvZKnDZ224n+4BWldDrxYvMved2t2JPiJ9R
thkT0VyvS5AzIfCj93SnKwyzePJjA9h+qkW4krjlx4Jy2J2B7gofVkn2PjeuMsVg7rkqYnJvjxep
fcVgW4yOnzMyGTyi9m+Fq41fIaWfLA7U399PbaCHnr0RXXN6zFG8Ct18m++Ob4o5qLlmVSx7et8P
S0tLlbcdGxxE/xoypw/onB1qZDE+i6PDUNZlXBIpw7nk+MOVBLVhgaZpiTVRDA5tJj4oewV4AuS5
l3vaAH/JCAMvwBDoIB0CIlvNeGdz9Tzc1VzSE5ZU3EGz2bmx78o4itd52dPWO2oAuZqLwP8Awivf
Gw8oKU6uKwcizRK9b2uR7sNGOszEtbBHgHRR99Wbykl94gkEkT+2uVfzQWPvqF1lIAlP5llzABOQ
ibght1SfCVy84ptG2PusB9iRGplXpps+7EMnF3biDyqttpcQxtfKEJ1HxlfkmgLMLvs5zlR84+xg
JmxNzvVBBlHnDSQOjIO3RHQZSHdWiP5Aw2Jb4s6XYwmxORcYP2w4XfTz37O4g8NGZXlP40rgfNsc
Z3E8gMmi+wCp0pGOo0cCv9mRvmhAnGpN+VPXJ6l66es9TNdYLh3yaIUjeb5aAhDv1ykSjhf9DHIm
dZrMtnXFjSDY0EBfjhh1Wk0SmU+c6bHXc3JbULBzpVMK+RT50kJHf3ke7W0UNRq8IlmvHBTvlsSn
tL1ZKbSu/JCeixDGjriW7k54gng3Vpa6LfnkJhVaA2Ahg2gYGy9JidoU/9Beg6iU5K7BSlSZyLIl
IwvKEwZL2BeW3hWvuNL6CSEIOKVp2X/mBs8u7Gym4mJB3JNEP/FPolh8DoqS/uO1Nux3Wv4+zGaK
S/DtB6bvSzThmYBLaRCJ1sUYBDJpb+Qs/vgIeDJGTlhbanSi6Te3Q5QTPGySNyKSc5Jmbjh3du3E
5JHsdEPgCAS9S/ksuDdoQkH2RcxnL817lgnMwpa3oladGHsA7fwzZXGwq3Ulfins9TyXnu7NrFpP
6bosvMVWfGWzXa3W02z4xefriWurxzzycxtkSqqVuU5IsAsNzbuiv2PVTAOcMD7IN6Kbr6kBsYsQ
NMVg5FW+NbLT5yK6HFqvu81q3PJzAPwTiqyHzAeS+5L/GwPwcnzIoekk6KhSf6VBqdmn2/XWyLwt
6xH6tldN/UR1NvQ8ssbzuvGu46QZZ/t9iQ+nS5WtcZqI8isvdazTsS5LUuIWPxYv5P/rYPMLplG7
nT1FPhxedE4rU5qHPL/2lO9LfgrGzcGEc++OaRS3+zbe6YcqlJ9XbWOqtz/hoPBbKFDsuoZirj8B
h+/tL+Jy61VYmsA3xe7Bku3vT4e4FGHT6t6V/fdbWIOppLHT9cyK9j8SnhD6ehyg+5cY2DJ2Bbgv
j9nxZYTFvLmfMXLeG2X1MuEQFvK6y+OwClbduHerNrJ5aIX6uk9a2GIVcKKRuceNOvI4Odk3fNBo
oDLbNZly+VRov4LzF/RdF6rggd+lzlYThjmpt3gjaCQ034ueddjAq7baK7m1+2lyx7rFwrKrj6Rn
xMmL2/7MUY9EpyP7wgEWs1HdjJh0+bCEV39VLt1RhFmkh6pXNYjMoYzkA5soMzn7KYtWqXAX294Z
QonWoktojSR7VBPXw7qO0u4DcradEBJPKxDCXeWrI9NJMOH3yhhsZ9iZzAwEnZAj6qr7gKvzZtn1
1uZO53SA361ZUCt8aO1+qdKuaWG1j8N6T5RhVFlOdCpHWjaYdiTkjAcod+JaHj7Gm6nd0YZMYk5v
Yd0dw25zlUY7eGr4WZQcG6tRUKDrsDGF+jZg/Y+siiihPxMFeHSdG8LTqKPqHUhRTFcM0EBJAd9g
T80aMb8HPXyP4r7sLS5f461Eub7eHjIsvCvlYRK+kQFedsx1RzRfP/LFgyC1ncOrNDisWdSbgqfd
YOt7AekTIxBWhMWaVdsVV3ZH3/SZwhQINLQHXACpEK6/WreIpsxjpU0AriCSOP4FpzIvJruQplbE
+TYizSGk0eJqFBRllAPYmdfYSvsx3OF3bQhByLSW03mny7ewmhlh/grkhS79Da8wmj9vM9DA2RoQ
oYhnbV5AtwHyfJMBMkfLvFGaVNMh+NRY+TRY482ppg2Bx/yg+Jf+iDiFkCT4OO2D05MZkSRgWoHm
YxVkM7mGtUztHnruQKCKuAhE8rPaRBwuuc3qVGLniImEFTkx31Suk8ta9jPy1DXYHeREDZ0hMCiU
26x9JNLet/fOMOakdNi4efSHvLDs9KdBiLQt6/twp1+5nOTaeEJeZ0MUzoTgxmqEen3lmoeLKEzD
d+i5FRb1qNDs8jsIxJlwxuS2Dxq4A3lAIn3UEq+dkZA9GmIBi9mzN1G/uOIIjtAPxgxsUs0boyK7
Acsw5uLQUDRdiBn9wGrc9CgAy5N/tXSnqS5D1bNv+efWLsuLzU39np7tLetVgA9Kuae2kGWrlReQ
kLCg3+X8H5fuEuFv3y5w2K8UrVS5b/SPE/AyOkm+vDEpvqBSb3WeVsQE8Ccg/Jksfc5mNIH4IC/h
n+aQMKmk2bYPxq3z0z21+gKkTVv4Zglan3IS7tf5vATn35NQnzV0ykvPQDSRVaj5+BVVmSfpHqmz
znDCh4MXWV2mMvC4KuQkgWip3MYawOassMJPjEJs/1d2Nznnp+hKTXCJWS5JSmm0lI5s3SCaLD6x
dpmtTM+cFizt9o6Y8upVsINdP0UXeVgH7PXTLYzxaJtODoZIIrfjK7W4Tod8OH9biXWpZL5VZoIM
miuI2+IIK7pdi/Vs40VkSWIaLnDb8KzWpTiB3PqCALD7Rqijl4Q173RXcr9FdPHk6PYP+bPpSARI
dwzkwRIvlDOAGtOR2kLXN9PHHBFdxbLCXQJP6LGv2CPNC71dYPnzUutoMLINgOT2uX+bAgpQ/gEy
2Ki1aQgXqcMcj6tPyExpz5K5WCR6pgqXzSk/Ju9dGZChEd1K0tqt3A4lTD9Eqkjd9qBOwiudr8QW
gFaggCBy6N8INYFi7xu5oippjW9uGA3b0r8h1erZvxh8oNBsATGK4Ryh+mkafvfM/jB+G1pDrOmT
cO3HNNCfznI5/sGuVhxXbGruYctPuWd/PL0TKZRJ53cFQ1coJo6r+V9Ik/H9FcYAsjsezEoPt8XY
TUMj7lRwjLSNBWKSl+xGiJNQ1m4hJWPwKdsAuJBXi5isCVRKTUnCBSadQkH1jsbPJ6QeENe1JE3A
A2HXQLBbwcs7PLDVH4xfhfJlCIoc+21vto3s1uvXf2D6hJC2eWeRhbOXoiZHhDIcEsqly4Ax+cUR
S8uDLEOLZV88L/epRGmb5ti8X6BnkBh5RYkz6wQj6GzYktw1P1dBpdYuNpM0DhvpPDyaahoFZx+h
dShnH70t9FgZWWihoiYatEiBds/kyn3xXU/mLdI/AOuMuCtki01cm+13x+CVuvYHgH1LcUVMlK/i
tBBpqSz7jNUIo98I10/fEhCGoCZ4pDFeCaw76rKckJRgajfWrRuB3ykjDSOqqbBVn+kNSmsFnPjL
XVjqCoOd9q/dxNwP8yan38Gfg+mQZYiKF+8uBEyOeeeQDc9UtvDoTtdlwpMdEPYCfiPN+fko5mqI
BMLRUO8VdnaI1CR5FaovJ/qgoNFYrAITKwMMhjhhraMUNXlMr14Xk8+3wlTTm7qYv5nDhOOUy0kg
ZnW/2WzSvGgRuIdBbPQnWGZuWLbKkxNwtiPspkfY2XbV28v/YwsOGSoN8m+ozxqHSlFCWfivqzgz
plvedHjqqXKLjg+2h+g7LKDS4uw4meiYXs/7XRmz2w28q1mLZ4//CiMLf6foJ1Po6nIBScKG6CRr
A1Ij+hnniWv9WXt/ZutDh7ikwBXtspTct+xkA8+Z2wYglE3IWET/Pc7+lvEF+l2hMxihqCOiTN+L
i+FnmlofyvrB8FbZ69xhpWw/TdxWbJT/u0QVkEWb2t/DkYpjCjGcJklh0Fv2Hl5DiW6b7/OI6f0B
9owBfX+198DTQAIyMfM3LSuhdq1AGa8Oqji/rLx7IYJLQEOc19pBZD7dyPBfNYTpppJegay8+iC0
2dNwODuGSRCZ3cq5EbT8oikq0G58Uq+U6ttcaNsXDmghwLmIpu5nHBJ89j332sWaeiyjVng1jccp
CEhVhSgiDq3AGuekCklbZjnsn6HgwtBKT441t5gGzIDzesF3fPh0/pqPA667divqPVHeDgNqN06u
zcCjHawpL4pDatP1TfFGVUSOEEBpVpWZakRevsgFdZwLqHXYsI+SXaKywsfv0qLQKIrsVsystdxY
K7QPz30lY3F0o47IhuqmckYSZpo5BXLEtIqdHa4PMhlJhThkEQJMEUVMdKCHdGlfS3BINuSGAKBh
e0Ep9WnY/wQNwRWeCQydJK/btuU4RWF6UwMSgbVzMZsnU/UgoFXlhwtc29TmZlCQJQFtQYpBjBvA
4UTypp2dur2jY0NTppjlvgHwgUgBMgRJ+5vXtWePi40CC1CmCq74FuJGRNzbfk1aOnNSbmHm95lz
Ea3GcrGdeqrCQ1VcRntLcsgoPDb/DUCtz0F2Wy13u9y6htbAfpKu2dvABlmC2Xunvmrv6oD+Uuzc
MS7O3GFmKeMh+Ozp6r8qsEJ46NNRdpDzGT0KGP74G0MWV3dAd5J+rFLDQ6WfhoeBnSM2iFzdd4Gv
yQu6XQUcHxajytyqQmvsTbC/eS89sw7tk65FMdztWcpJN8EOdPUUyCEpBFJAJ4JVeEcBn+7tZorz
vj3Fk0CjXvTWpg6mL5LLeHVx0mTLLddxwGabgMRdSPgmiiea4Y7Jfsd9EpTm900tvqF4hNsEHt+Z
cSVxaHPXhMPhbgwtaEgt7+Zs+J3SWERxjm8iGR+apiO3tv05R7hZS0FfPmCRIT8DUtek/t6UVpTt
syR7USCOBfN0OgxEH5DiqXxXBDpCsW08VZYgH5WPIsrz2/0HT8a+kyMtOubRD9q0QmySW/2wVMr+
ulSr57W8G2A1o/PsPoZiErJnHbcqfGttRKTqBx7EaSsoA2x2H5sQZvn/M/SFgwcvjCaSf7b5zKsL
h6/QJ3k/eQalsnmINzXSp03hIrGEi+5yQ7Jc12j1lz9/wE7SAaHE7gcZ4xsDQ7yiXgQ2PG3s/V64
3s7v/m++ewfjNwQ4uknIe3ZTfDOSNgBzY3YT4E3+LNKtewtR3FCDTZ7KgiVYoxdHulUe1QU6c8HG
WYpkb0LoMt7vaRTfAjjS2WQsptt5n2QoTntQtIKstH79mr7D2NWlt438hFxeJZjBJuZhVEZ6jaTl
J2FR9KBihR/FeZTpk6evzJ4Pp4ZCUseNA3SmIHBzH+MfGHU34WPel/OKJmC0b4q0JrbBuiHwsEmw
XEfPXfmAahKGk5ghAWJfZ7dmZfwT86tcgvKuVj3vYCT9gVSWB/XEX1TUceUsBSY4PdMnEXx/GJNf
LbnveA0RypCBPjhZWxryunCNJPGbc3NcxJHcju3S7keudmDsxNG1SqoaKwQlPwI/cx3YhQnMXGFd
nD7VRhZzffFmrKf6i4doYXArBTiRDUHEdRB3fAQKFieLmEp8vPvm8wEfUjIiqTdD9jNYgGvWyRNW
odfYVcC+XiPzqEQBUarBvnWwjHI1ul420uf3v4SIrm2vwcJddYpZRVD3b+FUCKuwFI4sUgONnyTq
uP/pyurg7dcqkz91dWaYSzcnoZC9rQdsvOIrkz+7M0tjec5RTkpsqsskpAYjtRyVKgBw5FRKwoBY
U7uid8LWkp9Q0ciVoKkFj0p1dVcNoMAS5GZNEYzTOFybvJMgKGshM3n4UhFvEIaH3MG2/lk+lW2o
/m/5Zt7Wx4xoMCvtx+xqOdFejSR6o8FMkbB/LyqDf6tk9GmgM0jq72oUvv5QBiXqPcxllnPW1Yd1
8Ym1LLCENxlGpunr2VgbiThWlbTLUSw+yOuAUKilxERRqpWvyON/YazGyPnksjJQDPJrqsT2rjmj
94RajqM3gwA5IGexoXObEiICMzPC0eSgN62/zMAnxWOb8TNocbGGJLAmEHmZgMF+V5RIqzNHUL8Q
A25mLryFUpOektqRT96/ZkOC+4nVOFGNoBFabu232cuBA0R1jV4CbslSbS4dIA9XL+RcOIuTH08I
qG3WzCjQuIeIwx9dh3s57wcmrkM2/tdgpibRYbiIURjagu1+Gb8wT4ElBKgeeVWo38mq8tAJmF56
edYuTS9jRzSoS7tDRhC5YLgUFAM2WFJiUEkx+4tGc7aNKrWr18lWlpurpEfvufGEGmxaiAbNpsfV
8w/gmRfjjgqF2udor8dNQeEb/urvewUiIITlrs3YuLBFEhMwa0Wij9YcGigoV+ZFF44ak7bivNpG
Cvdk/VtMQ2ctQwgOVQ2ukrlFSP7s5n4ctlGpsY9vpIaejvJFSnGeqZl/IIVPfEIftWhxnLyy6+0p
PjCX7d3fAu9tolk13VBVxpSfae+eHpnaTuieb+HiQ3kDHtwcaBPoKscAOlcVQxzMnAHoBPCjEBEP
7dY/IOu6ZjoXCPvO0/s77ZtkHrbXRJFdBelp5MlDcRA4XkQi2Y73FnSEytrTscrOWRxSuv2s9Jhg
jJ9t1t8YQHWqq/g+E/bU0qDBS72/sa8yOb4Gs/Xjhv2aamMC/jAsfslkeyWsaDqzjmlG7AI8fLdz
L86wsUPBhqmoputnEIJtKYH6m4WRWVuY0ijrKA2hiRbDCh9IOtM84HjCNECWqEbpLoCWRqLUQj8l
kC2vdHjMasBaghF6skyoPiYkdZOxATZETC2mirOMoJMcLRQSguS8v2foJPaR/LVtih1yzolnmRTV
AkXH81ue0Zvd5tlE3/bLcZB4kYaDHce9lRsUYXECwoRFMP/wveoyyQV/YDCHEOQbccvsQc9mytwd
i+6q5+I4k6VPtQWVV9oHNKyufx5HlnW9b8cA5LUHSFkYljPPBBHpZ3ME9WKBJ5EJi/RCHM5qP8iP
jt9ATfPZbD2Ppefqk0h0aCbn7QRn+4vYL6KZUQeLvwX1wtgxFaQOVfDJ821vwmuZvR3wz2YvxKdg
QQpO7IkAsNLnc4LWO2IwoMi0FkNVqvMdsuu2qweu8ymN5BMQKnbBZNCKyuWPYHlaW0xec9P9WkyN
EF1ClDwhDyxo5R5C8mtzqRLG3K+0TVJvxSZsHenkS1tcs5SkZB/lismapQJKMaxYGQfMc/jDihAy
fKCtPbfZhh/jDlS1F0JMnh2DSNCfW1VrvOnUIPnSl8F23PFxFt36AHdXHOUqHu4LbVAM+0TdQbIn
RjVUxdGNx238NyHADFns1DiUa8wV4W/ngnZWhA+4nMPvM5+YMKuJU/iHS1gXiQf+2mQADcYerFHd
9c2pq2cT2bBS1FTQYuYTBhtRsfW+tlpIxCA6lXPdGUQsVQ6GwpB82L4QMP9jthknwWsQvmMTyMeB
gMxSvIGlV2eNRUfszHWhrJlgz6KKgtBlV1EYglERnTNvgxYa3cw7ncsmGFAulgBGHPDoRp8rf18Z
h89mKroB6uJNZ/LQZuHhMUMVBRewW6HPleRLPmlZU+d6qyAbb+KofercYunUbhwdN+0QnKjW1EAQ
hhJ7upe3KIlq+gkDXprFpvguPkogH1+mnqfTqlkJXrxVXpZh8rBcMZI+uFPJQzKIPRLPqYJRWG/i
QhRXUV4eWIjaanAClNEbyCiFzigFa66JnYCUDIW9ZoGOP8Whh/EuKlup0mW0sGqEd9j1MocCbnY7
5288/XKWUEJulqvGCxTO0Hxf1ueeMD77Uugt3hAhquCn1hmPmXwCSgEwHpP7Ot1qRxj6Yme24Noo
z5aZBIiil/bk7rFammKebfGAFVZ1g9f0pf2T/WukuOoKVSqBup+09WbPDN6sQSlf9kL0HhIkqK6X
gClKy1KW7cfSr1QoR/komaO1eqWgVd00fU5Z9zKOCmTUrI1+v3SfmFP8LtYb6Hb1E9+hu56x0vWl
HaXQGbtYKDDB/IF69f47nwDDolShM/PqI63h/tpF/4p96SNPI8Cyp1WktVaWLdYtsYjm+J2dMi9w
4WQKe5NFpYcal0vFRR2/8rdDmruQ1YjogMYGxjVAUFLZ6lbq96abX3+nCwfGPoEWdEO3MHJxVavp
dexsC2nUNoFj+quzQ3NRz/gZ9AkexjStlZFbV381ehWOl6+GNEH8+Ni9Z4Tqd0/LWlSixfdXkQ8r
uPSBrae/GZ/gGwOnqiCdX+CwoX4/bnctwNQ1H8cMDQFwSy9jj7DzLMB+r7LgI1XzkqAvsjjBbllt
ct/odj1v8VFAUkKmpmc/KFd0sAhwxmTDiYEa8bshKFER7v0sEcv6Ioo/MXZAvUVeOsnBi6tKoLWs
9MLq7+5DP2JOW6qXKL7fSZBKpHV27L4i9RsWpdkMW3Cq8MuyYQx4hDW3J9G/+SbbhwkUrzPLdbSm
+XSZNJwcAXfKmnSSAuHhyB0cHPKv9Fr2NhI9TeHLm7L1O2Klik3CF+Q0ebA/8vtGQhPyuielbCeC
iHmE8Hg3etdrjAp11v7+JS/qHwQu2g0IN3vjzIEjq9/rePphjgwpC/cizQF8RquCVS3y9Sr7vcaG
SAaH6hHYBxegBSWgTS9wUKQRA4Gy2dTK9WbzgqPNkIK/RxRsbWEdY4vPBpljMgp1dVcNVO12YbiB
0aAzbvahiP5RCEckz5kwIZz/CesfNFYh35oKvvVrGD6N0L3LHyj3TO6a/M8OWYK3iOFhglq1xvNX
vYOWUBglu20AOJp35MdI0Z3l8Z3x/2UMTyGyaiIgtO4EKWuy3p3X+K16rwzykJ9XX58AFvcOHHSY
j/tbTBZamvShEWPO9s4CKW4l6/XvD8fCF3EoKvWqA3dYXbSnJgx9hd+jLFJe85aW6geZbijj6327
SGsl6cB1+OSptoaWaXZL6Mqr5VCKxtthARzZoZpXoXomAkG5d+k8MOPUeDtzbDdfryMYLmpqrekN
tWZC2lpEl62yfn+rXH7+k4M6EiJjc8vv9EpyUbceZi0rs65wwQ8hC2l2ZcWG2fxdjnjpi8bIq4uZ
qz6rIYwAvIbIGuwrHvWPQjPwpH64poxvyfkes0JIC5t2edbp40kqnOpVmyLv8qcXN60gTk6lt9MG
TZLw83iGtUm4erIpbv2xDOH4q11YJZbPhp8SpaDS0A9IZBQ6Vw+orinPacCyt+xkVVYRGI0bGN4+
RAyqy8KhEoW+Q7k7Qxdg+o/ugvX7PMIFXHWIzmotXsTGfzGM1z5JMgq1QS2tVOJ85JL353HMZHJp
x9DshXM3kpqTf9wiBZmf0s+5Ty5P5Ab9iMJRJH0nsRN7dcqZPn8Aeq0pTiQBFfijabWuNwfFLbwk
EimCg9whHsIgHGTcDAAZOff1dbGAzCE3Rnmn3QfVcP4eCRUec+ViQ03BOxtI7PLg9zpNWWZBIg1G
eGmkbx1X9ID4CvHwDPuXnTp+uaWzFb6ghVzcouXyhYfum9Wo2OQFd2YQYBUaSrKxLLufrcdhiVK6
JO5uCPWsgmJrEDjdswucK5o2ecxIFiupe0KVsIa7mlkoi86kcBt9Wo4ymO7ALGFXXMgU/sV0rs5g
U5gouVK7wgGfqB/EmcgbTqXxBX2pMj69/aVkGAhxl4rgfoylvg+MoGj5rMDctwfKifnbGIn3uaJ6
Qz4rXudryJsBQmGJgkkMgte769jgQgt7nQ4SwtxHSc5lzGCGXsuGtF5/KNwD7hch2laEIggSGfbc
jot1h/80sozHJY1rR9KSijJPSasD7Y3Wv0QSIjvjRqseJSf1K4LT+U47fBa00fovjyksK/MJVcxm
ptVSvu8lpv7t6MLqI0jF/rqvmxxCfVby89eWjcKcku0YAJttGXMMgPrOGfEAPKWqgku0PtshY4tf
tJuOGkWPtyH4H+vKF5+IvsPN8zt/UMJ71x5IOveUjrRD6l+GgKmhUdoRZYp85OE6On4BWnhpVeFX
rFMystkbdZ+zpaeuVO1hU/KO6XZNB+28FLd9voVo25xrMadVrGZP2BATSTjHTlDYDiQAqYh+BBm4
bHLtY3TOZA9qBuT4dWNUwmiwAXo+MQC2ObkNyJ15WxhETGZjYAcSCVTCInnAPyfcdJgHDChc8RQX
QM+1CYj88bDYpUBl/yMUc9goYz+eUG/1Que/Ok9Xm00chn4/1ZZ+YZEHWpVg0Vh8kYwz/8N1aEgz
mPiTOtMRo7MdrpkRfJfijOVPqgVvidmwFkKXa0pfenZY2dmPZyGCJSLYV4Uh9QDjoPKTmfd7y3Nl
+p52uVQxduwk2chFbOQ0eXyaVPXMXgRFG48i5fWPzyWmJSxTRc7i/CHfihSgVYQCuMDjUY5GfzMY
EavrkkFRFXqdH90HDeLJ0iIImq0JO0f/shxx+EBf3SzgW0466v67uzCf6B4y6YLJDvSmRKfloZnQ
4Ucl8sGQGKi5+5LmS8LE+oJVkGpjTJKcCTVoEdGAlVAMoSRsi2aCzJ55e1zhMl4RKs7ivM2Dlqwf
RXdLMORVc3OyMIYTu68DOktpXtLDjB+WAO+PAUPiDaKpHladNllcUidMi79wvJwrbOKCbmLFR6B7
sqeP+WgtJ8saF5ZbEPd59N1y82yMYP7pe7PWFF5a/u2lzw6LXKGVjyC4r+OSobI2g2Y99EUalsqw
yOhxUIzuEoYbZA7jZ1QlHTi750+Gvf9FPs0wjIrciLpANHoy47HyJfGhRmB/bZY4kcT1Fw7XzSWh
CZcvf9quLGOV9t4Vxx2C8m75rzQ/f03lY1imbd8//jb2nq4irnX0U1t9w3XLYpZGrHbUzKJcN2xV
565IjDyu2Sgn0ZhnCFB3/WVfqSwVr3jiTqOCwmydW5HxB/MoaLl/LFEzU6EJfMDSpIo9OFi0KuxZ
WpCU+r8CC0c7iZXkvWKEtAA1wImtmT/pZTHjCFwrJIqYbA2IQkiqj9PpKJ4qYzFHzuCcg4HzV+xF
YDxAZiYefEW9i1Ls98C14Fozfja13xUV8wgcQXjOzzHRs5Dtw3UpDmMICiBN6u7BfZgmEd0lZpYz
izkdrsryDJ3Z81OvFYqfC4j5UMUG9Oy6yIe/7OUosuW7T2rmEj5Jlw1n+4B2mTvNxwtBt5SWYta6
vfV3n+8OhbNmq1AHfm5SuIATkQl8mnQkNgyW91qjbEWgLqXaIHPU1j6/I5TlaWQiqb9x9SXk1SNe
iIlvJvXimLMT++HCFpV1X4mQ6s3CemO5DO2lBF7fpybV+mOT/NYQruONd1yARh1JeDZQTuqPOHEm
h84mRN/X/NZUb2YgDQHUQCtDqoW54II7yyOzk1RdG11xfCSqEu3IAaPfCGJN7jT+/wSs/888Y3eC
HdW+Sex3eCizG2wPNakMlCP/y4dQdNIlKJaQsk54qE4J9FTirVrfyyGlycpYRUQBBb7pU/n2jwwM
QjfCJW9iRd/0ZAqfyZrnAEyIcQKYlX0xVBYJvb22O4Kd+T4a9ejmMPYrCUS4rCiBURkEVD9Raegl
yxvvc8658CM3ScXcwhewTvywJdkVI6UH0kDRN8Um4rFaFsf6wMSZmbUNHBOY6NPLq2Ql43SS085q
3ewWcXe0Xy5hUUBvz1J3xAIzoSFVOVMQXc83q8CWaobM+GMc9W4C1cJyGxRwUneNoE1O/R14Ehas
D5hOkH/f6fKuqI7cA68iTbTqEAtWBLTso57Y2WDr7cWcjuugYa+BOlbNqA9+IFfrYya79Qb0W4CT
Nv7N9W1YfYRbokVIzDq8SlEo5Sc2OHQhyRt9E5YxdX7ROqaRJ5MoYEWgXmRaw87WDt9KT6Wdhz0E
8eLA1CztqejI+nrzgeSsp4kXqr5xm6kA6JXw0cHISzv7HomGZAxnFeShg3Dq0dhfnFqzWzealMT7
kAyqU/twNItR0BfSZc0dodAny81f/i2PZBFmioPmGgrGFumOeiBgYYbVYPRVR/CM/Mpoxyqp4MTE
hf05Cj2GveX1EZC711MC7w0Z5a4LRwBUxzlThL8QiyyyIQrNgxikHn0Eo68eR2jf83tkf2koaDPm
D+pZHrTHmwZViiG63rUjEULxrKdDTRz2EcvP465sv4SAIQaT2U0hvkMQlDwocacoJNIf+Ldcu5+A
Z+a2gOHV881PLC9SdJ9C1+4FLjdOXNZ0jSvVBFrvPxqFTeS+oa1t8+iul5UIns6E/XaoxRf8Yinb
w2TeloeMJOG95/y3xwie6WqZFacBsBlysLcBrXSKj6yG0IfBGuNtahIoXZtjDN7zQCI05Zp2zleh
qcq5pFglKRCoqrHMGsS8pgMigQO90FkDKDb9AgjMTLXx4zyJ8TuMBneQlmTf9Mi7XVEr/9XIS0bU
jQ2WprTeoZ7tN2ZIRlcHQj3tReBISIwwgRDuvSJ2chsQrLTTo5tXnSkMVlAQP2qlArn216af1trH
c1vIclys5B8JK4AsFK9IVms2nBkQXVN/ET2aPbpR8uc4PeGvhOVK6jB1W4TyM+kEJuSra/A07/yd
N3Qs0ED32xxHhyeKxVjc1sWXqWOWng1D8MWJO0QvBwbkJ/1K+gqAYUbs6PEL0it+z+K1dT9Zfx5f
PAUgrVMKRnO/hTbdNmsVPT3aRSFpv7HqjzbiO/7YzZz7x4gHc8+k9q2ggRznnG6pAPULkwxEqDkq
U1NrRNAUTJpezWkQGu9o4F042wDCPHtIILOxz6IdhZuDV3OCleyBF0UXboP3nJAbFwsxg46Nvz8H
P8nrqYo+WiNZS+/7KWgqj0SMytht+Ueb6zR6/2hRg0Ab4Y/f7/R82L8GZFInXnSPPJ9seE1supI4
NodqbiqjOBzEQRLhBJeD3BlgDHh0aTcsGtUa3CMh0AQl0oQKSDPSFSrB6T4ULRvSEnGFVe9OPh5f
BEPR3fodhQ6ljr2ZgP+sXfmmdfyieGgoiq/42oIGZUKnzhr17mLrt8S2MIiBDWiYiR80H5q60RAc
udD9EvzGuOgs9ubfMVKEbbgADb4v6/ULoegbTo0XypFWOCYvhEGcMQIt9pkiaSSp+rcy0ujoZE6A
4sJze0hiLcllihJ0KscLWivJTMHwB9J/OkDH+ia6AGV1J2jlhsjjKbqF6GZUm6zz5SJAaXwV4FX2
UJov61c2zd5v3eQMpYbTOOgtbg2E/Vd9eCVPPKw1W/skferH2T8ODGzXMKCm9jvjXCbw7xedtC5E
rNT7/wcj0pstkha64Y5Cu0nOp1MwIpR25s2E0W+ve8jvxhYAKdDIvaNrbKvAbZkJtnxK7ceRxWMB
VKhykYwdnoodOxqCDweIAy0/arrzEsnsJzaE1Lqcey8byulS5Z0ZbyjmGX1PJe9K58FAzIpgu7PQ
lnuxhvzTu8fMtkXd3M4+V34EYILEgXi0TMeG1foBS48/HFtQLJzU5Qo4e9JrTIRoGz2VxBj5K+6i
R6JFX7v8E/DjdQzV04zs7nE4fUqS2FXvu+ncS3wykoLzuJ/s3k9KUVsoUVijj81770PfyxLJ+fgs
vvmECfuOipi91v8xp8J5/1MRUaCicw+76fkCVgIdIZovMFtl+RKcQSopMHhtDn3OFegrjOr8b/aT
4RwM17PcUCajk1ww4DzgFp3PPi3SpbbnZ9sa7TLNREsOhmnBEjV6p2Yvv9B9/MRPBx/SHx8UZJqS
dzWxd8IosvbEJquRZLYf28h62TTy7ovxCSv4u9wutf7Q0j8Gv1t8g6Vps5CrK+Dibv5CWfd8qCSj
QjSzJWJkBx8Xx87Rh0e8FS+Q/4mmUtOAJdK9kszQdEMzV/mVFsG69uqbmkZs5VndBsW8gSC+qokK
6m0avr4B/3vJ3jNMy1Xt3Ctb/LhU/13jvyvWh7+xyewP/uIwulvVy/vqGjbpp2Y+7DhOUKAcmnPO
VC+e0dbJVwhXL6CiXtAICbKq1L2XtrcULEqXY6dZi6pL3l/gzgolxBdItKgdAt0txN6QgK/dxtPT
hQNXznh5dz1g4OKjKT8iZw24/HtZAil/sS5JCerQ4cpgAbC4UN3r+fJSLBjhoJrrR3oe77cKR/rz
dxBV++uLzAShPA1fxBZ0hpvJmAsv/FOLwIXhJp3n9kJCZPG/Lr6MKcq9L8FXfbnh2bx0cD9PlZex
o0UkCFDEfyHZyaF830a6P1pERwi9Uo0U3Nbv8N7Ye2UFctbLyfUE5eHRuCEE7/M0cCWNnX7FzhAB
muC65NU1VWkb0WvgVeznBaRbrHmcTirbm6kn6oib3/0W5lumk/9InyUlR99WRFJnWbFLzSJNJDRF
l/S4nPLIsK7LfNdqHfiSjPvcRyp2vNq1/k4xc+xdse1HSe6xbTXgbo3DHm+PaBedT0ESgYbZmUGD
h+s1Ry3ofOzg/pNgRw9Vd5PuCbYf9D7RKRLYA9NqElbQSRWFMgL4mLnkv6JkmdEbkC1XsKcmbzuW
Yza8yRz5+S1y6X2p4Rloaxd7NfK8UgAoXf1Ix+FkqUvDmb/M7ygG2Tj5BxB/PY+SA6PnEaz2uXhd
VJjc6fQaSRoJcFrxinzI0xXgoOWgN+Zsj/Fjj2qm53F419WspInmzkOc5978t8e7UYbRXqiNW8ng
MWhezOpQ2Ep1SoiYhr1dbx3ohK0kA5RsFdMJk2YFqG2nxRQq2G1O7CbGNmIXoPhS/XPFEChvhHmQ
mhtBv9Bkpn7X5vIMM9kEvkwxm476Wr0QakOu/JsD+fqI18ubXWFD+EMreaCRRQxtLvTdfdA5xMdg
rq4mRjA2fh7IaJTlZW3Fn4iarxnUafu8DuGO4LacGnXrvG4PEclmnaGziKQZYVB4weOM4cDFM9tY
6am+kBuXlq2STyf7M20cCLfUTOTcW3KM5CfqVxwxdvQCjsINq97MDmxs6mgkDnCMuKqy1c8SSJR+
LcOwa4kV5jpL/Oea5cVoMc/wMSaTVUZjZXRaovIf1aiWVmUaerBit+/mRYrLNkuXh0ppg+2aavcp
JDILAjJ4IlkX3QrX1A0AKVy9Fe2gSF/GeC1/y6RYc+ppWsJ2XiKdDFxFEH654TarUKpxRpOFlgrY
CtyZiYwwpU2Pn985jCXdWZCZHWR+/nfIMNquRX8yh7FXJykchMZsBTqYofht7qh3yWj8Vpv88RLS
/wCzklTuY5xTZecxh/oo/bDcuiKDAfgn8dLjvCPDZ0fu5pt6odCajosulAsdPw88EnUGK+YiAqWe
ZH6/6473uTIgiGDmKbjfuw0uV3LFvrbeSt0zyIKK+LT3s4DmBc/7mhUCkr/uytYGcCDJ8mLYgIAI
o0uF2cC/uSFVcEi1NopJO5iQbAOLoGmColwzALywWcpXHsZ3qtKL2klM4sDRXfeT4KG1Pj0uFbRf
nKdGhouMXOuAo6A6Y9OaLUhR9aJeRBbnGl6TLXmUc9P0PdgIsQxFBgQsMX95pst3nildGLkZIQ00
vL+jrbUkokI/bXc3B5mPHEmvUAQyr/1zW9/JxX1+2cxh4DZxPzqeRm/MtA3cAJ99SV/M2UL5wd1Z
+l20pKaj1/L/xvJepsB5YiwmGN68KGfYV06zTD5sdecGeyYT9sjhq8ZRInlvRM7XA/sjhE6VsXYO
e7e+Rac5XoE3JiEHHqmr0Dmxa6Pzp2eFC+GdImYJ0K8czwkSj9MjfkX3rs/ofc+tmTg+dri7a7RS
t0IPtrZfokzOccJcmNJI+O0XxsSPjiTSSW1sVfj0zfAZAmK5efVmw+flfI6bE5TfdWemRCiGkEeX
NGxljhnvwIf+rNredHD2KmRDgaHAJVTdn9TcwU8CPr1EB2wOjr6jPTe8X1iAQOrRW+Zi9m9ciiNY
/WOQX+EQWi8eiNtpzVVKFfNhFJmS3N9jba6bYymW8ODSyPh/XuD0lamlJymcywYwe2RU7tVrrR9a
229HCcbjxd6HoWS6bbsBtFOMOt0SrujnSpHJq0jL/jSXbp7ep5Q5go9pwungJggvDoda7BuVGTfm
31T6nldqC+LrXsdNAjl8qkfSOIjSfesQdvCfqxSGTS0ys4dqCSQuUly6pE1gKgA9ZsWI6lBPxW9Q
Vl4s5ZlXVCLrjYt2BSll3AizUMjat7CpIfdQ4hiIjWvsdR2fiZxlDSHtNkvq/G2PRMWWwWOUYv3V
P61JCxW1WsTesvCZUt8X2Lfv/GCk8Jax9v16DpSEkyukl/2B7KEd6Cr2GIMprhKZ62IAOBOGwHVg
c6qB4bLmrQzCCijN6PQ6+flCBpWF4qoYVLeUgrCTGJ/nJXKfDMXyiV434cFYORLIPEoaenFBrREy
4O6qjEstH2S800iA9AZlMd+BrAYB8mHb3d+qy2FuLh0aPj4r6OMCQ+NoYp29/H73XJdTgNBOJVSV
s6fPWbGsymDAy/tSQHbOWGR8rebaOcXU7MJoM9fNJjRMT2Hl+85kQBu3PauRo4SM5rsyBgmJ5Sgs
UkBS6soKcf0O7+3mvNk48w/8BYREqxdS+LzVw1KvAkIeNfhT6+VvryEuJNMBZj2PWmW7axA37mMa
pTwIHn0ycjFVFh98eqf6dPP3XwZMI8q5Fiy0OQJGp0rZRzO6VN786wn2TAZ4/i5Uo//PpJOPXSRb
crGMRD/Tl/3bu4QLnDCVWVoPD4oB7aLAZ+jQf6TaXMjDEW96b+1ePKNCla7LPTxiOHorwcGcfpSK
qvSlpLquCPDw0MQSg5cW2SpVZa1dfsx4gToq6XnGleHUq63O6hOFTr4DovgIkTayKKNwvTneVVip
g5AIzcqFZm6zSrwUK84erNMVBYVWKMZfqQwALi6gRTWRiVnldd0LerOO2PEqNHAv6OXEgSBOhevB
Kz1cNcZg+ZfOcdmaZH6gjH4P9Z7ItJwjxt1F/RW+l2Fl2+nZAZzebKS2vJ7AGOXYf61IGAOqmD9A
GGoiYPZYCpNi7TdFgGmIjTjXBr5eMKl6BXV+Rg+Rxju+4oc+uUrINZzwwRLf0ixkUWbratS/4aRi
kgJArAuqthhF6XSvw7wa51lz4XLXtPacedn6C2KDTVsHdICEklKU6UzDvnftMpU04kHL6OBsp/Gu
Jn49BHz+lZ68A13FiCPe7jndI6Ouc2bztVYn2IMgrb4YOGLGs6OONFHucdLG3avC4bi0cAwht7ab
n+LDOjkFNsGfVJa5Ku/RUZSMUK09BCGOsg5W8V7il+uEEeNVGDLaW6GUscOaxB+dSPg5RN5p0LAe
6gaENnJs2F0DdZ4ps4ZwTgQQcDwcspL+mmzbx25XZLap2EHiFhcjlD8YIJu8Zg/0x0GwfUA3EeXw
qjDZSOMvhcwP8kZuhc6BvEIEsDkeEapVAX50EGLjY4N9mZBe3t/tWwqQz2raNTSmnSzU9k00T2qU
4m0hRTwopEs6IWjobjP74jxQOVUsI0fkmt++u+z4Mcyw5PdxRMa5o8UNDzQkJNVZSYZYmkTVJW/4
fV4kKV6iEKt9zhXyicRnBgRlCiemdv/+g139CUjmoU/1W3K7R09WGyjDJZcB52Th+6VaucrrlvLe
+QrAAlp/mq2KpsQZMnxEnEzZvHXc8RIAR+XfLpcqbP5glvaamCQIFOXK09sBphL/7bIu3AoBjaPK
f2zbOXFSxPi1aoaocjef4b0cw/NKYSt1Bdw/EjmxGTEgfri74zyL7xoOqW9dSNoiJHwzXHUdgJoR
UcCSol0yVCacSnEo9NDlEt9n9O8+kmgLxQI8BoR89TehMPXHC25wI7wNWXhVEh9ckb5XgYyDWxzg
x6lMwG0BQJAYMru15wjee8rGhYcgqIRqnkM9YNljBVHFXCSzO6rzSMAir+YNmSStx49Tvm5gS+FI
duage5rrYd5iuI+1xgf1OMWmkF4zT1q0Na3HdI+wZLV+wNJRCdbkRJyYDQYUXlPPHUOeyCGBn6pM
Rnt2HqfcKexQwumuDHFkLI/E1S1FDfrtDDL6GV+31XReN516eq8o/CEdqtkTlHVSU3gs2Ix8854S
M4wi9d/M0HMBqNIlmdpRQysSG+gB8UJNUbCX8Gvme5RVEEA0Opy8mvKUIUyk9Bx/+L9hXMg1kkxG
iI7RBjzEJ0zRwkeYtNb4A2QjG0YOMBi0PxIKiGkxBZgO+WN0ClbL01ZdJ3cNoVkVRrMV8j5aSuBj
vVdr7tC2hrVpEDfA/1Zqm6BkMRYQijgQNvmSDrmM5bITq8ui+u9c/aAyDfCfLK5mP2xCjtWSGRQZ
uh59x/cRyYhq5Jb3zzy5kPswi4eQ90bLj/atdsY2WIkckReXvf61dgW+l4zJNxAiivcXpwp7XJYp
dwJ7mA9cvZFYAScHkex7QuSR0kQo3rtaWfQwInW7JKWRTHDtN6/gyJw02Uw+oSQ/fZorFKJe6FG4
TCSQqvmvMLeExkQoTdZI4sy8r6QI31TFQgKOBQNNYKsNQn6EHVYdUlniBsgJ9+upx5tKn0K92aQA
hOnfmei+4cIH2Kh9YB11M4kkJaeS5o0P4bPjMsDQrqyEuLLWffcFoC6qOTylDasvit8q+lRvavAC
ghyBrBV0E/24dhx8ZqRL0ZeKuxknWrkCmsdvAVoJXfc8B8F+2TjlSh6fjjJjetzFDpRaqe/kEgpR
vupfn6WMNdv89yPFe4/Q+NN/VG8jlJ+WK8MrfFiTNHYwXO5zJyrDZbMEeFeSw4MwF4xrdN7NVzzF
4bkbiTe6mvnwYAm/QBccTv9Ooh9QA3qZw6I+rDNa7ojU1T+3ty/GKUpb/7osvOyBEPODEheNZMhz
UaW4MNHGm3TUEhA/Hc9n4P6JT1CtUCB6RduxbQaj4hQNzdVdeX6mMahGRukeps4fRlBedrqwJNr1
r2Ad+6A0l0Ao0ZSK9+SW8PyocrMGEmL/DZOqJ6QrQmm6uBvxsqaO7lI72B9EEylVP7o+aodMph1m
D2D4IXcG/jLbWOJtTv4LuqHj0VX9r8iOCE9S+XoInJR8duPi0hAwhoTU8dtkFqjna6J+CCP3h8Vw
KxJPAXMTHkJx60WZTe6DxfjF6h4edvJrtmy8SyVTV53OvKtRizGcwl5uonoVq8Vz/TOto4IN6yXm
+APA4IV7UvFw5UfZD1x4wAoEG4ivB+WGd7rVjTvoB+eTc8CyOha9fZDGzX9BW1luseR6E4n/MCwr
CMRGVW3VhzAbtuxmEmVdIfa8apF0s6naZxa5OVoBsNnPMyES8O17/SNO9VUUZTHr/MGXUJs7LQQe
XahmhNRoFbSuhtLCslR29Tv2iBQIOsnkuLD4RKXlZn/RqFGDIIgSvfHex9CKaSnainfc/m3Pn3Rs
v6N2rM+p7GhPuJ0ZmFH9b+ppIFdMJ9UqLst4SO245iO3GNv0AQzLOhq1nBmbM3IqqNI5EhYQ9crs
k7t7RWC0YQUqMl+W2/50pKQAeiBlOEgRECjejAu0/q00PpGz9AHsAbi2h2D44+pClTbsALv0Qqmf
HLVQJv2nmE1UKVqJj1dHjad1/98v7aA9R5aMB8V8RI6QO7QBg/LXtSiABWVjB8JwhxyI3pvLq0Rs
VLZmkdZyVhsq4U3hBstxMQs+vY08YkR+nyzQBMam40NiynwgTOP5Y0oCfW1fCbIJEDywXlIv5YKz
C5o+dvgnvlBtIbnHbTkkIw4gmGx60db294SmrhMR9RWGTJVAteE6pSBUlfiEY6bFTaVYRuMf5JTo
VOcpOfycOswD+ZDGuEuu1PpHWltCfIxYptpVXA1JqdinOf7t5E1VUvZtUTZ17xP9OZi0ccb5Jsos
m2vkcMZA7J7tcdtsiQ0rnDRkYzItzn3L/beapjU3liHql9USpt/dOmAdfvHL26rJNYmaXkPGD58p
9Kc3Ph3d2XDvM+9YM0Xifh+Zig+q+crQv2K6vPaCXloceMUcA2Lb815VUGD1RBteJg90e9dP9IZf
Jbj7399mkqddWWr6LM3zXegW8pThzUHP9xv3zBQVe/3xEmUi/LH4keA2a6ylW3egC+RrnmoeE7xp
TbMcC6rkWMeM6NzHgnfQeo1rOJ+DjKmmEKoNd5RdPK1qBBE/MBSKI/PDQibg7Qlt3aQgOj/RgNyG
RxGJ9VUQHwe+uM9f6nP2dezCUoFYAsulFMcBODCRVPY73HvmlG4p6I8jJfdtcAgNNndp857hYMPz
CNy/UU4AYw3oxIVx2gss718toz4FA26ShipVnNGzNqHINehbsQhBoiZaZlywIWR2Ex4kKGMN11ie
exWN9kANQnjOfo8Gug3XpM4pifIYQ0+eLa+wHil4zyZS7Dn8bxDjKVSJR1TxWgvRSrDOvVrFjD3N
NapQODDQ8NB7hglHJ/nsvpG6tijROh5o8B3ElttC5x66iX4dJz5SXoKh9LHqEircEgacVUzU32Ve
IlgIo1zXLV0PIRiNkXYdJHPRLFbMLkmm8towtPsHb7Lab5BWKX/0HlKMNMsOh0cJ1pI59OCfix+e
/9ECQ8hsjVfY5UnbaFL0w69V29Ugyrz9VoBKvfh7RT4uv7rBX8IjcnrbXiX95reFaPDowHVqJZ90
e9c8sGVypJjrYtQEt/aAgCrCMUlBGCwGIXhYphNaxj3qagtz5O7BQRYn7TYnXFmnMxRGVz7nWXGc
29Qvro51dt9hyS0Y4IOGNTEU3wMnvQFkW/0ZqOYp6ctm3rPX2VZCpwgbWHmS6RAykPZugjc/JHmP
U384aX1oapA/I79tu9ssXc/ZYJlio27s4V4Et5UvGhXpfgXWvY6QMkdJjoEhzvYO6s/o0FVe4zar
Efgj8afN2PugOHjOeWTb0iVYFW33VqzhMCuRLEF7oRHh6HiGaJgN8rC6kRPRiSK7ByB2fqvaMkUC
bBzHLCD/PXgBqmcFlvqtHCX3yVTB06KM0V1c1/g/Qf6/pWSfwnZrYf9wxgDLGjNmIUQlOAKR6/+S
2SvEKVK6HNFWAjFz6s3UauVDKjjytpsD1+1f2VPjU4krSc2CyHxb5DUHHGc7+7pno6QfvXzRe750
Vc/DX3P6nAvYwD5g+vk+JdpHkmIM7Aew8kQcGtTJTsBgdL5hoDtz/YnxnTB1ao8epbxwYXVqjKDS
PwAFT7Gx7R0Bk7UWdhfv7WgP/IJvYIpr7Zhp2vy4Z9sl9+874QJYL0jjs4gWibyhpVwP9LmvMYI1
2A+LXvqqhRxvk7yXNjtRlfwAbM38go1jIpMVNNYGRQG4caQtnoGsANjbY8Q3ntrfAyaFc+BloK32
6S/VFVJT97nsTvLvgFUXU4LxNHHGfOqDSa8rEePs61P5Y5plalilw61XR8t2faQLWjMxfTRx7clJ
5SGPj7VM0ROo9878C7mFH1qHa0Nm3ZMl9Pe7q1653DwD8qKh6JubQp2ZEvstgzZ4eE7qc77bzzuj
XsS3Sx00CPERS4aa+nvTFIDuHEgi2tXXMcRE+IW6R+HTVMpjrX3yCNgZ4m9CpFTY81LOmXZWNBeD
txpXMOIl2/g+eNlRzWB+XwsDW+gIVOSEbsFZMykisjZvB3T4OYik8cP1aq233VEo+/7NpYnRCkYY
vg/cUqaHCQ8hV+QV/NLrpXgQwKFNdp+HQ0ya3Rlj9mySiPWO+FXcSfZbAFYtoMJRvKIJpvIaSjIj
/mVGMD9PgLugJyVgl9iq8piykLbbIjUYULVLJ5b9HGKUJRHy1bDx1C8puZFqWzY+ZQsL6DGwI6wf
zYkGbCPsqteEPryXTAr5vayBQSVeqa4KVpO3IYedNLqur3ylE4raAWbSWeZL6UJeIWBX3b/Bw/mQ
RVRtAMb/MzVeRmdkVOP+eYR3kcs+j8GbG793/tVJ+uDnargQPr+ekhu6MymkEpZBIv4eFYmk+cZQ
VvUHho1SHvIeFMlRN2yD6vh2qXpeDrfD8wuHR9sAeNNe5sIl3phR7JWjZrefKJedQA4vs8XgPgYa
vKbqUOM4JAysBw3ulWrK+LnOdXXWMPI0tD+BOfwrPKIhawui+bxydfkp0/+okHxlzplqaHC/HKGv
d758gLB+dycrJNtvs9NFu5+aLvj2fzl61wEvVrEhWzlv/MC80h7vim7arzITmmEDiEfnwyI618qs
gyGMHAvUtxH6j5QHO4HaLC8BrG1y7Nfl1z7r1cNrSSlqW0ztKbpl2F63JYd3ELvV0PFr/Ovr8sTc
9+Lc+Gedxxt0KlY9tgjpgqqarrsbb3FBdzpC0V3A5Yowq8E9Hiff6fp4uxi9IWl7YB5+BkncTaAw
gSvJmyQoJ7HyLLMWczQvppRz/UiDjEIkVqZ3Z0ObEpjbowmxE1JMq5oq62nwV9gOqtq+yCIkK3zr
I9BT57oIbmYcMmiGfFE1EZcRWv9R5j44wuIWCSgEOzqXorxJcKvcVfr6WkODvOyFMhWt0VI4YZ7A
TCo21k2GXoNtC1K0jsh4sWvRCQhCOigG28guJgixdEFXj0PVWBiNCfYGiPdZ4KLX8st+nKGNxOFw
2zm3YNCEHi5iP6R7RaYMgJW3ixrvhRfDQFIa/sPOF+uo0viBhNNYhWNUDZx9bhIlJJp833YWuZ9S
nheZlACFKNDIo8dycA/nVn/sULPFaqB1ST1ssID++EJI8REiqb+ykkwXEjC/7kryCAfNZ2lrpdx1
ov/D1IOfFKVGCB10fklAyE1lj1KyjNoM2eWE3P/vzEFmFu6bxFFzsqwV5yYxwlR3xWPUQVyOORs4
8uGTPTVQavnLreu06V6l/8oD4f1cMjmC/AqCm6vmvAeI0/6j9gDdj9zRNxeIeywYdd7hUonaimoe
FQeBR2FuJ8NPWMbySkkaxk8Lx3aPIwsYnwhuKEglbfUI6cvTj3omXMCg+PyOMLkydnv2nGuxPo6j
Ano0GHY+ufhelzyHkYRfH0IYmGAGbyTT2iqMxYbdydyUzKnpa1tezkFsYKlZvckNwxx7MHWFym0S
Gb+bj2naJEqzauHPJlCvgbjZ0NB4D8MjHgQTvlKOvQEdHutEvP00f7d260MueBXE4u0PwkmJAHh0
qRNMMRK8yds1Jl/gNsgZXJxZTBot7VF3NiFK+vhNU2np3ybHp7208/8EEVTDyTzoLK4s9cHT3CNf
iG6D6PPbLKhKok7PK84luNdzYh2bItX5v9JDHbQQlHZpv0UBGpcbmT3vhn0Ah96Jn6zwFs1aJeg9
jryVnpEA4/CFsl79LC6gjBoHUrnISKu18DEgx9j3I3R3b5vHMCG8aJ7eZkweYkzdr3Df5t4V+495
wN0QedXtOAMnHSAEidsJeP+Xmd2o+xQzYQEOqa3Lc7KMWhkiQ6sQJPsfHHKfMoMNfEsudYt55tIr
8+/JjzYLDPziv2AP8CRBhKeuyjIdiLQ0rk22YasVOkMCcv92fq7aRumcq2sso0cdjV+CdFASP1NI
laXiVB8zf5/liLvsfsSwaWhX+jkXs80xphfVBZWDW2pITf+J5IJc2OrD16ik1E3wTInfw855GqWD
fqQL73TVk4gjW1LVDyvAlaOqyfP8/DwJJAFiiNGG0rRgXM7euIwd2iDTNzBYUUq29uGj5fXhvB0V
HFzmZNX/fvPx7bR7pN0VjNpFT4pZfLkA7P+V7N2z4rx3WcqcXz0cxq0D7XJy7zWVFJ+5+zyS+Y80
mZBpPRvapRkgcQjRqYidVxjD2U6JxIBo0OW/veEZ9LOfPkvypY8VoWdvdsoMpRVmBr0mP2VEUi6G
kikWdxVMnM8KHwLNoSWxpJFYUVK0iEYzTjXZIAFPImnB8V6/4HcrI06CS7m2SvAP12ODHdyAMEo4
dMH21Ew/NyXt/BEfTp7ZhAz7T/gDPovU9YtLByLPRNKCJq2mG3qXES8H1Wqr5KD1OBf5TXI6Vp3x
xgZlM80nC+tRKeefHy/CDzNZtz0hq9CzxV4h1ywhC/NOWroqqWXLejP/5Mw8uAZz4WTRqyFD2xWV
Qgr1MuxGykfSMrFmdalxHcInEthqsf/xUkOSWdIMUVW7HTE0B8yXkl5zvs+2n7ubHpHjPBp4f6aK
6YB/JiayrbwJSgDGLFYKQaqD22/aZTLzfutQkivPlnA2N3S/XfqrzGN3Mz/NnUhTRnwGeOH6kZ88
JWd4Ankb182SsVcHFKZnnFM2/KRtwBiUnkjDPW2orZa37UnJQykiusid9HRwA5PicpmqO7ynm1C0
TBuNv7orRDe9iENfpdEifcNoAzHaQ0ptAJ6D1UVK4fsN+u332xZfETv+Nu9VWwwNBrMvUtnPb6Uw
sp8vv+gPEnTNkEwbBYgqhX0N4janZ+Mk18sepr3fxBFBBqaXWSbqbkUbkubcI/baN+Vum3jtUx6z
opBRm2D+NrMMdOkiY72ruprrf/sQH37VizxPKcEhlO75UPTHjLser3Ruac2/Uz11Y7lMYdt2c177
5BIxXFr1Rg5xmxs2Uu1odIOc5jydFpdlFsQqI8j9tqCnUx+3UWooeDXZGOM6mCweLmM6NDJrvO08
vt2LFH0FxtFwAphvj+iooX85nZu1doaiG0Kkxt0G9HOWEAZu5v+q69TQ/ly0vUuuPkxKcnlh85DW
7VBLAf6+inOto8YnKXur7jgFISCFPZSsEr8gbWxQL8jlbOhXsrry8d+u4KL3I2JrDswmwdjqXryR
2/BmkG3McaW+AK0tq4s6zYAEKR4DwRfYHRDygUN/NgpIyaaQyRCTReGIhuZfBzSkp3vNs52g7Oh1
q65O1cRmRNxhwqItB+hm9I4k3Rpk6Ui1m7VoqIjsUnQPu90SAdvW/ZbElKeQxkBBfrTynKWR5m7S
GdSh8xCylaKIm2J4IZxmRNq4XopnORfGSANak9/ac7HlStaYw0TqVZ2d3Eq3MZqG8Rzkgufo7NsD
8IaqS4GAGRFP4NGsOfS4MEOXoGuGfCq+KrmCDl7tRSe30lFblMmixJoVm9QPuiG0264aCOnrR93V
M6ofkcTblmGTELXoS/D6QXnX9AHQoXpl4VoUXC+T1IvQn9FwRL5p3OdZ4sfD1WH3HVpxvsF6EpJL
ydFpkU8McUipgJV2+Y7eKbqbXTCfpJZq9DX8JAEW5HQpUNXDlD3yyW85V+mFeDuKMak+NXiHfd95
ZQjhDGyD5mB9Z0yAeX9odQ7vD1s7i7YJiceW3Fxs7l0mALxgsC4AuVjPkkPVn9Wy6m0ivu2DNwkK
L4QwMc5pZ3fmJaz6RBL7MpI4uQ6aLVgaw0sQnZ9VXSxUutIp5b4YowPo7Znp9p2xTVIXqhEF/2vQ
oBz8VQkbaFOcSMFEg5N/W8n4zhhefPb5KZTrZpP34zY6T9pfzTgV0KrMTakBoXz++Qe18KoxA0HE
Pqpkfrl+PGm2KnwiiEKwuzvO661XEatl+1VGeEnCd1UtqZ2NianK4FdBy8LA+EDtAJTx3wGHyARK
fnAMgrBWYYk0TujeCmGtkhiRrK8R0MY40dAWdsQ1whufU/negzNpfeFRZ7+X+zIy2n0jbLS9pp84
UdG4Zt3BxzUClpdSPDwvfmhM9YzoiSpscBDYZvqTP+AEVMApsyZ90lNc5nB/OGC+N2x8KkBPjw3C
EAkNzKU1y2/EGzBwu5hypmxCSI4EhO9E96O4V00ArVmUqFNclTgBj+AuUMUidlyDsFpWnDCYw1Ut
nXGTopiC3ObL0jkiB5KyI5HDO5sguR1/GGSCVIK2fuhfT4SdQ3m5gfRs1i08UKBvUqiKPl1zybqK
j44d8W8dkzTZkN85c9AWaC3Ih9n6l0RrDpe99RgPshlP/moZELiBmbPQvgcYn9SO0QNe3RIm2AOk
xmTbdy1o3yjv4V+8n814RNi3ecv6We/f/wjHUUqeCXg3r+OxEUo65N0OEiBA5/v7Ji+k/WQVwJqg
qTLsJn2xpJBxpRhEGAJZfCsNo055G2Cc8c7uJPJTUW+xCK1+iwoJYAeYLGlmQvAgHMVJiRd74Myt
RgLCVmfvRussSsDC4d4v0/cLJ4IBMsVmmDPHeXzIUEjhoFdIuis+EKsWvgbfqZ/wh1zG7gFTekdV
S4ug7GotS/cCEGknkLxEmZCe6kwPOJNC1M7d6lukbfwPTG2/b53M1rYSwgCt9oFHNUhYgbG3Qgow
eCqSZtF/mmEJiVV6xPGJfAMCtC2IgelVKQAO0Cvy23G/C8UpB332PMQjlasj9bXJk1jyTaUMxALV
W4a4oHN9YnAmTcFzCxNSZRNBUwQUhr27bt1jSU9cBcZfeg6/ltA1m71gfrhP4cXA1VSTA22rvN6M
UzyNxa7BxypNqDJqWmYIQGUkYZCihdQOyr2z/a6+8oU4BKuneHhAGTnKUo1GUNHQCyWACB533Wel
Agw3KHVTAQ+Ui4vEBo5Wtc8n/nPPw0YQ8oyzgl1HWZDHjZubqKb7NdODeZ8PsYd+N1UYjpuiW+HY
apfCvi8bYN9ZQ+GSTge9TFmeWtKxFSWkQmBH+1VH1srx5/8Phf5D74k+4gEjBTAYaWw4QALjkghh
nixa9P+dj4ILd0z91w+3usKWsYrdzW95IVtXWdclfK7a0DcPsj7dyfTNJMiEdQ1JVbF2vWVMeZ2H
5+hCDnW0Q5GkAW7oupiq11WsRokADYp9BrApTtRP0RPLsfir8PlL4rKhY9EJWNXg5b2yCFwSEaSC
BJg4GCI1jV9egpLeExcIenlM0H/9jzDCIDLyur+OCi1/WcBVvLGJ5Md8Sm4Ys9LnegqYicmOAH78
8I78JcTNlVSkW9BJja0HDaB+NEt3KPx3XnWzNVKAFe5nTR+qZ0pbARfvDV9MC1QpDhU/E636/R1p
VcH6/0FK8HzYO7R3kvC4tuIT9xflHhyEcQFuOw0Eye8zJE4JQAres4JXWE0ayFQHVpFTkXkW9KQr
21m5HcIP4hG5dRuahb67InzmPuZ+mVPtfWDDU99rjLyB4YflA7EQTjQZCMLgdKocotFC0mBbmol5
wJlVk0VDKJSkLvZE67pIzlk5ywFror/7wv9dDUulA2IXWq74ZZe86FgwmvXYVU/e848aJUFWRBOW
OpXEC9mcd/6tV2NUHr+jxIGmJqR77+sTevgcTvU4cbM7T04cKlDqyTWt4yaRZGCzQiUcqvtvTL4/
y5U+nYIY0rgTfTbtjIDkIPHcd6QdLMwmefsl4ZjgSozP0x6CFj+9fTQkHis8Yd1TbFHB4zENToBk
/GXCQEUr2rrnzyDqpkwjN8n1sNoGRsseR2O4zAhXUjX5AnVHv9+2dCIOVQExih2UV4EXynVWiWwW
xLItfudOgc0usrZePC5gzTr0xrmoPTSCr11Xt83m6ZckaQpDiumYlnaA6aCheTtyz5IapX40Taw0
VdTS4FrspjwhyYJVQq87Ea/VZiMsXasG5m2utbohIZNA1el/4BLH/OAEPC8z7iNsGZ2oJtUL/l9U
3vgukQ7x94wqBf+LYAa41sevumySN849m+fZCuBct6OKpR5fpOYhd3yq13/vq8ZaUDQGwjtHENy/
PKgcvdplrSML3Ru7HwjBe8wRjqSz29em6XEY4YQr7Fkc3GnTT+sldivD2PgPAAZQlPxhL848gLoJ
z0g8+MBDbUM9jnnSBhbx+MIoOTPdrsLR3t9bkIUC0Oo+z0oiEim8aexJCc9UiXEpKlpMk3QPfVTq
mp0AEZM7BXjZjbCkDWE2dnz7j1dG4ULReIblQzxEMJh1X88oxgTjNvcQh35Br4GGW0KLEuAdt+/2
DyX4sqDXp22fwqHd3qAzkLiMD0TKTn6h8vHLBsb/nfYUXNfHOOVIYXgOMe8Gqm68Xd+WGSMVuoDk
y1ZEYOCergbwOSK2kIfMMbQuOE0Z6JTz1aR1l2LdfiAilUJoJltW3yXy+D74EZpahx/0PZyHi1ib
zvmJeryytlQLKZK2os2Mb4ToGs5uGmgrTgMmsGTgI/0/hXOU9upZd8C9SnXDnex+ukU+4zRWrzsi
IqVYPYRnLQm8xJWUs/qTnSFjAqGZilReG+sbaNNqPwJzoCYuYgAe3cD/TG55FID9CsHamY3M5gmZ
vLadU3wIpsLW2ywCCJkDJcRKZZLfkK3C0Ublmg4WyIZ7UWCMdx6pN2zcaozVSEcvr4Mkd4LR3xRt
/4jdTCkMLPNLPvr1vDr8roPP7DPGA1yCM8fJzhcqXlLv2Lb0gcfmpeqdA/nHrCzqFhls5LYkiqsc
Rbz7mKui+N1W6QHXweteEWkeE97kDkXNp5E2DMZ9zKNL4oAtQ6p58Nb2vGg7B9aPNX0ZLOc1c5Ts
XSws/d/YUv89pdFrPBRWRol+3e5re4mvJVboN/145K1pz8UVyJT5BPHzMmcIpqmTclp3AlHiAnRX
DyE00p9AFL1sT1Rx9OZqHRLpdvzRc8hTaMHEVk1iyTor69qNHFJVdIvly3CusQBLxb/ArAsco/Dm
XF5+EEBla4f6Rlsnxn4j7UUEINjJQCFwBXErSNcDI6portnVdV7nti8KC9b149mTXGxdN2n+IgNv
j9rFU4skISX18+ECy/oy++ET1SJGcJmEeOqbxomUBDGMWswJuPtkJGNY71Rh7cXPAS5Zbu15+A5g
bBHBAj/9ddHKjgPTGGWwwQtP5ZvRctsbuYBtFVZXWsuZoEbd+DBpV8ySIErh7x+jm1qizulpEZA3
R40DNnHLspCpxClEyPxaz5atkpLVrryiLMHd/nfHJ+QxVb9BaxBmIby/29JD7UJ+76rsLi7626O/
1psj0TLIMruXBjzCMqXs33Nk1WgptGLZFr478fjID7jhXy1BGgCmtRrfz1wz2A85KbWtFX1+GWhF
UFOoJZ/UJvW/8+ee9ms1JLCBnNAZ1RfjJ6O+CSgoDvAGbi4Cl+7b7hDKxyzWouwq6YyTF4PlEaoB
i0Z/Z73OReKPVgBHulq4PWLF9qe4QLD95K605IdAJCtBWb3eAy2jXuKQc4MU2U12+3JN3KVskLyy
suTY1H+ipWjfv2mzxyA1EipieMfEzufTh+HVP3gbpURzy4Wm7LXcoqP33rZbSCd8Aktv+22T1uIH
uwzy865Hrcmdx31XnWt+smfHsp+fBCv1YgV50TXL2ixwjXhNun85Y8k/FbnuytVs6R3hCj+fA2vk
yNw82j2igqbmBYSWV93x6aT0i+k9XpWTeUCfnIu1+5dwxhmVBSVMKFMbLWCJfQ3/PuaZUz86cYp0
E5lACHV68gIzHEvRze9mCiRR4c4LqI2kUyUw3k7FisORS/pAIFRbsfwIh4hY4Rhfqep3/W+C81Lf
KwzcSS/H9plqsyAUPFXhd7N4xXGTGBFarJe5uw87VwRn9z6bAkVBJTetRKhn589u7JRRJCTYKUik
KoTJNGXU/DvK+TzsdXhC/sBoHj1OYNCwJMQb7FydRAEYwOqk6Uw+g8irXdZrt2iIxW4Bqxgd3WoP
dVIhc7bkARbCzZfelhX5XjGqB5ONyPncWnmYr+MLH/luEUpiElus95JqsoAzUq6L1Y1ZLigY2xRX
ZEX2gHKN7BlxYAHAxT9n7zHiM7FAOrCx2eytqkXBOq2aU2+SFeXiY9YHF/+qJ1S4e0HzVfvI/XfM
Rq0viy9Pe91Y4ui3jmix2Uvo+0r0qpKtiisarB/NnaRIofRTJZOIJ+3Nnhd3dWeH6stzcT2sw/6i
5y7DoVHpS5A1F4qsqqVM3XEqAXVjr7YE/A81pXrLAwwldOwlq++010uRauC5Zpfuw4dtlVBRRtiz
PjmOopcU81pIE7DyZGUCEbZR+tUvguRUxzKCRuMaCingGicU4R4GXAjhf5z/UIVuQahLUZLBC+3W
YuPAHTT6qJtmZGmdaT+4B24O3sbtAKi/+PZqsWKgkbUENRgVoXM/bqWXB59jd+SlRbp5MNQtvJAo
NxRAPCarKnJPilosbSIp1+CoW/jtT8u0et3mBxhhQ9lj21g4HzYG0dU9DjwtrvWRLT1oxMTOuOCn
b+wZFhBoee/hXEQoWq4b2D4CKzW16lUy8FDrSqypE11SdaBUqW98x+zhRvGHrd4p7Me7MhxFg++W
3mrwSui5x4Z3/wA5QenkeANuR19s69Htx/PO95+Tc4tMBz91jELR1n4pwW/lCr49hz9xM62p/ZVD
L5fU6RaC8UF63I1AMz1IYoVhoRIHi1cVfZLCg82hQ/sUxt+z1Hxem9lsztQScwhaaVKZMB7N0t9d
z7YNdXp4dl7VfMbkJR9US67YkkCBf+siIX6pv4pm8P6HxX1N+vpgA5RdRvbhNaGuypwQYP6ZWj+A
QwHrraCwG2+SNfoI+iCrckpEeYxpvGOE5+sD0YCivQv8txP5BgCLIFlaeobNk3+w7McPjgNe4Y2F
L2YM96SFEZ7v9VtVzvzW4SF49sQV0KUo01D/rTyq8ZuckGxUwCvuNKxUav2VTaRNQv0lyAr99asB
+Xbwg4tAr6/JimeIep0GUFFy7LE0VgNSkH/ST/BWrdH6hpUgq4FjwoURSrG/rlfalBZswobqcuqM
vwwVFu+tc4/xXtGQJ5R/fRLV0q/nDdxqXAmpoeOIVzEofB6k4m8GQs2HDB8FygXkGIi/+dq8S7Ts
cd68Oc3gPhg7zaxlTKaF8fH98+ngYdnOQbNj0u+l0Y1/ovZ+3HDAphDtC38gHBmuGCEsbiuVFnPZ
Kn8rJKZ6rqHn3iae6YLnUHRnWj+i4t2cMwdqD5gZo55Q+ShrgNPi1VjZi0rDqav3yVUBGLirwKD5
S+Q4/06IAJ7gx10VX7hIcaZ7uwQdPr2YKfCH7aiR4Xpq8DW9bfx6MqX3s14rlqS8D1HvCYN6ltro
GK3zKQLX0YnHGblM2+bTLKsQwzyeY+0K6YKILYvu9Np70zVY6FwSIR8wb+KGIQD6qBMUCnoFgnDX
k6roBjONoBd+5LmQQ7cnMJ6sKMrHP1bEs7IHGHoywPgnFRvnQYAZrT2DhOGao38+TPU7QDJcEVAT
mTvKMo2ON61q68BR1a2Z/rygpPW0x8t36qiSfv6Id/dMu+2BRme3RB6mxelUCxGLsLn9WWspVY/y
9bFnegTwMU//jQ7Ez+I6HwN38XDQRCiMSyuZ6r9FUkRHuBTI3ckvaPOfrVNkmkB6VS8OIbrB3UpM
XuAGDTWbdnmTP6y7NxlUxrpYVY6bqw5Gooo5iaax2xHmBc/MNxOQ5nvwGJPbvm6Gta8sxbFFLk/+
QqmX9mv0cuzzrEqRptoYB0kW7VLVPoX3AdJqUunJEqwBkjyVhVax0hqFWASFX4gv8s30Mhv+XVvD
Yk6tUnCT5sZiYS5gzQYNlTItITWknKDa9BMzvYjV7gKGIqrg4qg8rNMWg2VXAg9OqaHJ1gB2IJ2P
ihrBQwQxZ01Lv1TCEIXPJ3XNeakx41Br9krKJ9hVgcFF2UKzMcl5CRbkQ4oCqpZLRI2z7BLL8mZB
YBnEVvB2N5BueewYOt/KMe3bsCVJpSm9hqB/B9ppRFQ6mbkVLhLKIgGlyWCfVb4NGgBobG7jL6wK
0BMrjpLVgwf6nWSy907fSyqwCpz2tJrgSWSLSHnmWS8mJrAfR6wjcR16H+K5xexephcjils9LGWI
Mo7Oohydnj+iRC8VIUQmQPFcbNSH7d245FBD1rDd9R5JIlinJSBOxWHprn3pvJdXe0oIq3/gbHqu
9IJgygZxOQw0JGmSuInr6HtnepNJIviJ7k4BAKtbwOZEmOPnwMXJdpIQFzZizmD3bTijINodpT2D
ctq5c3avwBFxKoLufq/YTOC+kF0091bngS+qhvK/djCxWrZ7IGdXdcheMU/NRoBjWVxtb650swb9
1Kj3seY10ziiWY26zlbAaGGOrlqXMF1kb6Nh28EPUCngWo+N9tPUjF94T4XtBitwUQIu1kVjbOba
MUOoF6YlV2/8ar1rFIpGf7vFiAg057I7pJHgzfl90d0ZGpVHTlEi7puqQHMz0UWYWSVXtjLSUFGK
GD5EZBCPx0t3M+CblTsssVzKsoUzsy3eu7ytGZ3vJtXaQsUwEMKwheRTFwBr1UTQnkRJmT5DfQ2q
gIZzJcsLm6On/6XZR+klrHldJGOFCOHXZdv4WYdnv7IBZoEnNuynG1YmHztvHv6M2GrbfjunePT/
9LdPg9HOQBzT3RauxjJ/vjvfUcN1INbbvO8ngCbAGW2umy2IfeZYElTBdbXl++UaaF6JkWAe5Mgi
yEbVjk6TT68nhl8J+PzqkpXbFJ/BV2Jz60iuaJRw+R49eBc9MAjtjPiuxtEvvPekIQ50RX4MAedK
ybsYuu3x5iGyPf2c0OQyT/dT5Trg2JGya099nXCLiXN8DnuyJEWeUR5O1AP183JJAj6IPs7gRerV
XazrKImN5wUa+E2IdRG4axoB0+Vw/g2vmymrBKJz0BYgWaUcix6bafZGz04336ErZ4+Y4yHmMGJl
2s88QfsewxXV9+hVLma+lXQNNBl465sQz4WHL+PK4GJudfbHRHw7Kav3ZyIo1GYV9/Fz4Qbb5mJo
VDqjpuo3jWB+2kZuC0Rie50sDPkKF4ARDT8VPzle553D2xe0ZquZMKl2DwfauUsbhO7VGEOQbtvV
hgexW6MEK0ZnWozxmojGlITx4SqjM2ieC8G4Tne1mc6Zi6bDWidDxPa5LksLBUTZmfAj3bFbuVT/
gs5IF1PRxWCJR8nfkWjjLRwA9VYQGH30OaNit5d1E+9EKwv4v9oQRAL/q4fqhAj8zFH1Eqlo4FWA
2XtrePFhpjYyLBBDtbzni/YYoeyPiC/8TdIlYNJcXLaz0P9DQaar4kIPsIexrY/HPYwpx/QR9X4G
j9VMm+/WTUda8B273tWZ7ABzGDdWQBb8vdvoPg5J6EF2LtGTrvzHlgeXL8YvGlBMOoSX+m59p+BW
edLk/3BjEW2PKivmtf/pD+jI+lJCF8FiKx9HIk+hK8Gzs3KFQVO1KbhnaSwWSJWzfxFFU3Zh7BUg
2Q890keorPJ56DjBita7uHL9MK2eLBgZ7yNSgR3VuoliW12F+6AsKwv9PRuZBV7Zz2eKxeLl6ozc
PbBljGBMiAhEDp2Nap9MR+/B3kf0VXeHXZil/ZFCeZtkLgi5rjum6KgoqkgpUajOHKwxAIrwyOUr
e7DV05cbViv662Ck/HFpBuO1dcVIWI6X9e+kBICca4MUUEzUjczYCJZY32RX9mu/gzBoGlVC5XR1
HXixcPEk1vl+Evh9bneZtej3oPnTR8GndFLmOVpqW6zDg/Q/+bgVb7Nrt+N4m3vl0T7hblR9IZW9
vXTKGpcWVolAnXzqIroMpMkelkDtN1agFYguszIp1EoPVBPGT1M2IWS3Hpppf/scZki0B+3BDs1Y
VgGoB8GA54pojOj3FbXZy3P2zhufGV4DZ3/oMGlX0knXqbx+ae1IKGhr0guNaA2ABcyylnQdMsSP
m3DjsCc/xVZy0cfuruFjoPgYd1EROwWde0HMpyeHpKLYV3oQfC7bnpkbFYcO7YHfy33EcSR1dvQl
IFOFKJBkMBcMLIbJ/tP01YAABNXfEHGu+QLFvn5pDFYyP2wMx5Zw7cWFJ7KnkBRzoatpA/JGdYW6
zs7mRmL98VzWOfswaEiwSK6rlCnZjSGbsYzlLqZpyWiYBLYwbJxDWtUj3+55GevtHzh6m4T1Xy4r
remhYjNVraxR4dFkP4LDjFhTkIaYFb16CbL1FQhQjMxvqnIKdbVxoPBcEUNvqTazfzdz1YVJSFps
qzWfDbUgBi7vWz+kqIGnDaTqUhOu9p4IPJ1P5hGhueUcAaCBvaKRtJAAQimOndVti8KGrgF5QayY
LpPsEpq2zUGZfk0Ew1JiSgHTSI6rbUmn9Tv2LmoJ+2h0KFEvFOOpFlsYIR1uSIk93m3URSZPNW3N
jR89gTDbxpa2l0e5XNbR8dEAAgr6Vy3SCKwmMf3d5ZRWAiAmIwCntSDwnPJC+V2Z5OL5JgHvWbbI
zpTZTvHSVE5BCI9jxS2xwr+Ygwm9Pxzf+T1mzDORHWQxCVuebUSyDt5v1oDD+zmSkZasNHW6I4z2
3Aw0MqW/zQV4ClNIEuCqoAco4us4OmZL4egwD5dQ3G1bNAPk/38inDl8k8wa9yn1INEZyM2xAREI
hql5EwVxY6ZlcrsCE4Z4y+BrXG7JzXQlotF5fW9UDQbeI9kbmUSWyp7NyuRzIc1vXgsvofyQ2JeL
wmP7D5J16fiasNqhlDlxAZGIXQHzKubFiFhjEZcJn/8Pk2QZEDpUnjB7vNUzv5XQu49ecRf8dNeS
5xWrLri1pTjMAr/A7ZW1oUZ32o2o4zeac72gLroSnszIr8gREoEwHh6sHDZ0/1pp36R80Yw/arOr
+HQYmMrtrwO3T7sc4iFlYf0RmhyGjyJemPeekb4zEcQfakdako8IYI8nrPNy+Nl6K2JJwSk4P1pl
2dDpiUKywCLw4w7n7cr352TCBXn6CZzTeFSlFpMGJS/8sjmtUkmwWK6/W0xsqQjbQWHJMA3WtcIn
55e9wXefnV1r08WQjrhHiH+YjEwRI4gL6qG4xb1SfI97P3QEm0hoqetIdJCFnW35PYFFo+9ObjEY
D18Us3AutRjuhJhL3K/VVz2Syc90Huef3vxT9pUlaz+m9gh/S2RBaaosvN1lEa69J34tObROuQ8N
T4NbS41zvz8uJFQfmYNDXi/hgLy4oJmxTvLJ60thJMpzXkBj0vBDaxGI0l3UczU430lwAeyJfE3N
m/jXArU4E1JXyoB+V2tluP7h7Not1/4iHQx+UXCA3Htw9SFowxq1STs8r8I5QSWQcyYMjvOusjCV
ULwnPHfQO0v63aHqQDnXdLcdna4qt15NbfH9V3T5ZI6QYMZeGhZmuGK8k96gifs3nVFdmpOmmfo8
ICh8oMgUCjqYtDymxIeUFGYDuKD2Nr9bPH2Z2fdV3OY/Pr9kpcFzoFMUhds6Pj4cFSXJNL1LjFyp
M3IQGSdFu5EMMp3EZ3uLQMhfdXAtQvi/KCeeY3l9NR2dYZxj30GU5J81UsdXSvZMwOv+p1JpZGhI
wGj3v4izhBTSmtcNb+fbWT/X+9mB9HB75OcjsyZ73XR95Rl3xKHu/CUsfcRKXSDAj/MGx2CLM5t5
asU/V/cP9nezQVugILaF4TtSvVZfU0KFyKY9UH5Qe1adurpdnO0k2Dw3iVmc+Gp/BAaeEm6J0Jtl
epXK3ygC+klTzQRUq91hEI6SiLzbWkTn48olNhLEsdbT9HGvS/8yLzpIih1HcMBOrNHbtkP9zIzx
0dvjdsRZhvXU1o09cveo5mGJdbbNI7/5bin0ruJmHRgLegKSWzL3y0sPq0EZxxC0zec7/YOPdh7z
rO694WeWQa4CVfNTpMEX+IoIM+cpRVDY+laGuPcXHoOgu/1yepubRZXwrSl2/bMSR8sZT4AS2hEX
bsxbJP6nLc+wwarpXUVk4ZoLtZ2i0F90Wf1hKAFGVNtMSP/6juC504zoDlWraYRQNY2EYHJQwAOR
04hSjj1bd5rcX+Zd+1itXisPguxYi+Tc/IiqbDj4Qoet4HGsPJTiYagMvCYDYL59nStnhaUepUsh
7dYi6A7kXpm4Ix168CmiuzuVPiB7JkupVbOZPRpMg0mb+u342T5jrEC9ERpKQ2fvTUonupXS5i+p
MTwGZ7ff8KIMjT+hgBUOWpEMiyxBIw3N7kBc8y/gWVj1gnewvYgzUtsszychxUnuzTm3TRm3EJQ2
cdm9OWKs2AN+E3SgmcbBP4HENgR5TMgmkA+qBHoWabuisz29tLwGx065a7w+CKktSEXce4QIBl6W
eGTSGX8ZpqmI78iFelzNz4EnyXd5kcqBKuTT72ci+CK41TaY9whE8bcWrfLimqF1Kqov0vQ/nQBm
SS2vkHC5E3GIyRyvV9MOQcvuUjd0giiW28CMh16Z2a+Dwtgg8wtL43j4KiItSh2woKchxAsTiz9z
ZA4BApjy4DOzMZOSxdJ8G51GO+H99lnJ14c47MT9v6hjg8leRYHM9IwedIXC0ygDl60RGOfLfNe9
QCpLc50W95IRQ+YQEqtqQlWNiPhXRg03RsMo1Gd9DmDRC20JpUhyO8ayXQ2s3ANXXuEYXxfiEX8u
3MfJEcfcUJKpdX2UrlUo7rPHEgFQRvGXQJmFI4o80XNk3H0dLyaURyoMuA9HKd4Dplcvvo/K+KQp
am/gvffKObUhgMono+TvgxnY2ziY6MgWCW4oaLDWU7Tmez3dHZmeK3q0X7P6jxgt0DGwsbhiEqnI
E8+FPg4KEcgiTufPPkCa75nv2vFVLIDWkeQUFrSwFsB0hCjc3MX6Xg2Vcywjz2Dh612fkH0nx3Bz
E9/EPRt1lNu7fNbJzl4PzDS1fE31k9tqxtVkV5+6biAHeQi7JWv4euiRVuWMGuutWsbyzSqFhytB
HohlQqoUjMt4YQo9B1sD2dTPxhg4OeanE0Q5eD03WQ0bCcyeH/blR1j3SC8fqtKTxBDFQM6L+uL0
kkA7rEJPO1HJbOOz0/OSuL207ChJwilKelVBlq3XGFvIdcKTf5E+BecFS6suFKK6mvjkmyfiU1mi
Nhi/10m/o+eoQ+eRJeFvJmFlK4e6qtxVfC7SP8+37Y4dnR3LRBOd4zJafU4SjTFalS4CmgpM2cVU
qQnk+qBh5lggDuKdSNx7pBnLFuaIhGmhIZaHjgu7vMe/3FL2uRC1IiowTq/2v+jRQnBymN9ji2pf
u6wUQ0d3UkzUddZgmggh2weQqn5346ALb+POFIQOgI74QJg8yszvj42bcv2ydVfBk+vLbZX138as
0NGZ17N8y6utdNMgw5uU8YVNjcsPlWdVBDSNGNhLIxcEWOnCsUFs0GbfeMPmNRSk9JbilH+WGKNW
7tvzZNVXVl4LV/WBJasI5gin0s27ptyogf7RvflcfKk0l9P2/NXa8h7GuB3jurOvrG7i9dW1Dylp
e8gSufT6s1vdGPEAELPurtU0z/SFVZp48IXJqUZqDjjTR5ZWcAocsezSaA7yk1ZjW3tqCXilJYtZ
IydHP1cpAfXLtLsiJWwQGyOajGuynl0Fd8rL08dY1ls/csAxVqUijfdF6DvYpZdqq3UWzAnH4Bpu
U6CLbHYpDBYSLyl5e2h0uFpF66CfAbFf0X0/PJD0qQJAlh/OCoKJvURIe5HbLr3VQj1nM7bWCpCo
eFzZD/Ae5tMRFO2HplGD9CcW62IPcGfsEEnFPojk7v5/vWeoS7SC/kBKsaSKsHdX5/UHPqx6/GrY
yyX+ORRFS9TdVglPfpvDk3XgSqAxOuuznVkQ/cVYXdIoa25i2wGPEG80Diza+jd5IAS6qkLrwZ/X
xE1kHt6AGBGMcsWM3ga6bck3RvxkFB9iLWkxTQ+EvsykVOE0BJhQeQhrT5F3si8ZFlZcdvR35ltk
FjOAIG3lJDagFCGya1/n6EwFcxeUi1O9Jpf/Dry6v4e+qEuho/rV1a8u6tVfDk8khGM2ggGud8kE
5MoJq91SidRjlnc0zj78XFbotQBUmEqT+FsWom/hFVvsEVqR8xfcSzqP8XJ0oCI4o9rQZqNfQmRz
b/lMD0XgXwrLSysntB5g3eJ6AEOiOgZWWtUFMdDS4zgYfH6KaFMt+eksHuNb/zrqBGA8Aeckaseq
LiQCcbaQzTjm8K53P4EGZJEvvvBB3d/oXviyZ28bfEyJWEtBwe2yZ8crTHgii27VElGTKWh2kn5x
LDfNMHL5TIa+s8tRnYqwnzulucCb2Q4kxX/tdISk2q5SFQ8evcHldTp2TWRwwvFZ8T8PebZw9AH+
RZwpJhHSOjJhkErh+cYzNB3ZhUHxUgDAIhs+h/E01K76rkKgj4jR7LfrMBskzf6Iuvc7dmjq6wlZ
J8zlCj3J4/Yz57rS94QhFGs5HEnXS/XLPhOQsPZt5HdS1nbrKGWhKdURPJfi0qr64J6TXyVLgv2B
594CNavVTmQwW1ij0Ekj7euIiWC8Qww/7r8Y4O0/3uje/DpypGprRDvFmOucXEShr9CNhVkKbaBu
jNWUOvSE19obvJEqbBdbUrffZeSH5tSliTGstAL7iR5xKWcPuwTrz6mdaDs91zx2BTvyRBlGnR9j
XBP3FlUsFx3NazWf+A/p7MRJYssq+q244+7xxY1TjpuMCUvIWpShTyazDcMKZNERN+jltxk4VqKo
dte/qkuXLl+lGjt0FrwG5J0NyZoiDBb7NUYHtQq/KnoV+OA3wfE1pyrxO3oxb/DdhN/LfWsbgRwa
wugUuvq8ikOMpmqwKC61Tcg0qg1+m2JsFgs2Tr2a3lmg+Rvj2H2JRRarex2G2ElR2c9XaqGqURZr
O/m+P3qsJ/jaX4qem18cbDrq9kfN00GhTyLkRIL3GnvzE1u2k0SIjsRjCxO/B9My+hIq68nMGndT
DjlTab1/80imI9uheBVD7UYFtsn2WsghofoChJVjpx2RiW20QbAUcg3U4CO26Hz+ZhZtKOKIRsQw
14me6fTpLAyMKPNJzg2OQZj8jP+lzS0E3Hi5q59j7IoAHjINgd0SzxMbOQRfBg/mGtSzK5ommkPQ
gu9368ofjOTiorcCEM5gDxbrLjLT2q4GRsQcpBPmxnq8jjLwY25Qi70nzdXIn8D9aCnCwYWK2iLv
vWqb1J4F2Di+GNNct9Ew0EmGTJpwYQSJT4qLiGulZ4Queun6f4s5Hdw1HqJpGc0THPwBNTEvF30a
A7gn6Orkq1dIzjgkJzH4lY9ypTs163CHunkovZuiWsLberAev1IT8n8ymEGyMvsZFkPtnEN5SMcr
ISfGHwtUDprzP9LXKBirTE5TsX8QARsAcVRwldpB/TEXxj8MH/Ly57gedUXT9DNinL+LQ2MzPFj6
3tltAVPiI7WCiIyIzGc0BxbO5SjTGqkTHRG5VOix5iL8ZaqwtbVL5q7g6/XEFWiK7Dv4NpJc7Np3
37AxJdlGKp0rF9uNgDHAjk09eXM981YQu4h20tdR/ZDEhL9b+d0bpu4fVcXSNakHXpfknUG3YSPL
liMAqynaLC/ilFM+ADMLYb3Z1mrdz2PcrXmH0tDGtqjdQ3NcoJH2MoSVhlYLspUhnJoYvaND1TPj
SIh3kNN6Rlm9jGvWhbD7cDp3lALWuzwz+NgI5+qgB9IHeJ+29rIePBZdpxOXhWWVp2sL0f3/RTML
8hERO0GRiHzvABAAQ51gP+fEnjjDMxypAzGLcTQzXUTRRCS2CmeCptpU8yd/cFIU6j/CgDfB9RLE
yVW8HtBZEB6C6LzGvx2MDJgye7pNg16437E0hXvhdxFyOgfti6WTueX8NhC4UnjPJMeM2/egp2zp
4BeT0JrvqsqYbZonYlTQFTjph6LTKmS04PlozHM2hzNBXy5IzE8dQInAslndxsB/fvC0ymoJw2lQ
C+7rz5ET1vZQvvvtAe0+cPrAkhBsJfuJ7GAH792TrFXadNZtpcnLNDZ0J+PvTuOu7oj4jL+DDbdy
nMy5aD7IWrvo84Cky8SRjOyFN2jQnkVDxqPk+6bOfn7ArQX0WDGylIuKRysxq33kjNObUupCFmMl
VlRISKVA855d1WKaTvdBzamXR4iSR8/itC7AjvJAjjBJjz8eFeQNOAkWbkTCPARcHC6/FgMdIwPk
I3rvGhzzNXI8OnLfquxg19PANYCMZZyKSM+xfPkAweb+tDCLGUVqzwmQdBwBmabBJMRa937jCsQ2
9F0qZs8L/KtP4lBBbwGPhS9XM7qii9ffy9FuFuk+gxP/MI9IoHIMbCldss0kHAPlFNjGllrQ8BQV
+EAUoN0zD0Ev4Xnhe5pMzPngCB+oL/4ImAENDSlc9hN8pk+I3Uu89KUcZw/OZaHtIOoM8EXLtE5F
9GhmYo7ka+pQL5wC7iHMgVNvdt+7G10nUaZhuFCFFOTm9FTVyjHe55OXnv54xx7C6mTuLS7VEU4g
4AYBbOdVFcwf2cDobJgT7B/iGx85Wv7OgJnhJ5VtN5KepnyCUNAYk1ni413ZoM70fvyP/grVkG0F
YBEBM1Hf0ywpXpHHK1Dha5ibxOI5XMO6pb+apIC+euLXckXbaPCZlKQDanhQu2PIUW0LvL7Td4AR
r/yyFas+FcHApD3H0EfyaLkzcDrkiCifQkKaC+Uz1XXZRqIvQ5sLzeLd+MGZKOkk/q9Aq48TRPXx
auxFLZVQtC8VB+DxY3ryBVjBjvKgjrzM/TwOveEMnTditpF+D8/3LGPAo/4z4kkfa20m5xpXfA6u
EE0jmNoS17BSlths/S+GMXJ4jk2AU7UffM02K8pSdBR/YjAuRBf3GxERHAn0uQhXny6dfL8gWLVq
f8gruVdxCuOOncgsphDqhLXXVnHCLl/+EzGq3tWmSaAAPLoSY956yGSbKYfrZbIBxW7wOetWnLF3
bPMoSwNlFbrG5ToP+z2Ih1OFEF+x3dMmtqUTxlct0pwjRmZSk/ENS4MXYbfoTIQz9frSFIV2W+s7
Qjss2K3Zd6J4P3/vP4Ixeotn9JqHtx7fiISyy8Rl5CyreuBw7MqIlLphsiv+KdFoV0mVHcsCbcrr
h3GY5qQr9CbW2MDKphY+z4zOvkvQMRP2Aw7UiJrcT8++7I9MGytrmTNUcfFgHFntOKJJBxb1Brob
hOC6VXqtD5tBKw/rMdpasTzI8INc6waa6k51pKWoHlu/qrtmOkzt5U3CQSbTjWVbxCvlZswCqDha
n4TYuk9ezHvkqDJgdr2ichTEZ8CZGyxiN/i30NKoeACxqwW94YprNHcnINCqA7grd7saYxN6i4fV
FHAUQ99+UxFx9MinonvZdRrSb1HkPxLWMtenh6b07mYshVBcAcqv3UCUTaxLaoxsLeJWgShi38rv
KdxFblHqWN9CqI2s0NhgRQM5OKeghIv4pAPBCRv1DsA/v854F4HHee6RJ7ZlYj33Mk7wwG+qgLXS
Kc7ehF+ErA2PMHAB1ETZMoNXQ/dbYAhMbo5xYtilleA9oSkjSQCukmYseLbZg/Y5bnGWjWz4NacP
l5p38/Rywz8FT2QSVoMIBZEJWvRFbNivRWvE+AWJI+scDxmllbVttfL5LXH+67u23FGsNhcVY1gs
XBVx/7QZyo7WlNkYyZd44IS/4vNFk0Q7RqIj+JGgFjxHTCXhq2ABIr4FibrNRV+GGkGXKljb7+Ig
wE49ZALBdNB4m4XGeJARHXq9oLl1b7BqM9VqlAvmCkkYlklx5vzx1N41c8vXMZd/U28GcCQBUkoM
WAEjrhZrfFzu6FNOZiINSeQaMAKifIPo/OA+R2ReMM7GYVm0LeYXXl8zBf8FKwJOcJab9vjhT6v6
MJo8gyV9bb8l9hXH8gsYHoyELByJco3iPLQD+YrckldiT+x6Es2Q8FV4xaX44dlKvVdhs+IOo126
wpWURSdH9viCwg5cT92Cc7M7sG7FoBRf/iootnmhfMD6yHmUwWx4azuPGpXM7P3B+mKiyEgbA/Mf
6TpD0Rkii9P6XC8RQJkjgkgZUjf3Frm8G9I/EOSdnBopKl3e+KIWwUHx3mULFmrTRK1XFlvqqjVN
jDxvVrv7AJB4yHmIrhVVDBlkfel6Zp6/faNFinsvNeCKfsvMvoccldnClX5kigOqRnc2A3DPHiTy
tNEI+6aREZV3ROlwyU8PMzoYRM37Q2B6Krb5DeGyto6pZcDnV1ShrFV48o3tkgGosRLU1UfH/t/v
qPsRy/1QjCUaQAs3vroW2fjvaNqGIU5wVj2MMNam6cU8xy0mWeqjxqMusc2N80k6xnmOigWFwWWy
Q8D3fRbyPffRkVFzJpyWvw97/SXk/np/qmhrnU60Z4rP+Qy7avkKsGNGzeAJDjsVtw718pOWKAa7
LqRAMJMSu5aHpM7I5ecH8W7TaUMsyGa3Nc/4dISPBqwiMv1q5bWiXScmxWItqGziatcTauNYQjz4
NOukEt3eN2nLIytzak/5pffrYW9eo6DexbGrrbJgcN364rHFsdrv9K7wTsrk31b2QnTQ4LSFdSuC
6CNbBj6qbSV5VlrVI26xsJgBJ7Tq4kZ3QdvbFEpm+PGEqR5rw6A6ZeLhW6Q3wxe3zdclGEqoXfiS
MJ5jKYdf9b/+puXZ+lKVW0nHWt7F7HLnzdtC7x7mAIGrGKTiie4gZPgbXPUQQtgh3M/xFtIzLGPH
1HZ6zoRkLolcYhKW4XX56Tc24xIq0k3HnccX7wPTM8qeBo+HtsArpsC5nuOHd14E46UZb8W2fFsv
Vn0NsKRdJVt7lhGrUm2VdIxgQbZIF/yr3ol8oNio3vbE/cK6xkrhDcPe/FwB3iktrZhAi1jW925e
TO53ht2JPMl0UTvubS2eGE8v2wxUiDFnsUfxmBLlPMWn9QShHetqiywWIHFWnkNiFB5/qXwF5mW3
ZRgYHO1vW79BYpN+IVlDgoTxpo++XH6oWiiUsyURzDKIMejnf/5VXFg+FIkdUMCNJb7G0OMhRe4y
jmjR0r+PrqHg+Opnqi6319uh5TX2APtTWoZT1xU+Ds4TN4uR6XRYA8S2+NdbT8I7n8B/XXUFQGrD
29/OfZ2tAb7zTilkG4Bje85/t6b9aoR18xM6Cbb8iVVp1mOYN37WZTxvqPDBDuU+FdXBlVV8m3Cy
hQJFw9o/a5PYZYRV9fjJYCQvbQp9OKCQ5WyPm4hdE4K/tbMaF6EL6KsZChleZLJauGr+OmJuf3ea
Y2t4IYv3/xGCds9P5RHSOlZeHI0B/wqdwxAzDFX/pK3/ADZT34eHxQAxxJPYH1sahSzWwBIZNyRi
S31SF4AN+uZJpsYHcJAAuYHeVhxk+Zh8aV8MunVbtTQNeq9Mvl3lHSWK/wuD+DxDE0gWaQKXDS3O
tnYVJyyGcgfQ4+g/ElqppA1n+8JZxK6NhzhOfc6T0WuuxOd9mUYz3XFEmJZ2XXFBpYyLuXL9aMiY
mIr03ox4tLDcZ6NlCAhx8lJuFqjePnc4OQj6V59rP6labSnWtCW8hgkF7avnLXKdyhmcRySnApDf
gxCjQnUbbWqfGgeFBhbxCQ/7WhH3bBOEE5HjNPSm5NX8vAQywMsmB6UMp2U7uR3nq3yHVfZZohKZ
VpuJrREt9LfapuwCfpjAUtVBgA5boSx1E32Xk25Uvu6g9LEfkP9fYTCW4gbkrDsZROI4cYwb77VW
tNLycskUFLS5BXHYuoGkECkeqj+uu22YgbFCQI8P0PYnBriSiqR4BnBN1aAQr0cLZI9Wc+IOJFVH
HZT+bF1QNu5xFofIDMAJ7ZI1xAHykIKQqQmYUl1ESL7I/CXD6EChT44CvFM3TYObhcXid3CXsL85
ikdZUsa9r9ddmDNtmRBNy9zp7z7lL+/+a5LbxK+G4sQbN7NVf/SdJe2HcQM2ao7XO23bQqSI+jLR
Y+0wNY4gD36xSKDtwkwqOZ4Qnq2WVjZYiOeS8DQHMALnq+enDTYg2V3/sXaGCMGLmWva/FUWzhgG
lns+izsxUSBwQifdj7UvnBTSlrhsym9yAuX0YSq2c9QTVwYyJ6PuLpz1fB/DYqEzgICdPCx7vSAk
8RACFrEq897OKujSWlheLT24hgpttdMC9jVyy0IMKn6uXQTEupsPJMEcT3YXip3df2VX0lwxSYaI
DOEwCtygSFPAQpDgflEp7xfhhT4cioluaZPXaL7kBjuqHBbg09a3N3zVfLGZFLlBvEaENSj8+1Jk
GXnYOHif8UCWQP6uDtl/BA08cJLzLE45u0mqJDRSynaFRc/w/IxiWR3yC8zsD0WqnR04jR4ZzQ6n
wGBFa6vGvZZBWRrqptV1lSXV9BylSwG+PksChThVMM1sP3UT0rrGlGl0cWq2aLCNpgO3E6aZMhUZ
bHcXTq5bqkhoWHaPzULM/0nGOmyLuch8DKP8uIYCEBucwe6y6+068XrjEvIlNbaWg30RYhur5ZdK
bPGhyB7sI1xQaN62KFrnP2IIhAQXjDCduVPNkuM1dXNFe1S0EL+Z+9iVV90xtWybwOeq5hax3OuH
0fiAAEdJDUxwOi73chMaeKFZksdTNuueAgIPQbotCB2iilmmJ86ty+iHn8bbCyYD+4UMD0phDr3b
fDDDifMFj0KfXlnjjPnlbJ6vs7O2cUDRNuEYv/ixlIQ3DDSjlIB8TarK/8MCQwBprdNputn1u01L
lyUhzzBihn9SS4HFmYV0IsD98JNLyedYLQUpICNBOPah8eSGw3n3kF5RFikcm2OriS9V7kZZtm8x
8OxhKSJwJRs8XNZMgq+1O8gp0zqdhKKCvO5un6lCLXziNpg4ld4EZaOJMbzjamcTeqnbkd55sCV4
VOch3MuvVlWchscjGzneHzaB+1nlNuqOZqzkfcJprd8/aPBXIOqM5F78/fzPHwA1q3EkLcmedl4a
+6Ot/qnIZ0srkZp3BbW5tb61F3rsCoC+pFZt5Ulrh7LTRZF1kj46JoeDG0oE9DR/wgxUvF+oulxq
a1EWlEPE6rInu/JqLXPo8uCzbogL9Ga4lZ1RSAfkL4JxbOf1uNpSKxvouWntngpuJr5sMR2VUWap
/hrBiVOF6k64AlhWj+dwdoZXArd8nrbjUNOGor7/ve7NzR/oJ8sMKaa22lCkKiKRs2eEHTVX8CQT
KQWNzNFJPzkuAhWwJ5lmQK7lbXpoT5PBmmZAPU4lVP5LNRhmuomcuzvvVr5jYqaIaQ8UnSCN4GxV
/35ol9/5NuPRiD5xBkxbjXgQsc3rnCDBeNC+i/xzsGUWRbrC973vB2f9o69GyfcEdeuGpdbAwxfb
fxoxMACAoq3jWbmXEhAHF7LhSjzoYWx4cBhZ5yPHzEG24dm96l+gtYxayxX73W/gwjeVmL0G/YKt
34E+hhiD1Pl2uR4DGyJ5XtzWtyXkiAdUuH9/2tSaxRC8T4N7ukE3YzuPvFiofn2Rx/STV7VxNFCa
fE/o6myeAZ7M8YOnQj875LkRmzmltHhKclc1VdvPZ3kEA+D0ScEFgbncM8uvMK1VgVQLWRgs8Ayk
8nKN6pp20fMGU3rlVq6T4ruetXWuKfMMkZFmcZwq/P1iZG1JeYtpZRRI+EkkGj6zYdzxVC8y5YnK
c+e5j7MglU0H/jdhe56N6MkKhQ6pwuwT2IZFRSjWELqeqXqQmEPekmaGEgFsnPVzd6Jb0L6yOv5q
/ZgVkOl8d7Lyy6/0HctSmwd7BzmXVZ1GckvLKZHfETiz8cixE9/MRTYlmaTvBWQxoSTWmGIRSBOH
y7H71RNL6BErpayFFFgSxXfJNvS5u+3lTR2vqIItQsjH34hWkn+kJflqmFz4sZAKpHx1SgqZOVjD
sjyiFWt68PbUhGjfGWAsrksJmwAwXOFM8Y70VA5MTBKjuXGN995iGH0xXmqF73fmzy01x+iLQrhl
URrQAU7S42z248x/x0o9M5kxLmQdXzxtLE3Z+0ooCqyQFVkr5YAK23grcTvXfRcOMBuVg1v2BD/4
mu1IswV1PuGVlGisgjxhFITun7M6oSa6sXMThmt3AtAX9xA5JiMgL2tiXQw0BdlC70RBDGdh69dQ
mX+CSBoe49Gwun7smHRnHK9gSsjr7eqzpZrjcyvF5/ZTaC2yTip0VIsZBk8C5qQJGnwiae66oa9I
9x2cQARlpiGe+Eo3qoS/HoSc0QbSh12RprLwWwiKMdjB/XDTYxXXa9oRS5jZRcO5wUQBw++g9x4t
Opxs5Pl50Z985FbAo27tgG9r0O/n9WRQgPKaEoM7Ynwtzoi8v3j5NBYBd1scaJXGybCCh1PM7S62
01u+HkIY5GOQP0XlyoRk6ZU/+VMUUv6ynI31Diq5TUNdH/Qyhx8MXxDPwjH4xSk5AJvABOXq+M/9
U0S2xmieqK8l7z/WRSQz/15Y8WX0kPMYMOo51JSCUbTY5aeixAKiBMwu/9PbAb67q8SmdpIM96/f
2IaMzl3m8/ZLEvs4kAHpRCW9N3X5dT408KqTtTZ20mHeSOSe61zJ4HnGRjgXtCBCkHf0/YP7lr1p
t9BrdMKGV2xHvwFNKxEikIQmTIRKGH/pHhpqCYipAHBr/ApX+HmYyk77NPT4e+t/pEP+FX3q3kaP
GejHGBG5qsWCabPbdfNtxgR1rod9/Bf0pSQFvhLDBkz+gs4Nyqxchyl601BIA58A3rJc8t+pA1Pj
v8IR2Iv+9+EzF/FRm+wMlL0JEBzOls5qYg9EeFp/RoTrloW+ALg8ExqyUFFOZzyZG45c6NXvaozq
dssEQWFcWaurk0sBrwZCjcQw41VoctzB3BHcEK/7RGkDxv2O5+oVXzJteke6EOVu0rhfA0T2/75G
m44fD01tlCIOzmIaMJNIFpYPpRfGSbWpCx8u2ME++5qY1BRtuok1boELKkucgqFHMDIFkgHHwvQL
uOVOjBKN/sSasLRghP+Yu8gs+aGY0q0G1Eo8Dt4/IE61FmdEpxGXse1vtKZgG+B62UzPE424ZrzU
EdJKOioTlqJ+7XnHz4KS2MOmtP00kTBgl26D8HJOhP8L1IoPfyojlKFJzsCTT0CJ0rHE4eqTh3P6
/wy65z23CN9fTFgdnxaCghQcwQ4KnELHyhZ7061GvUhSrUs2HLNxOLWgrCixSxhdiIwD235fUZ5R
KivNti+ke8z2PP7Sxh6V5O7Te6poGObg2nkRbCeAoADYZmnMqHq2Sy/SiHEWHbyMd+kTDGkLJrs8
2ObG0zyVQQMROIQVvGrTNXJKn3nAIN7Skw3/12AOtTeC6gY9efgwzM0e/YUNqoszkg9H3UGZbSOQ
usvGjd5nAiHCCj4Jc9e85H2gfB5tW0tlKWT+F/spkOum23Dj4hWaR2loeYBEj17Era5Dcm89Xdxp
ckAZtqoNmeNiJiddmdL+tfyzd7kVa3SP1r6XX/VsW4/iYR8udy+ANH0rye0VnjkthU29jx5CNGdP
Zvr6GnHi1JOkRYNvuw4LHonidhY+o/5NAGURdbabo7qYCUnytj2g4dgYYIRG1z4vz8ePm/LTLALv
eNS9hLlP+aP6HZi+PrZ0WpSHZxcXGIvn24qyuMeM3qzMzywqjTt303D3VBDPz776HEnxPuNwasy5
yrCuuZ2UxvgAPjVWOf/fEdqVbYW6CdxKOaVm0vB6Z32VzKfSGhOgMoQwUWTwyWVVNY5ePbGL7DwN
a8wAnTtFxZuwp8KK8sCWj7riut4puDw9m2TwiUbsGHm70Qo0SErK5C53n/OMXGJYxE1AvjRxOvDy
0CLDyHUIYzL+MzRRveo33J6IZkXVuItn3M5+RC1vWam25eeZLl5kZDhkR4OSJrFXzKpmiNo1qUu2
l03VftELOfhA0CnArvPKvJaFmnrXKA64LOMT5RjEAMQPqLaPKTcGztS8yhuvXpNRKCgrxrA0GDgo
Nk7mBoN+hSx0L2gdvqSUYlozrqFgo5cxjYlJvkwkBnLIPERyAr9IuKnwPdCjbYXKgJ4avo0UUilh
0uTFIFqy8x30pquSX7FzWM/VUh9tDvEaesD6IfklcheXTduK4+Sykd+ZTDYrVEgHW0BBq5/5R4ph
nuVSQ27JY+sJbu0JY3FnIOwGnNQaf44p5LjKYFoxminnbBaefuafHp0OquBXi2cT0esWnuY/0g+2
RftL7qOLoG6F0HdDLN7rLBoBFw7NGjmhc1J1/IQGAMkW21fzxrhbZhZLinBSnpR3TOljbMOtFedB
ZV0Nb9+469JXILY2N8eZ2RCR72ZUMxppp4Jn+TzD0Fngqo0NONo/qCVypOgaAsJlgGEA0PZrBUhP
f2K1y7ZJB2aRZTiU6Ndjl2NmY5vTAW0PEF3MsV20vuj5gtW7RbfT4Ny4UeZU+E744igv/Z3MDyFR
IzArpyWRfKCJmWhQfdsYfQW3Gea5mbz0MFVZfskDRbpog/KhkEKu2ISYwVsgM71eZ8FDbjrsi3Mg
KTyysHb6BdoAdtJJ3Xn8xBD9pmYLcnibnNfr0fkCECFTeUT/PIrvNbZyDvH77PoxMMuFfnC0uO3z
qghlYfQ2i2u3mHfot3xC0k/epbucxtNdT9gjg/shjSHUKmAhRrGUf1ppIt3It1B76Htt5pEEIBvn
RX0XIJ4ufjbWA7km5MFgVuLQL/BxdA7q1MT/EzHTW/MaxPAuwMHnbT8MtTCqT//w1DJ5WruMgA6e
j3a56sVHiqGABOuA2o8OAhm/+odLIaVSgccyBZkDzOJx1/a9+PvS1ePodTwepP1CKVyNDrk1oPtD
OWV64d3JFC4riBvq94tJbsJFPycIlzSSSDOBLTmUNkNUoKHKWwG0dFrl7mCefyhkuVIv6WZsep+f
LIpUD7+hrMaAoIFDL0ARi+xPaIBceXMX06GllSS9dOorZw0KuA6Ou2iqp2vH4n3d6vqB+nAOByr2
GlLY70K8DwQCRhtvkRhS+/Lm7WLruNA+Gcqp90wcZ7SW88/KV0d0U7HG6VQCLQztSprIsdYqilFS
2mGVPHumcNKVn73C2Lhf3NG4fxTH+TnxZt4pRr6LuMQCoCrCQAWmrEZILuGPUESIWKZxuFAJLqKh
Ko5lhgFRKOSNToX11RgooGmH7wF5HDSV+nKPPRk12P58sktJJv9YZ8mla/9ri8Rvc6HxWW9uzEcQ
N/ZmT8YtyHFz3hPHbU0b8tJkGag77kpPgFxifyPE+blzpzCcPTbVyc+1/pUEfd8rRUtjXP+Pjtio
9BJCND8VQ3BAIj86WeXrkntx04yzOTsnQP3N+4XHfX+14I6x2L4JU2thYbdqzQnJPmR+DwyWdF2F
LZSk6pfo4eqPgbvVfbNDJ/r6dy8WSNs46NgKLXXCN1HmsvlZa9fnOGNNkAdvoexYopxDVDcfBxkj
mNP2w4uW5sKdiKvx2GzLMEJGPbUbbFCxV1TzpJB+zYiQrGvx1tRRLLk36+++OG0tWGnAmBf7Dpuj
YA/o55UxDEQBx6w0y/xoq+jPYbsRfUfMkO0BU9Hw+LVtwI9BWn9CEsm6NiThtSYHIzcOjE2Nsa1C
Tfu3feEPFrDCbHSSMogIFesSsgr2mNhJqAmuOWP/VfkQ0Rt9D2dbOIDLNVacd35zL1140k7ODmdh
b/8dM6lmo7ufBfO0bm3AimArltmFeyx007UC/tPEnBlsCokXnq5Mt/NKU8oW71StiIiKOhBXKnNs
QS0PNESt2wSPQZqNbEbMSvWuHcUkNo5HNR5YxgUQHFZdmvqzS0gRLXSsZSMPzlHHcFZGvmFkJBxE
WcL0OGfcav5d7kVM1bjWOIm2/uXypSSMNW4bjt4QFTJ50UpYSpttSuTBfZ/xoxy+4LVphb7MF93F
2L6Cp9QPpgATsZDKn7JrEilqT4BMUkGStaSpS5aW/MIVKI3lVrL0jBH7qmuiFVgFJBa29t8xN1ap
A4tDUY222dHzVwhQMPvDT97aZ1ZUQ2naQHBwuTl+omjXQU9wC+qiDMCDOVc0NstipVywNZn+9FQK
hoTafN3HZkftE8OO7ybcLAz89HpCjl5YAqqyDMUpjPEWpC8Q060BndUytra7d+cGl17lxt5/UmNQ
9zJErlyOOejkrGxU9thMWDJFU86KJSniZKkJ1/kaLdCUO880F+LPBpiAJYuvYssFZAf8eNY8U+9/
g3erj/IPnGpRzHfI9wvKVtzStNC5CBDTM3j3irHNzr5ljzuiVv6FcfyTkjPmGh3uoAs29zKFUCQ1
MMuBzxHfzr3bMSm2czJaYY+QXWTlNJNxxaXa25t3uTkl5rrfT/IGvuCeuNFddOYcGOBdgRsDTF5q
Y6Fo4NG7tdEXHIR37I8Ud079lwZYxo4PLk+/td/8T98xehqtfouDW4WZGbYFRGwv3N2rgMtpF/Ro
35k3PYoPkJWY8U3bm9X5o6hXbpp2SiAlI5I21FrwR6AvjUTqKTT5ffsUZKhfB9F/0PiSXtkoRM5q
JMWqyqOHTL2jkB7Eb+0KSWvCvJ/I7j6jhMtd0DCaoNv+BVmnK4uiZ3ULH7LSBbXRkXV6v3W8Fe2H
2zraxxhv97Old7uff2lHSeE61JEV319s/BuJXu0MpsRKh6OZXg97N5Qg6Rkin5b/zsU8W/Xn1/aQ
kdlhUhD0C9a+bRfMbEqvuJWQulgQxUa9OdgwPHa4Ebog9WdiZw8qrXgupQeyrPIp8Jqfg1mtPw6W
XHeP5pPlQNSDAMA1/wqgYneSB7lbFEWzRji4KCXmLj9lNejvYr//QnweNNeBqEPOIXOPW632SFBX
RVw+b0aNLwnL5sTYJdDeap8vh8FnZUXHiMf/dbuALD4cuGCGX1d7kd3tyw9KhpsG1UAYycrX0ORV
INQTbaDrdE3Mnxj1a3GVphAmMdCJqWGgeqi7glu0ugEBs/ZpeRuX0OFSJCtlTKWNC3SfmST+nUD0
4xjdvXLLPPyu9nRpKm1O5iWumkYpytyb399JqcHaKSbcRIORRApBLKjVRhhXeewESDZrNNeQ2epD
9t/2bmnt9pPHnUlsHuqKoiiP/fK1nPT3g93iQpvqrSxk9EC2dNkGzx9c+rSHfmKfrHOH2ZcyFYHT
NpaI6RNtzd5mU0mcT+fGwFnthBYBplkkrW5vHEEw1xIqo+TaLpapvjI0NOHUv49fgUrKQs9NokNq
HWX/XEDdMvWP3DlTMQcfFWjKJqxGmDIxJADmqY4d4S5fGnE6/RwUaIkrsyAsNYBsV6QMYkUd7K59
o2KrRvEU1Dz4Q2B47loeM7JXNirNaVs3lTDSKpMcjrhxwo7Ga77v4xalcmoLTWxk/WPZ5nuwX5fN
HrU5WO0wC1NY8DN7QfcqlmNyhnaXamhtjjLTyKxMcBrm4jA054q5C8Fz+UbmwcLpbzceEMWmeXJY
oqGdBMAoUYcGUgonMRaQdiz6ApsQGaXaFJrOiHMGP+ZoD7+ZQ252QA7Z3ss7d8k2jBaOacoEb0VZ
8YjG9TxAZqo72wBletYHcgbAWN3im3LP8rLM/d6kmPRR4934DVHciRDJ9nE7uun+PTTOePNBQBJJ
S6dsmlbnpWnF4bS6wJ5x8xHr0SSJHZfbRlhm2c5z89HkYyFxWNpPJ6BrKBPyMG+lLcELkPHr78F1
DD3yga531LjzYjOoFPwPBdYHX8l3/SXpB/ixclxvBI9Bsi2Xthf+hvPsZi7Hm45NKOddRwNYbROi
BVtXHY2lmfYQVSl2LYVaOiIPlFFAsNalUDdz6TYyoj2I68Yqu6mL+xf7eJVXs0D/tAmYCU78KEU3
tada9i4Rc6NLGLXBLKFeS0MsQhD8kAaFRtM95cWZZf714JrFo9izer1OG0VC9KJPujqxb8ABWFaH
mKFcGjEdnEgGUkxqz5+nL5VlRReY0U0pY6hPaErI9mwg3OdhfNjvV6So9WZarAT2shqlwi6EBYIb
yOdPJ/Dt4x6ctysH+i0Jb0/Y2eGqzNvdpECka2TeWn0D0cMgzPbQ/IXiXW9Tmy4/4hmbfGCmGoqw
U5tM8GK1ACqH83biXONGw3/UMWY3fYw2ekscxXrhcW8+BiaRXMu4keyNdE80ff74NgpmoxDj1+Lf
COYQOMRdYOsIHZRuHXu+2rb1kgR5RGU2A5aZ1Bk/FO7dSN5gIk7iKS5oWNiDsxG2ow0OADjZJT8s
ZQYtevNKYdlts0Vdbgx1qYtugKTuUVaf+pD//NSR2VfAdbS8iqYNS4xErmMZjSOCByj1Mg4t97ER
LqpZJDmNXkOBFyBXDY/3uwF0IPZnu/uP+jpTG+wn88CdUS9QFomsOMppxUKj2czwuCQh84vEyxKn
+vmQWdbWfQT7OYrQOyom9gYvbd7PC95yEtMRE7IHzn/MUfXik3ICJby3961MenGtosZ7rBVhK9qN
S0wGge0QeCIUhz080qaaXWVTNreg6xDyeJRWxIFVTHu1LTTDEfW5GKVnKG+vZ29FlbOT3BR7bJKc
9aK+Ppa96JMYnvs7ZDb1bu8UbMoKCQivwgfN0EXw7LZ9oSA1zJzosfgGFMM9zIbprmz5pc4wTD5B
Hq5Pj/jnRznj22HxmO15Cp6cY+DrBa2kBJfCDDF3o652n1G885ZtXIpWmbPyo1FJqVEZ5flLvxnr
SNLwqsh9CsRm+0U4YubZ+NUI09Yvdt1nSgmM7voI+CIUn7JPOViFW/tKj0TdRdXEoQZbO1mbAi+1
nTLGEQYWsafDl46iruBPv1PL8Q8/+LydD/QQY1khQ8dqa2HLxazwgKsB7CmlN3kw8nP4FkfdghE8
MkMiX8Cq49+1b2CJ8ScpvHnQiB9cBt0HAZSGZtIYpfsyz1INZYHrftVWAxtRFh8QAPQCIguMFawn
Q8N+C7GZ2MeaYwvEHWmAETY0AV5auNj7f8T5kqmPFRWOHG0DgYcRIl8bj1PomYPaHZoVbqySoKKo
vUE3KJJaxlf5yKt4/s87AELgLzE38amJV3l+JG12sQGxosDz49iUMlW8CTlG95Y1leiGC/9Xfwwr
NSPiOZdb3Rg3y/BbglyHhz8b2SgTWqnRPSUAHMQlM9gJXMvalIFmUhq+Rr9OanRWfIjgI6USwtPR
qOM5rb49BvTG/kspI2vGBxQhMKVmAAz1972dUBxWhvei+VseQc8pkVbmkxZ1l6zYo9Jk4i0gOKZx
3ctfQ3K/B3evvBJHnDGH4RmnBFn25I7KHOIj6p9kFVfY8qaPdkyczzcwM4wzme9gy2B9AKt5k5Bm
+krGnP8dwdSD6cP/Q/G9GEhhNLz42OsVRtkK0lrTEmnIeAkg+dPc5gASs8TZYvh7YT1zSy+MVuGa
j7GZBSh3xAbcGN6pHdcch8CvMeNUFMlXDmfROhuHxXMc8XUX90GUkmCsjJnmAlyiO40SUj1hYqyS
nzuYvhao5Yp6+KzxnHTnso/8Gu+Y7ZHgkgztfZ43+0KXbgFSeyqM3LpMafpgMerakQmhqsrrM0vA
IJx5sgXZJJr+ECrat+X/jj6Jb44sPKuGLrKqY4mCeqUdLgYjNkowpS0qDKenGclfm8sM7POgXPpe
rmDE6ITkdBok0S3gKVEUuhkzcYEVMcNCgOGLawvEtL+smcJ/PLfRgTR5OaWczEyAHbUNCBkDXuVo
n5cQCDjTPQx7wSAbiaiEY3LvPnZf+dfV8N5b6NNeBBVBVLwfKY5a+TzEbwd2Pk78Ex3AOFF+H7to
IuRZEqPtzPMB0YXqzG8fvTYUdFvqjXJ0q7StuuRMbiYjW4mxfU88FoB8fOlf3Cs39D8oiYtAeDCJ
oFOhq4klM+mmPsGfQPP239aMaebkac4FFZHKm/Dz5aif9v1kBaS7s6UqbSVkRJxJc8dSVsWLkbi7
z5Ye2UunKreSrgpmvnFl608ObGpFc47OXfui9r1kvCy+dJEBtTPQbkJNmymKPh7p9qKU9agsirnw
oWaw7cBF8Tam5eJ0rjx9j6siqljcx8yFKKL18Xtf8Oht64bFm/c5U9wT5SO47VbgJS7fb1cDTUxO
ctqPAy+SNFIczRC3JaGNgxnDOFl1JM/F6aOmAz9SApmlNUeHitHflpguAwzuFwc/hVGsxUKYU8Zh
w2R6NqeMxmjU6ptNVO6kmOF8NmeghaacX3SKrViPRuabyYr4DU7tumPAXdfv9Vrl6c7XYN50LCV+
wN7082DYCL7jByf4cmM0nGjlGGHXMvvRcK55lnTXW18w7PJCiBEw9hDSD0Fftr0Qw8UE6Aq7BOU5
fTqH1bzfCG0Ty8K5Kq0Sg9nXrnTWt3Vxl1nTEkVrDjpPtqOOQ+RUe+T6RCZ5wNSjjjKkMruA44or
cNWBLMP33GDeqYN94CMV8jaCtr0N2AgheABUv3094lFUPuHBYlpC896rI6YDUVkfbzFl/q7fHPXR
wtN2NEvKA6qYFfsf2PA8FNKtrT4Xd9HnMWIpBsBACwgzI3PMo/Afhj8UlYCUdNgZkRorZDvEwGIp
lX/C18SwEzOKKmLes1MX4zGi2dLfUwvdkuQeaA8pracyuceWJ0wBjXYnbWAM0pXcgV36KR8dxpdd
moySITiQD2KwD0NCabXG7fX9L5FRtA33vnavNqvWq6/7gC7UTbSD86vMOyYMD55JZS+aoesAXjvI
S4cPTmTRG0W+3F0kPx+PKY/93dFhSnJMtQJiIC1UmsWKP13e2y4KA6iH1ETlJwFZUtfWcdbT0cRp
4pN0QkvR/LRlv/QqFebD3d6sg7RKgvhqmjOWCRVsC4ke4ZTeB9crr3fCW3ZOy93sltu4ZD0/NdIz
+lPuLVgLcC/Y0zZljOySdoj3CrCA0OQC6R1VCsWyfTIgyY1k8Fu0c1M0WCiylx7C+9tkWnyVwn0W
7mNq/JczHKzF6u8+mDxu9MpHOne4cRvQE7faG6wwGXCf8byD8ckCMTCimYQzYDncFBAkGtT5IAnQ
eyivPWHv9Ht/XkZ+iciCQLYu490PyrkEJW0fpPcxzbmYIrN0xtQ4jW4DAXWWOffVN2LaIHi+27nt
GIUJeIT1yknkWMFNjO8bFDG/OgQSLy3GSkEZ+AoAFBWOtVHptDd5xDEsCqQtESn947nl1DSRPwod
wAC5Ud6zld3Qdw+8u1c4W+zqiSAj8XYlafFlwgnb6UtI6mudd9IKGHdatp3oslf5j7mDbh77DnuX
KYCTZzB70Awp7q3yrg+9R3d+X9AgnvBXksGy3Ku/abmtueJZgT40h3iCfVFrwg9hCyJ5iRjt1Yxq
uVUsNgPEhUghrEATt5PtVmn9HJ8P78PHoKiYdKOesfIJzcgJOc7HKTZ9eMP/yMv9HJoiH4e+lEi8
WKHX9rxvmgF1363c/dhDfXQfc4nvnWicQE5/s/zrc+seOJiXQ7K3dGgmHEF839tSvlQLp080moRd
ao36sRYKEgEJQogbMf2N7mgBw83aDPoq5qLhAdfELhoFOg6UH9sqeTHjtBSn02Ys41TfHIsYZXZ1
0CPvyGdemjiiXYJgWcouiCxy+LTzObAk/So/GrENU2/0B+NEJCudFHpqPL0aVp6nFaxIkyhgKMst
E945REzHAJcjtTPxS/3pfMjwYMHeAyRjRxxTe5gTshjXZeCmzWmlprQz1tR4CgHUlRKyhKjt3Tsq
U/EgqxbKePLiIP2aSAewJGN6GLt4NpkW7Atg1KMp1qXQ/RdxNQstVa1Q4+RRfFcDvDF7SUNPfH6y
/UDQNCE3IuJVfvpSeVVao/qEpecWx7mtjzEEUenS6MkOxEFS/heio+h+NibXOj6f7h1h0lWm7Tlw
O9avSuD6esT+hZBs4pU7CbIjHU7nxxjcdtRklLOnt6FeJjrZh6v/ueAQ/PJOFHZsmasBJNE52lcP
jc7yCd4M4T2NSPn6ExUgt1zjAyuw9pBSUaIH5wnCZinYytWpfyVPl3Fg667tWchQGLjSskpSW5Mq
siFp/T8y6tQmV1aGAJWxm2fEU/Q+b9gOYLZeFk1obgQInkXPySgZ4PoYxtakmAnNNRKXXpG9AMfl
7HF77H6fuO6dX316QqJPEC9fKlYhbKeoYfEc64UADIv9zLwrlCHAboxEaKY6cCrLc8WZIU76IWEA
CK5Rgc/Xam1vCxffxuUcx3CG1ZkHH0i4/rrkUR/1yxXfzrsjoQGXB0SpTEwfgxhb3gchUoQA8XNA
aP5Dwwk0+gw/6psHzMHE92D+0IHui7gthaxP8mty2x+RpomNzm9mnhiMpBqaGwpAiLbok40C7/3L
Lktm87zcdj3HcX49aWnaHFxULdPiAKJqpfqPtbOJBhrVgdWblJigxxWphTafd/hYEJgwcdkthtHD
yy/mRxiZVuLnnaJSH2TUe39NVa/ltinzq2B7l5fSVGJD3mknEUwvhNa2HYC2jyR9+KYOuwmgS4FC
6OsF+zdZ4mus80HdsZEQrxYRuJiTjnvJM4BmJneiMGv8qa5Eml704OQK5iRAtlcjpuA9vJL3I541
xamJS+bEEEVX7Ua6tYMgej5lK77gxIXzvpveXKan4xt6VW74Wh+suBOzUW4wB9xCjruDiw9WkSlb
zrJ0Ka+25p8K25L3KcE6CPYhPSW0+qmfKcGaYISGkMFmU0RA7W7o3jDuvOQAHrOx6adRY4kArH0E
PC7BRa0o4ArFZ+ljugqG4XoNgelv2llr2JJiS3xTs/Sy909TR41l4n6Nz8Zm9HVMoCjGfMsjgP9s
nXbQM56VYSuRsHdhdpjd16IKaXeZWglWRm5/at52+R0J4ev0gy8Zdo8qxdNn+1rWXgdGy6lsPu9b
MQ2aTsBm+lioynnMXdlt1DNaFjQBRIJ+m6E/zsFn3WRvmdV6bU9jP/L481NVwh55qT9qX5b/46tZ
Kcbb+7zQkfBcZqQ2PsM39Hmmhb//UeKeydC/5JCa+ZcJlVTxJB+73jUMGFTsd2o1wb0qeLZ5N50R
AczyLk8v77Mx5/FmimhqsrAcr6oaTJQKCWC3kQHrSbYc0O4dkwXGFKRAXvUFZ5HuApmb5jks7/rF
o9zufQ/x+7Dgi0i48bBYUayhJui4WL+M8VthG7hApM0yKg6IPOMchCyltUHCTgu/aB/qsCoIXa8A
PekxGpB7f6+7VRMSmeXvj9RLwsoGrXE6qfOXWMZVNNvo5YnaywVzszFSm4Y5ZT9eVfTnbcDb6g9I
5Y9OVLcrNSv5zqJltMhJ40g2I6eDKG2bb1ZwMm47yWYGwrOcvGGP03hISSGH8TtLtwR9onGQG6Mg
bklU443NcXJMIIDU6dm5+tlKojeYd+GCAcU6+w93sJla6/Uc6UMIBUrNxZhVdc/SQ8VENJX9syMh
FAGsJTQ7MpIPCJmRAFa3g0M9M5Hrbzq6M6w17u2UmdM84BMSlF6Zk6LE8mPa6haC/s1MVjkccvrn
OQ6MPx6W0dW1oj1XDK4wRvwI/GLYehWpc85gqT19Uk64+k3S0LoNUWK4t4/yOT7cYS7uCt4XW767
IZpEvuoDVnFGdUOSVYEKpbYsWW2lUKKIPOORByD4gmFsnV7wZvCachqMeVfahGGlVh0N8gPUN3/U
C3C34DwPDcvMOWR+4O8rUO+mzVVnKXLGKTlOZEGb8+bpRZnt2tVia2RPezIPaSnK1ckIZlHje2R5
z6b3HWfnFkfrna5ka4zAbYv9iJOf2oQ6ZIMMqXhyk463mc1x9ah+2UoNku+gte+Gm9tChUbZuwk8
FB0UHJWrsvw3CxiVvVQn3QodwlERE8sMWb73laWnD+6KszDj4y7eZkuCRk8kBSpc5IG5NW4mMVLK
Quh7O+Oy2ZAM7A0L+fplGDuunrSgT0/Twvbh3xonlRemrDduQFr+HRaIec5hZMnrVc8gBGMeGtYl
kqM3i/O4agU/YkVM9+jJ7ZeT2yYSYSSfB3NInd8Xd6XdsWHAl7QvvAATkHCGwn22xHLeO3xmg3hK
GJKFHSz/8t6W6BBJ6pl5099F5mgBS+BmWi+EPcKo6M6PRGtKxdePDiUFTE1gnRAxPcAfDjgm7WA/
mecBTNH6RkkCaFt+D7ewjK2cpK2dNHiTIaDJN478/b0mGLnmizaxz6Y6P+515CTXwxHk3y/gJnAf
yUMpts+b8wFZRXP75fIvqxhZPQEcu+fJUTE5JemkpWpXOQCuxn+khPjZ/4uGTSj01IrxOKQaswLZ
Ik9fyrsOjIRIvpMOt00Tak1F9Q3NIxY5suU946PXhkBpahohnXnGB7ClZYy7jGrraUP7SBtwtbnp
B1owmGDX8/1JmHOdqSByO6qj9kZMNNAO9BnTiRsHIPeg9GoMag9PAs2yh4OHkmppzvKxpzLGIAD1
h/2tkWNlB7tbgy8PaqLqjsCB2arIyJhxEtlb2OB5SFY+dBDOLm2/uCm8nIH6lNSc+foxoYXr7P74
ooHYvxG17YmQcAQM19i0D5NzLoXfqkQep70VcRJXMAoTHLpc2AtGYATlxCKU6grTjveUqrMyb5Ra
hi9vvfNkZjWrkzUsoi3cMOR8GiIqWD4nOIHe0hnMBmA63tefQZkKsBrNXYOMEU1iQD3FsAn7OwLU
O3zHxA5h05Aav8y1xryeBn80NbJCfz4t7IwXItX6lbx6QN7P6/95eH2taqn67KUZ1gmkvkMopxcL
tsWruyHXOBnGLeYDTDAsD5aYhKEYy3nZU749mLeY1P3vt3HO6NQZXVndpc2Zo+vj7LXZWYHs8YqA
kOVb+GJSssZ81/IDJm0abYJGVZSLF+7AGLM1cVlePTmYLZPuTh3QgjTw7OIrTfknsaSlcnr+ilZu
zw8bnnLnXWCejh1VGfleMlozsAl3UtBbKlRvzWvkTUUiNv7vyqhClVsxrei7v+mMamc+LBIH9JP5
qQ6y1h16KJSPYtJfUO+be/CIYiGoJqq1p51sfzfT0wYKsSpQxxnGRNV0iZGTKY6PAkVCfH23Si+I
GZEJ8Z+2eZsWS5ndEckYxz9DI04nLqCx1r2WhYDJE1JdcQE83I0vOBFi9OeAZcuw5vKhGPFD6ISa
WtGMs5JiSsd71eIKdqBTKaDYHWwPTgmXRjRiI6ritZYDrqbsT6XntmOUwG8A/+ga0uVypzd3EdbY
Hgn5XUtJMXOiRYDBUg954wiDiGYN5a2b4y2YhIUHvVs8QEgUUoLc82r/otlrP97UasGYTaWmd0bn
exWwY6G70pd/KHwocV+we1e9lhUyYTz6CmwGGAU0JtwK9AgJHjkV1hUb7039HkMiTswmvp0D/txN
lFWv8rVU2OqXwhQWt0FCT/GSzPhh0mHrfd1NzPV7+++E9IeEKnk/DhXEkEtOuN+Q4iIm3JcLJBl+
LSNvgYn7BiQTSbtVVMbCLqZVN4ceu6SApoodcneJwy1G+fA0L6f1tURZ5yQF6vWq9D8bpEGyNPTi
uKDBLjxtUZpTEWTSx3u4bX7ME3oJMtjldDQwyJXungCfXmFV7/YHZTvZ8d90AvrijOuT58hsNJJq
KBhTHFeVa2BVtwcBINKQK7Nh2Rij2cT/lP4dnwlvIunr6pZl++HVWWTkefArhdrnghP1Rvxs5Eft
aZ+zvQbf+YMOvmoKgyttepCYbRA2UwgunRfFUkLAdDxt6UFATSLjyFYEWKb18P2UOBaGZvnOol77
le2wPy0Oefuft0hjumizDP4hdgf/3ZOalqxWcPD/YdpqurYDZz3sW9L/Ce+/3ZMc+oEyRGAMO/fA
BAZy+CJSJGjpwLJw3LmKn938OCX1ya0QA9y3VWQQ112/EU4TwP9NxYaqGu07Nh9mr/rsnPjSJSGj
F9M7RPO3Ba56+vaXwJh8wQEXXcuJU+ZX1nvz0km6YOVxH40XJsKVL//TnNv00du3vWIJ1ZWhPmDa
aE8vg6ZmRV9SLRN2tJiO2ezUHGrzBcn/ssx+2jELx0KcFDtsC8162E9XTu18x2GYU2lUeKszAt6Y
JyLfy2HkbtS/6mwNXONfLXSFC5fxv90Qra1HuJLU9YsPp+Fw/9QG6zfJBcOBXml574kr7DwyYxmh
wd1zUmoGzJXolmruXvAwLnTXv5HyAteOOPLgVPk3KKT1rHRZO2XxlORcxFZVM/nTGYrExbadDK0t
ZEkvY5IgU/U0GvAwsx0C5SrH/JmIU+XtKdKjjkUGBH/Nv3s0/C1NXsiUK5eJHvW7JK9TjBbBbX1t
qrd4nVELBJsrnZiJjS5omZSAE5eyd8O9Rg+O/wMKIgmhBkvcdm58T8i8bUheLo5wTNJwTzEkEFU9
pNRWorTE1A9mZ9+OLCLo0p/vLKh0/nw7mP2NF8xGLlEBUPHuqZ40VMqq1GSr+X0Qwlz6xzHzKjPM
1QzjI8iuVwWv6xRxqd/yISVOGqSAshhGugsedkEI03+KmaGKDesimfADLlb8O/mrfGiiWFS+IAIS
LbmqfkwhQCfACt6bwqMyf0tn8GbzLRK04/VfYGqz9+JJsL7ivTTjQpHiDBOqgh7f/IxXgOL7uBVQ
r36FDvGoPH092/LMcsjvn0wuqcJ32oHh0Iuzp0dvzWCO9Ts9tGRk5WzdtJhEUUYhAJ++wEx8mxeV
zqBct1NDQcORru3AL7D3Y/lCkQtC0xKbnvqhHk2sXPjByej0ddurBH2dQ5ITwx9PvDy8QWG6NMeR
GS4jJoY6r+tiEQ5pYpIU8UhlKlmFWSbLE9V0f0EnlMh7FCIeoqgpCnTjLfAkMTJ4u4PFPVM/mcoc
+5W9/QqApitO1R80PWmEC/lD7Jd+f0gxFVF6ejcHX9KU5DOgxzHS4/LUe6KfneIqfaeE9JkZt0yb
qi1lzPLVeN7aS+xfvKDf9wvGdSjisxn6Et2A8MKm4rBQbRfWdbAH8z8CUW23rkbygoRjHJhL/ZCb
pMAdFk3101m154wGQi/YZ3xJqfY2/ozkq1tOZzrsdd4LsW+3jxGVcXTcp1IY3BSbn4eLf5k6y0c/
M4nW6Wpw4eXEc3lltB4wF5YzPREKVR1HhhoUyu3pt36Dah7nyTRmayRDHn38daBp1JJTHYyF5pM4
76c76DyfUJ1cFjBbQVlwXqdZ80NGzH8kVj4+m/j55Bz1xd+vMy+8Ty0LHMnB9zEtnwtBdgg+93BV
7YiHQVwJFizMSXfebxnpLZ7SnkfzT/poUEXkhGEXChKHRM4xkELkcxP8WFsjq/OXzAZKTNZSd6ve
AEOIoUSIUj1wO83pln1encBd+ABnmd+M6zn0hjSXYfaRXbmsveWbSS43UNuo2ApxufL9vkJdsGkr
tk4Yby3aYODH8BRkAQ34DfP0AW3KTgJOTp6lckzOOf48ESA11ibG3QJShQXMUiwSZ+GKDBRvzI9O
z/PQj6KeNwNXEzqZ6iyTNvleSrjQj5a65WQyjOHlahaEcMPDx0PU3bYJYibVQuiINidn1Ofj8ZiS
2GSSMcGpwqXkzPiXK8BXzuVKneEB/5XQxxQp3b62TLJhyskDkTVycy4W17r4Laly8PXHD5JJsy05
xJtGZkAS0NkSS1+WRxn7pU0CPgknmveBNNWd2UqhsqlvTAKxe6dAZH7E2RVZ3gJTMjY3MLEN4KAa
t7Cz0VrGIYSD/O/okUSXDY0E96dQfDJ9jFwcsNlJhFM13RFJenbCw9fhTYVeVgcji4rkx986H0BB
v5BB+4nF+EhMy8Qw6IuaY7vkTcM2mIRUD2h4SXxhLc8TwboFbJwPMr8zp40/9b8eXiGrVULpMPMS
fUKWKElFPzMs4N28+lgdOuQZq8w5l2WygN1yDZrn34GOaa2Wo8DRk/V+dgACcStSK8pgDWe2WvzC
qP1DYITOdcwK6R7p/YZmiJLwzbeU/6933cy2aTfN6YQhQ3VagCtZMREGRuGt9I1bNn5vGDNt28kP
n+R/5H0OXA/hBLGOAi5J3NYxuLdAjkJk980Kt0NzeSSzL4ubPmPFOiNA5Qf/kHXJor4XwSrPt33V
E1ofcOnsnA09Ea+BAu3WmmgNkARKucoFCzqWizMYAmq/ctOrijrtneF8j2dy07vtBA8CwcItwWm4
rVJbrlMjqIYMksqkDwzUQ31IhBV3zzWAyED5hLbmZ/76IMvlr7xv4OlHBaufNtJPqHi+MIOXQ9jb
geJi1gbNs/wjQ3hlwRV+LBHaOwQ4jnBrCXANPsFknSu1JvdFc3nHwRuZAXAcOJR4UUc1a5L3IMuP
tJyhzfQJuBX36lNmoMPqYyoD+mzGlk+OqMBsEcnEbGaTtHkk6bTkNpMixoN8f6Z+zbSZgGNkJo2X
+9kedxY+YNiVujgu0oEJD9ZZGywBISbV+j00P4j4Hlmv13P8aN2OAmOnztfcyL0GPNwxcPXNa/Qq
l0HB8t1ErLi8qDzAY4jkkrrfs5+18iCfG0SuNb8DurnpOn+aVe1pddiNjqoZvrklswnYqWdt2BHm
xbeaSL1c36mXErw0RyiVYrYnDriLBVwLKB7EZvtaA4qyvCHfhTlfTheMsSV6UqfGV0eXzUAYuKKc
+vfY0M0KQx1c63I2zXCCwZQQ4I4Qte6jUiBGrsBFgP+SkowWDpDgNDeEJ+wpSGj2VA0nIuqFoy/s
BLuMeooi1VpLrjwVNRJIdp019YVqy09YLc46xX7zKF/96QHEardFPKIuGKMpzXvBGWBA5Ne77yzq
20RBl1/xQC5DLLCxwrJCPmOxf+h2/fphceClgTehfW6cKoN4SewctbIR/Oz/2MxU5xWKfw3RwCFx
A7VaTV8wT8Ut0SWcLij90MqSeJ7lo6Oz02RJYgiDfEci9LpgkDMKmVbvJ9C8TgN5jXrpvUP0j95Q
DsaT+WKPFSfcrqp+tg1rtczLoG3XYtjNVC9hbJSnZog9in16KixmhC+JXOhsZ3BvhrQQo1cVnQhD
r4MOq97sq8dJpIlIrSI1RuexKWgJnkxjpZVm1UcKlBNdmfeSL+D9FlgESkoEYgwl1tmeX0shRZ7K
+Kchln5HyPuOx3SwDWhgSCIHG49d8//wyPExYohL52IqoTs0Y1jIn5a9p483Zl24bT/nwDsf+i7n
1gpt9N1lbj7TtQ8HDRI4Axuqnmz9dynj9VPGFvPVs0nwLEhwh9w33J3yTw4xiN01AendN5N01KBY
n/WCGhhQVBwH8dCQA2lHQfKi7zEJUeBmmHuEvRFzmuQdsa5Rr/0lnI/YlhhK6j8L0F18nIiqBaGm
XKOFVETf0ktXVR4RBFmtYooWOxL049z+aZ6j3NgfAfpbUfnBBe1+TO40jdq964GLQEjJf2LhPzcj
kPITA3Xip7kinQtbL4HmgYg5m0wOcD4jS8+AjufIDS48of67ByFd+Hs5d53JxXMwJYSUzfvQor7v
xW+//nV3bRnazpKWGLpChXPHUpZTrtyrfOe1wcHXKJUkk3lb+QwHTo1HOq7m0DdU4/r5/x/lxKDA
yM+7xy/QIw/l98Y76itbusvkz/PYXewEEuIuX68R0YrENidEwcxJXvdONffldnEt7VLny3BWYiLe
W4yRFR5jL25s3LLLiBRlL5HnD/8LRGT/6RmOqmNSxWVq9I42lWaj4I/VWYBxsylkV7wte9az0i/M
i2szLEX4pUjG7iZHk/fW6YINSLGKC2VPNToNAINVTmHzl9ui2k851JTfoPHJuAzc29qSwewHxZfB
SKLl2BWT0JN4C0GebZatT17YOnViJbUaha/daGsAV0Jsrb0o5IC1aZu2A2UOpzGxO1hVPiRVlKj3
vzd4AeNdPUDrbjCU9fy99b1rhbKUW13l7aTOOfmbiTbd3l0SMUj+mj57ryjRTvEadUab6yC4J9ZE
lx21pyitiVg5+R0EWAXxYx6RFZX+NMGLDm0savL+285T8d0CqggwpdvHiTmZeumC+umiukR4MDom
g+FUH+jXvD1Hq27tYkmiKrAG2bm6nC56Hg9d9T049xwe9k4KjN2AeToq9Cn1teUZj3TDGhoRk/8N
8TZ2mk9ci/BrxnhIrFnBo/yiroL4Ojxz1Eryub7VNAoybxXPuM0k4ylWBrYRMeYSmuPD0wxlWHKS
p1m+SeVk+EFAkqczFT4x71skjEWlbOucKRZAFzKfTQZwUusLOBxYAlrf84De5Ufe40qVIUstsbZL
M6P3roapvjElxzlA4zf5+J0R+KDKCue8ujPRil9aqXVG7BsNoS5eKRfxaB2QDZt6GJOSQeAapj6t
RPi4cqE/Tyqju3dBSz5uucToiXh8z2S9BpgLZrwH+cPh98xTiHhI9XhipW11dRffbdOH2wnQX21Q
1yZPZfRFdzbpRQpZs7Ht/QHB8TPeGeeMBryYhcwQeJtcBM/Zj8SeHfJCuUKYI2yzZM12f8ob7DU0
UXyiiWjf4Mihob3k5aBEBS6e98qRjYCd/QbCHDhVC41ITl3cvtLahDMfBsGB//kkFk33AZM57R7w
08OQwD3dD0GSPHCOLIpCOrx4M+eCCWnA0L8G9i8liG2DCqNXMaWvvzQ3WMBepYY747xUkZPfrpmQ
My5JfuTuf31yi+qi6qAmpusBPC2gHTFMqolEXlW2N8S4oNzMZfdnZm0aSV9F/ffe90ISeEp2OP/D
9yu3j30LXx7UkIm9S1ALQLyAmcBgZ/Tcai9lmYQcMPQJIHqALmQtsGpNqkw+owNhjnwWWMqgDuZE
NFOU+BAf91bbdIh8/FRmytxdOC8QUkC28d8k0thIIkl1YZiPihaBs3JQO1xTrwoUF77mrLcmB9d+
kFRLFnfMTcWHzMTbxjxmY00uZ+dx2VaX9CvHeu/Wg2psTNtJt4aoeO1a8gc+rQsAkNEtXQhrJ6GX
pi75yFghgUjcVljMsLEqeYe9mCxXHSxGq0PiK0ilr2S5dYApOokIyxFX9wM5ScBo6VAR87kj7ZpZ
j3cHL1+lTWjwQay3D2aOIc7ypVgofvFQHg4pVQPFt1jeQWyVSTgt0xiANn4C9FUNRK396aSGTIOX
wo3QuUjwUcj2p3XUBF6tyIVcQYMsS/Bklb7kyRbhuG2CHnXb/Yuy02YRPUnCSKWdHnRnuxOUQ20H
bvuWeZVGHjFla5sOBGLHGbaXC2yoJQtQ72fIbUgyf0bfGGplwpz/Xggm+IWJESJ3QIMSLNWS1v+h
0snAQ2JFwM5JYoKCAY97fNkJQvtn5tU0lnNSTwOdxalCXdRE/WWnjhsmjlgCJjfGDT/XjrZYm3TH
f8opXciHAYcy2Lf7VELwS/zn9cNRqn+4byE2X731ygb19QgF6UzhNYhoqn6ntaOFAlIUvbZ5socU
W6lLUUqzONTQs4uUusFJ2TgXcurGvlIt3p7h2QQZDLV+PGSzRQIkunXJTyD8PztgLv+bx2X7vj/e
BxBFhrz7n+vnkkSaCI2LkGGkvGa/OxTekvVGeGy+rcuieRxiJWJB8WCQsrAwry0BIX/IVYWhqt+b
zSpQkdl8aGX78Adv8NTtQrymzDRMwGnaKy2I6YR0rPGpJ/K/WHjOx/5kviXmKkZGma/QhrnyjeSf
1ZZtPElIctpG5OTP3q3PU6rmtmfKDUe4JXqmx3NyifxPL9arjN08o6PbkXEmup4kT0VyVDbndhe1
/eiJhM96QVZ9kEP/gQWLc9/Ke98bpCf+Mux1q2QdSa5mEG4zulb7A+yTo72llqT+jk+uRC9Yhd0F
TLqN1iWyEF79eQRYhJwOZGa0bQSoCPdcfvZdGkwyZ6NbkvhTeG9nijCGY939owDhG9aiaCdn78CD
KggkUo3bBDvSQAmuanuhNYDA4QxD/2kMFsuFUZalPg+pAjV7DygSyNGIqIgyPc3chiCNOI4xq5KP
Nm+L9tSo5zwKvqTaICFvl74M1I/e/FggIdq/txmKd1+5ZrPcZfQhIJy9SB6XUhq5XXGLb+4VmllC
mVZtqPuR7v6pkj2n2zzR/yDRuXIyNnR23PKY9AgxJe97uAvpgYuAevohP459O6AbxfnMeRy7azg+
rC2z2HBpNRj3ZFIcnhlD2TybAmhoE1mgm6QJGjianH7eh3lALhn8lIxVpXbONnVtrk5yoAKBNLy+
HZ7Hjpj8AVfshtQz7Pw0jRW3EF2SzcovQB+izZIU+m5KR3sihkKO/v55sd49vVBDTlKcd867XhB/
39OM/1bwpRkBBGJgqRsXbJK49l/e57JJ8nZa4cFI/O8C6mLhfdTzhsOdJwbdMWRHXZ1+v8Xd5CDq
Ibc7uAjOgclB2s2whbkvB0aaPkgpnNr1UdaqnQJFTUaAleQDgKXtazB/NENdcFe+rdzs2EgliG9l
vrW/1oGKFHKskPJ8z2P6X52/G4Vh8Q1KA3s7n8Aorhjwwbks77cSKRocjWRPTtaLerFP8OJG6Gqw
5If15LZf8UuBo+MDNI1dJb8ILxqWIUQeMG9s/Gw+KbT8Oz9vqWewnzvgqboITKmWcH8ewgENqOXm
ri6jVmG+xzMHiYpRz5YCFHnOhPFDVa4D5CLxJKyUV0jKUiTZ9w4J6HmLCja+zLBHQJPRMtAS9Ojs
57r8sL2c0QgAAZiVODdAtgVstkogzItRi7nmglGjJ5Mbbg35HnI2IufqzIxubimeFBKE1AKDxIXM
7GMhOLxPJSzOxXRT0h8rVm7XcQ+ZRYhKqeaYvtk//V2SXO7dpjjydQDJfsoJcR+EI66u1qtskD5/
O8nwV/UR4Vo3xU0EkRhhmUZTFdKjpppgWOqLg9+wP7Ohb1QmelXDzQ7OyfCtzxa0gQK7zz9VS3ZL
Nq6tL5bUqZSnnxRTYTZPk4JjR9FiKufvBHtAU0Y6lKWt8/hOf5s0crLdgbiRC9sdAGldDuK8j/6I
d2Q11jyg0mBEy/8CJ85j6SuJG4HXpFKRwm7Qo8y90yzNq/48Jw7mfPBPFVvVJlcEtEwM7rpvfBen
FJx9fIEYvdzlPHlUpga5hPkP9vMMfapFE4rdfj+yuuDKGdrCGufPSsrynOUYX7MOaQpS5B1HPQak
LR+IwcawSzu+Wr2hbDkY5pugK0myRoa4tvQxPAcfwrryxvNW4NmdiMlH3P7S19egppEdzu4yo2AC
fcduP9gdcTaZe0f3rqUGwcw7DBX0vY5FCq6GitecAF44Am4rh4tY9PVo+z1dA46j2RuD1pGg5WKo
00U7R7spxOVamRyTFXH5v7M9usGkbjEEW1v0h3sEPFwPF8F2//G1wFh8lq6kbRHOGr0IZ+DVm01Z
slTA0irakAoRUzFRJDtZFsgThrqf25c7cUxhK87ZkdBSVTjN6BEGrsLkeajFymZ9ADKTc5XPxtf+
UAiiRBeuFlegiEXhjzeBZE9EHeUgiLRMcOIZSwLwRcSyUzRUKdq10qzxpmevjLojfj7Ug/DVvHLq
a9k8VUhqeE4w49QqqnrY8pj9RsHojEQXB6tiooEgObeL1FhjY/B5Qr8bJ2JXc/s6a/aLsQ1Bcin/
58Kj5X9L7iox4SDz4NqL8KpNfupqvLGbVH8qMaX8mSEpKFLkF6vjJszr+4G7jh7wcAfSJDk47/PT
GmcD+BjZttmG1L4XFD3ceV2SQJhdE3HVn62x3TJhxMJ1GBibCYUmDS8JXfcgBbPbBC8bQW3BsYF6
rBe+2CTqlHTPWoNIQyu3NKwMXkuH0L7TWdMjH9Om1hTP0/NUwA3a2qXWcflF1lBp9/W1o1Miytnu
zUrF3ZlLX6vTJgsQGxrL4mKZNBtvp4AZqmTWrsvggNtYJ4BZsT2+SKl5t5SWcYimbGxszLpxtqd0
cl2jiTZ9yxHDbLz9RotCbO7HhR4SwyjcG7yJKflyAKTVWehnqCZsHknScrKzerk/IIaIpF35fMr5
Jv82F93PcEnkAQEJ+u5TFzaWtFvDmutzCwSbl7Sz5IBC0heNd4BKC3HA1hsUSbX3d2E4hJye4qC/
00wy8YvfAlkFokSgW6Oq80Df7LTZsNUYRzbvdQ224px6dGlOZGJTCf1KM2hD+gbxxSR/aCMOtqri
6ngIUmEV1tsncbP9NFVcwbK3JQ6G9Qx7PUTgnfN/KqX1DYXggpqkoW4q4J/udDZ+geMNlLUhyIOS
QXhL7sxzujo8j0D0z0MOGDdQ8nZtuq56ck0rhyYlmRHNaOT4SmmiW5OW+hhYu4msN1oW4hcEifY0
bUXrrtCZ5UuND4stmdD96W7ihp8oTknta++hzPh6xj+rABE4d8tZO3igXN4Iq/eGxFB3Tc+vVFgA
jh6sRcq4vBVmWuaDQJvohfyjWlNc9DrcyY0o9PGXusHmIjPYd/b1VtDVLa4BFzujKr191aIw1oPe
d+2w/hEOZHY7WxlqS3ZPhyreMNLxmT5IpQY3TGU+RZprEB/JesJyN+DuUMw/hpVBfmx+yWoGHHNc
AgYIsaJG+bcclhsbXX3+eQXT9q9EXXZrcep32VxMbz9114ttGOhnvW4ICkgLBX8HdCCPYIzU0J9I
TBoGKVmQ5d/tLpKd6R8qpuw3K53uucFvIbFekPD9IcfowP4/mhgp8HzMoKWgA8xJ/IDTHcejjIMf
U08Lb9j5D+W9UoEzFxCCbx1wHr0eBwOtKGEm3lchvJtXOsBTbWh5NpiurGOmKsOKSTdEa358qnal
j438McF5uXjTcPnTTbRK/TJciAWtblPXUWS47FcPk8Fu7gIEuxFSwtQoJ89JdWAl8raXEEPjb2cy
bU8qXh/dloG/79fhBUlJHGimQwglFZUQba4Zyubgn21BtqZsPnFiam8klAHHPvLXlkJDald7c/xw
ys5Ksv8Y2cjTEq8no6wQ2hMNEceOPi+hcWObyPfAEc2Gq3wBKob2gAcrpYBlHbRIY16TbsQ1WzJQ
sNoPLGKB/n2gtBeG1nOyaEzLXRDEDECB209+qgKWIFbPnXvhi3okQJL8RMnTynxW4PqxF+pFei4O
DWFy4D13LOUhWgjO2Qqvq8H+Q3g9Eq5Bj0dN7Twc1GVSlh+LBdTzYU6mR21+pH/thrm2jOKiLGTp
1CmEykmKzRS3g78Gtn74OfaFBQna5UHiIPswD/cVuIhERk7hzs8RpQwS1X371PrubSaCteLZSeki
7MOhUGxcmSfhhCEF9phKeOnvitPU3tFkZbXLfvKEaZgQaWeEA6e7UENxt6jkcoM4lfinpzNtTOjj
XPDVDKRNz/BdzXmnH0YKanQDeIjJUMEINY9Lu3wmkt3VozIvMFfUbinMmosW4n2V7g+A4ol1Gcj6
p0ep4773F5+Of0rcMNsuwlm7s6rKd5NRkSdlV25ItNk1NriqlefT38zo2VogPKxduNBIyEdxXXEv
UPiXJECPOb62Kqm5o6B6n433WMGDcZEaHoWrt+rbHpWuo79/lJ56SRkaxIWcOfs81YgYdiLUOK3K
aFcZgot2/CNJeo5myW5/KVx19VG9LTiHzl/c+0CyTafjcCAl9VIF0H9hdyU0BtVy2oRLrGlCbNQl
hrQ/CQvCT8VAJ4EUMm78+n16voBS9H2HBcGOLsv8hChWhKjRfMiGRGOouzal0KkR2ngd1Q//ADqO
rx+YwClr6lvdd+h6lCTgNGgbVOQcgQoVHF60Tze1CxGEqGBQ3vnKE+W3Hyj+NQbsSqnwcWK2v9Kk
gB9Ig2Z4D672mPgU82nvQhBFPkuyc9amQMhWHTORGW4uw6JudR0x0tBbvrAUvHfgDx94pbdmqkLa
dIRlV/47udNcEcqioiB42eqbtaMc633d21adqv7M+cVtT0+d3zfjMhLC/ADcoMWkjS57aO7bImdu
88FNFS/gl9MmiH/B+eg0y7Lfzmra82C1nKG2mftfXaC4peoFmE7UxsBJk70aEF5TF51MLiAMGn4N
kPo55cqhC0kedPdA1Gt3S/QqJI8fZ6NSHQv9ZS+67hX6xqakTC+5rCA2cuXpGU7CTncGRrOEiIJW
0AUaU/pqtaqOUjn8v/NuZI3ezPmqZKcc2vrW7vw8/CNvbFBX26Yl1ZFwpDH1QWgdRllKshErL8gz
CITwBBKRgDNlpbHir7NhG4gAwUXXoKAarDbD+wMttqPDIe7YM4TdL1crbJkVFDqK/07kF9u+W6A3
yIR0/mCxpwy3xb625RcmSDCeBFj6fXEGEhBHnK/f++ggPgmBJhTvDzCETdqr229hONg/YbVZvIZK
44ViVPlsexcvM2fLfotewt8FM+3PYCcc49+BQs0ke2k9AbVqKqA+/h6bICZGlKlBmOj0YA1Vn6Vy
lfQSkjf5VAiC6VkUZ45fIt+N+PzbJrkOj3Yeqoz51l5VboHMBqQrbwKog98X/G/kyWRHXnQD92SV
ghWVGm32pYhKoBD1A/Ak2K33PRuwPB53DU6gQ6BqFD+pV2UOb6/0eegBkNV5BDKLYO3Iac/PcQLc
2GgoZ3UREPdpTMRO0VLqrqbLlUyeP1z1/UUwrVqxws8bC6plkD7EdVAxIY5a7hDtamZ8Vj2UnUjr
vn5fp2akBwVVqlQMMkW2ujupi68FHJ8Yb/tOtlGxQSeONA1vfbXnXD7ht+kt4z70l+RGS+OMOGRc
vCL0BOZoWv/hNc44NwUlcR+0dWZF5LvFKFseiruAKMdyuzTuHeF6fWsQ8iFlBv+kCK+DtBeHimrD
qAk293SUA7yK0KK3uKu8EeJNo6MlUGa4KVgu/f++PePSrfpyCGhqBqh4Q9JrIbIMj4xpOjF92IaL
VdJt7dJwkUKuYWVPBepKQKw74v9cmRzvLWvSYpkJF4SxCkWE/hBc20KH2U28ktImsCKrCDftkdYs
xSS298+4GPfN6mSclrC+ju/WTepoXsqiGHzQm/oTKI1DTHa174uM5doxh9cgi0Xc7S8C3oFJ+DH5
ZSvmDkEWBJfz7WYqjMaO8gySZlIAqI1GZmfJwYz/IkTi9X2rByH1dPryOgxHIqwEaFJVEQ5l4xy3
YD2aUiumQiuP46EDSISToweaCxGr2eKJYox52slfvbYZPHKs/6rHsUhpIoBb/xo6GIaPzC3dkLF8
18b64SeF2iAOEXHPn+E0s8pEhd3bpOoTzG1B9u2ic5jznPcPDsnE/4ufjldjZ4TYbrgE3EnMe5vI
DNz9DaKWf60n1O7OgwHVKgOAK4AM2hEzhObQqWpwIuzPtxli9woEVJxqQEcDoeUMEDVjqK6nnamk
7HsCls5cEMBIV3U9yROqcm1hdyPaSpHAX94nmDtMIroqM8k9729G1Pfw0ZEef6Qk7eLQ0Ql0b+Nr
ycT2ZyRjwGFJYma5reD4DLYh6uTTxPEO+V4/qu9wgZFMhz8fySLQe4C1RiqSv231TBJisGhLUOPj
FVD+piXXyO12wrJMGKnxpTp77pPxLy+acwSExXmNfGF5gC6QOkhp651a+P1FwPsJX8DVtPQTVTm2
kfaK4j72qyGCOPbUMVMK4t3d3vdk/3f1rdVKv+vU9yvf07LqC9hP605HFhgw4RMCfRwWUTMSaEJl
k4ehV8NsylLs/aGgJT/RVwcPz7EXfLddTc6JKc3uH+rHKRgD23nRmZTrFiGOCQkltrYu3HJY5QZ3
vCIwO0LZAhXLpPcVCPqX5L5fyOtrWgAYasF75yodq2ej4vLMtCvNBAYho2qqlmiy0Nml9ALuiKz4
cCocCZvI5StvzFZ1KNHFu1AIy5p0L2z1tO5q8z8Wls1C0csRnJ6xiEZ2Qyk856LUjg/4x/V5yUDb
w7PM/E2d/coqw7XYFoHsS8fc6VESEGvwf8HULwkokoFWrOF64HXmJ794rgYAw4hyWMiqxF7K4I5T
0T8U7dAyTH9cU6k426HP/RUET68m73Sb2dncElGkPS/VdDVHKRdHqMpB7iBybh3i3CIAdhrWLuJ6
G76Vv1bCkzoRrVnZKe84L4cCLVxK5pzAF/MF8xjyeaY0ilMtRx45gWhQ1eXsFxsLLXaEILtAh+Z3
+H1XYFpXfQqt38tTRG0pLkUZ8l6fxcTbmY8h7uHKbjvwEvAfYOo2+DFf3YOn4tby8vXJ7e2pQnPg
HLaul6RiDILvBqXhI1gehh2FZ7q9W5K6GsE1cTGLP4rGcwkDrAQ02uNfLySTV1Y7G/J9sw5E1Asr
tMfH2NrQNf7hnpu2suhsDpemj5RPcSvs0r9XBctgiybB2zQ5XFd+TEy71lCwnCfJbwklYLR6y/ya
rLrKzlSYentnNTWqmdGx+ixhzCp7gg2F96ux7zOgzZOuzn5Jioz93JJSCoWdE1HXPhDxyHhG5HQR
yWKAlGZtI++z1fpGIFWQSaAE/GTVQ8aCDECY43ZwCHFhTZMR/aPCy9NCtoxkN85Bcu4fgD6h7B3s
EHbBtk7lP9dEjk34LBFmI5q3DPLTwmK37PzqvbfHnTMSMGyAH4WmBh2w1E4AV1u61qy+f/3tHXUb
2mL4miVClZn6fVrU+hz8m51psdpjIEpbcBloS+ckDVvlFDLz9s7yTm2sCPkguUFYsXdh4ZtlD3My
IQu+ht9Kvps3sYbclUW/0pzhMdIViG9XJFF92gIsrpgbEkhFdAnErZ/7zzmSPHftLXJ6VlKy9r+V
MW7sOR4hVnhUlN+U9WMww8gEIp75FXwBhpPH8oZB1wdbd8uOyXqHK1ronPkKp3ub5GmynFxmabx8
VdiMKpslM13OOsFqhvnIeDVp2eJjgMdRatrG7nzH/mPu271RazTHM5bdPH46+v2wmQLcIr6cxrAN
sT9juF2e96Sfa7f1mpm/bMbDXEOWwIfKnSS+0W9TPXh8vg1RL9GuhFtzMe0JN2vBaj6dDo0gMuQk
EbSTEvXZJ0HZW1ghKvUytvbftQ4xfxsCGYVgpngfaa+yes5OtLnfXTAdsQLA/L2rttynIEhER7lh
wHIMlmwgpb0mIq/pQDWmmNMtjdh45fH6eBlVrBT5UJbUsBMxRQLiQsdwl5zedsfnX3ozRiGtZLfx
vOBw2nMzCVoplp+QszK2EY6qiMOb9xzWc5r48bLJB4o3ofi/A+D2KzMsxCiscrPQrAQSDlYsqaRh
rzLGmk9L/nLzWwMnPMcsQEg5wLatpeQjnMsVnZ1BctnkfV89C93hiVboOlnwAOXz2jiSVrC+kQPt
7s/UAEloMGzOb1ZFNQbcMR44fxZCK5QLXbhzgYFhWWy0geZ2GnQ3JBIS9UvKIPQWsqcEkj8I+9zx
OXLIoC8Pnag6AT0dw0Lguf0eOO0MhmGQDLcYsKiuEqhy1wI+h31BHdgnUGLQBxV+kZIIwgDiaoHS
+ynlhdiHY77kZR7Ij4jvgj16lMzIz076amaCu0lJo7xAIxMq8QtzuUy4rftcXjy1DIaLdUbRJYpj
d3S2X1xxQpY73qAS3qVcop9Ibi9eiGCy07ulY7ABUo8OeWwRUuplZsUGykMsnzTnYbcqquEqCIHr
UuwUsqvq3b273enIEiyfJwnt+Wsmza9VZuBtCOBsuyEeHj6tuIBIK6LGARafCbjbjuUjVYTG6mUL
yAy1CZhZYM2BRZkGmZ2Staqi+qk87fYB7i3yfJG+AdpK4OieVGGT2sPT7kPZu3G/U4wlbEDzo2MH
D3lc13GqwdpvVzi1y7aKEbTZNtVssNuPIc764PufqfZsjPbJlfyyJ9gpuOQ1ACBWGy5LEnt/3jMG
SMMaOb65r6GKUz+hq3Rl/ubIFitql+x7RWwsAUg8GK+0Nk+W+zzJB+sAT6mLfHutO7DyXWSBFWW6
xxGi1XMkeHPgmUpk3PZYSQelhnUh7xWOkAtTSDRsd04TGwl9O88M0GLrqPBj6OBnjUfWKPKfQURj
Y64kxi+dxwP/59L37a7dp7+0Y00M/ZYNebrqb+bZ1i3EtfcAEVf1msAfoo9lK5D4BeErh/j3PjoN
GSEho8wb0n5qpSXZl1ORCS5ahWEOW4UqKqS3lwOOTctMHuSlerlIV0H3kZZ1+rcTXj+qCkP0E9Pc
0FIZxJD/Zolqjq/fXEd2KJ0xWToqtnCd8PGrgm25i/HdcpMnQD2BO13ErsjEWU8a3HDebRz9MJ3u
plx0EkMUydpG0FLLm+Q/GKJvl9Tge3pnCWHh02DJqkUJtbLCquNmxx1z0DqQzc149KSZ0iuBjHUo
+FwFyQuGA7B4k86MD+KTYETD5dn8rjtsSK7fUQWEIXqozBqovh38+tVYpWTHw/Xt77EnqOo00gWz
QzhJ+TIJkw17O27rdK9KUfJQgJjUcahn7oxu4I3Kkb7bZf6TZ242HCUUTi/BthVa6fCREmgGaGTT
3BnlR/fiJQxVV2BMnFizcIGA3B/BDVi2jxUJTW1MAE8+9Lc4zSWaAXTZQ3dTLYJHsysyalCjcxbt
H69a51bB/YjE7A1/ckGczonO0y6XxJEr39CAgCWaTARSUVxmt9Twlwj3Iq066NqxGj0ILNsS/crk
xKN6qxRtzzgV+gDDxZrxWEES40VtdvDQdBHLrHwBJ9EHxKeC3ltqg4op874gMBvZGgOT5c63Py8H
KwbDU3gCjQoTiOScYS4K1SSfC/yWrwcB8Q2RZ1G5BJsNuAtZvp0RK2vrksOnqz0sneKs+vNC1u5B
wMt++NkhphyqqbOJ/IX3yOd/Pb1yI0GpcjpG6zSqtn8I0i/X9mbby4kIr+4Ylu6ClQYvFfxd+8CS
5Gln7Coz7HgxpTkYdx+nTXkj1ziuRCjcezhbHhp0x/FETOhjYBWnbsKEM8PNpivZ7vGmRAwmqu9h
4KDZatEGBNgFfCJXvsoTpsH7tuGsPftJNHScZGo6ubkgB9C7/eyBUsewNacw7Mip2BnpnTWtNrt5
8EeQaMpZHlT4sYReW7EVZ1pghDY9MSuIFyMb8Ohp8+JRIUzon/KjH73Dr8uyXu0oFSNUFb3sZ7GD
gscA2rs/CWTuvoAs2hUmygwDKgFoOyxz9dhP3I7fTARiyz2a7b17FJZV5uShs+syXh10Ns8Y/IYH
U7lY4wttQn612JZFnRvMD2e4BxPkYy+OjLFigBwDOI+4rvhJhwwIS2rjRvlLjloIfj4ZUnGSO3DP
m/IJ4Xj3os175k26BRVa0TfyjcS3yrrx5mHKxfIZDLdxh0irK1tRKr9u2FVHbiIPIH5ISCapDQaS
3UJYggO//130SCQrxjJoP+36K1CoEkF/cUBs4sDHWum5z9BuczI6lwXs58V+9d1jLOD9/iU2SFkB
s/xbfHxLMQopOFUnhC1Ijof6fZOsDpNDwI+L7llQeCXnIo3LP5ivAAh2l+k8+OfkKP+iJ5vv/OvV
KolbM+cKp3R1AE1tsp9ip85CMsYdaupguOwHms5tYerYzFHimjrS+S+58Fot8HqvyXCUq0RWVbC0
fr74nm35A4lm9Rwx/rcdMP5lcIl9reZ9ny/O8iT45BvS8FrKPTUQdV1A8tnZwJu80y8tG1gKsek9
QyDPlZ9vib8tw7vlZbvqZlX4t1Hs7rgrC1FR3uGCZuEJk/JR9PcMkANCX/7MgJMEnLUJ081QKOUO
8olniDSHQGeIlmtEu/BoNDByj3/wIFY1IeNkfoz/GQF4a+mtaShKt2qvUbza1fgqELcNOTDFQiQk
XMbeAa9kI8s797jK8WSoc4k8t0cwqtAkmILWXwILFnuZcXQybqDdFZCO1G1d10nPVdwQg5TpW1ok
wJxBBtgvHPVffwgxW+6AklNqOE+QifrZw2tmegBqCqj7TWabSgMt8QcfYgg5TqnUoG9qBqzDC3Qj
bNj0ugwhDQXFXLzzY8UAx/xembxfYC6Zo3ypQtYlXX/nDvta1H6ulG64FIa8jZnlupZEL9Fq2HNd
u7w6A3j6iOHdtoAjkVLo8jGfTP0q0RMEWkXakL+dsFFLyMnxEDa28xuwn1q2NfANob5SgprWO7zV
E1Y2GmXirIbiC3G0bQQCsilZBUlE1ibB09uo3J1VPcaBJwfHWnuZydx521rkTM5f4zhKaq55oecO
9UECIsIO4eAVW2F75fbMRmM+WSW0EVuLojlSI0HAmAuJ0h1/nf3HTF3pheAhL+CfepkRbxOzx4tF
ZdlIHPuoqnx8xBWmnzF4+Ghjx8LhlY9HI4zhH+E+EVeGABgNJyP20pv0QSTOQdKnbR0LJ0zSwLz0
Dzw8D5JAxSKavdBQ2C6KyIepI53Tbk6iARZISou3Q3l1IkPBznakloJe8oMNYSkFjupv2K0ijgY2
4og5TUJ4w5hKkEwKPewi9nUWzMB4GXXYR4Uxwedh37XrpOOQyHCnbxSgzMog+BYLxIA+A/wCF7Le
mbV52TyC8Kvsp0zHG084ohnnLY+UqkO8L+9OLEJ9G17/y+Aj+uZxMn/iW5y3koBgMs+Z5NqqeZx9
6ZW0zoyXX0gugOq3Zd5TFL6fVSm8BPhoV0q0CIWqv24uQZgeQ33LDPofJlIs2IOjTgGgNVBE2jwx
YXMTU9InQB0dxCzSO/eatxcvcEPHI7c5VJqVdOXNH5uLYOmIiwFDsAjDf2oN4A0A3LFBiRgjwRgs
5PL3+3DBLU4jIsHxoHJgZsda/vom2QMnfaR5/UNYelcLZHLFQKetOYE+UKeXod2hDbrfiGi3fAoj
SHp3A3quKkxb4W92PpqCuvZucawHWGKs5Ox8wFblf+ElkHb9lvVnp9k0xKEqYiGGIJjjrifFtrV8
4AQxf7ScU1UBZafd1zmkdLV4RbDLrLg0cqxVgXt/TO/VtCmsyfMfVdRyCAc3s/d9Qe7GPXIfeYHm
MDewJu5WIDRQ+e5TItztHFyR8/Q8+nSNx0caIex1dkORe4wbelDXR5u+j4EZVhUjyXg26QlCz6nS
U1D1IUd0P03GVs1kjmKjn/1uOVcn6/oxLULEFn537gSbXU4fEJwc3FCAHUPLi8JVDCTqCCDbMHLw
+tDPdYbDXS5uBP5Zx8c0HrKk73nsPTFT46Z6uBfp9+FmfdXizBl74KcEnQ9tnJ7VyjWPAOmyeCuQ
BAVCma7sx1YbtE9gBmkSt58fLKw1Cofb74uUQJU2WVvzFcpxZ3uktleNmUUvyqUcDyggamyPy/cm
M0KbDpwTejMCfgeJ84AVd74xaNhlsWwmlMJs/PSTI9EwlUu91mYaVS+PFzBBtjhkgZ4kHD1b3KOJ
331wwHO+XSW01qSWvYyPnZmT7vlVZT2BWyROgIEY9Z+8pN7SijW/i8uRb8KmiBs+debUq6PesrRb
FL5NnJTQSta37hX8684RPwQRJ26KOXYw02yRkzqaNS4F7y50SffZL52MbqWx/MRYj6Xk1eZjedqv
NYWk3zGxT9ZREFK/HY1rtXtM5eVFaUHP6EbbZAoilER2lA0NSz5fQZIE9Vi6cn8ymv9At42Po4pT
23gWgWDpEwaoGmWKHeuUkyr5Bli3Za4ljzCP71gsCJUOgpBELXKaDd23rWhpsyMq4gLWrnagUNNh
OunPPuTdRg2h3bCQ/JUqaxOafO6YfygrvE8F+rxARrvF/MXVRAKuSyglZ5nTj7hviAPq7yYDlB3Z
hUcVqFaB+rflRHtqHm6P854LvxmH4vpIP85t2u8SYulEHE1CaH50B9D/S4tWIDB5Bd/RUfsOUFw5
Bn6TbVnqCXi3j/5/p1uQ/nIh9VSb4wf66ssPbdYEfgLrgDhQn4fqGINKnr7PCpumW/1dd10raQTn
qrWvCeq1/TbJ+LtX/3Qyij7mASpch6rXTEGxumam8ssaIkKVyDwhLo/ljL97Xifxjsv0p89pLcOt
WtjWs5wbvBcThv9YkKGkg4TErbwPg7PjNyPNCpKvE/goPQPItOhLHsm4Grgt6S6Ici4CAeoxvRkU
4QTiXhQbGIxFgoSCSwoLzT4ZMoY4CL2GGJ8n8zlAcgakjeV9Zc3aw4VFLJZEs8BPu1r/kH/qTjX2
TC+b4EICbXbyRJ1in6Wwcr2HzGYnEbiq2YbhgKEmnJ1VZJNTjDwIb4ZuS4PGv5RBD3DsG5kK9IsK
VFpb5V/5sPUAgm5XUREF//DAmuX0eyBp474a4et4xrlcYkKmf1DzDQzE9k7Y5SKH81EDXQRjFGRF
9+WVqj+EIm6QSBkI7ktYi5bGYb8NZwjk6+p9CkjDX55J9Btb6ZYFoPdT36zFGFi9QajUT/FNNMle
iX09urjq3Ij9BW+j7irARIg86tz/ByXa8jGBU2B5APMvXg1J4q7CfNRDCX3cngz0NKSghzVRc4di
2ozJn9ELMYVEJqicXOKMmKVIm5o++eXlSp3VZodAj2OdvpzRl42FFg70ouRnnaY+3JAmfcv4Jk5b
319aEzHZteOclqsOufWSUXDuGf/Kg45SFVoPGpf6yM7tYZvPLWpaebTEfqH9ac/w2r3owNlPZz6E
8qsnOwt4/FZXAPNl0gp/YDc6moTo631u6Jj0T1wlM/A5Bi44XQeNIPSGuRrDuamQnUfxBlrdPSOK
yRA8BTpRAuBm5iQzdAOXwOv1fFxZ/vRGYMCnkMe8w/QcGfXSLzLLIIRdTpR++aIfh5Ko/n9xetao
77ZmtMEKm+xeGTuNKM2qbeuVnxaHySeVMXJboIHeal0dKEZyDPmL8kj/2FFQnh0Miobr9zBEQcIL
zEMhI+eWtp+UHPkQNLGVbBCHNdCG+ULB+4Ph9+JojzXX5iBjVBIAP6fG6sKCSsRr0CStEkV9l31m
99+Cc7nXJCb+RpsRj/08B2PPrV7k9fiA+20wawcFKm3J6KTsEM63XfKk0JtXDWeBwo54sVRzEETc
Ae01JM6ynBpvGUdscVXEZoBMnh5qqUAYThChDmw60qV/QErgDYc6TwtK3FXotz8+/fDo4yrYJnmy
DoelKjPWPd9lGBZ4ZoXNBD9w895G/BvDTm3AfSvivI/V2WcY7qUcmm3GI6OqZVkjjHZrNZXjuJ1Y
heZaTbeQ4WBmLOCBeFBubAqr0qysIoZVGce/fcPD3rlFOUZA8pkHx+TWXzAQpIHIkqXBOQnms6in
ikF6JrW45l9G8UcX7bv3zkC9iHlDjVo/m9siHTvk2SQjkyICtZlfZGEkw6Se8akef4rp+LDSNGd4
ZM/hPwJM99Ih/SyLUdBjGpYqsEsjPziiEXejWFDYU+HajVCiYGEJ9HTaDd7DLehNu7nXWPlBZYIZ
EUe7yqHbv9uIkUuNmWLAlVTtaWBlSk25csOCB9MfixxYglfO5iAUaaWEQ0VNubg+j+JrcqvL96ms
WDgbm4WJS9Y5aTCREv/ybxdta53eVXskdl8k6LYUmkcpMlh42dJO6WsMpmjEZUXQgw+RP9aJCSeq
fJ8uH0QXWgTK8ZAD1VdVVt0ac5YKeAZVK+zJ3Om2phJ+XyR5+eHzI16OzeH1uSpC0StcLPCbGV4f
CqTDFCKq9TUjXuL5zNiV3bXrvZ59PqS0tK5H9bXMrFCkQ/SQBsY82swqpbm+L33odCaNx90Gvn9b
0YPhGILwsqCYQLtYYgqiPn/MMy6e/T5lBSKTbGuq1eUyyvSK6nS5CNWN80AWn8BMeSMqj7SG2sIP
CzswNT3M7lh19M9LknLmm88srUDj4nNO3ZOKlPad787cd/2xodGRrprwu2AErXaZKe1us1xXGT5s
/IHmfA7uhzlbVCmpI+emHbUHvU1mZwvXnOOaA2OIaxJ13zMzQvgYLdrSdf9OXa70Tat2yKXcWD4+
p0kH9C9s9gqCsHJ202+YsCT3RQf04EstarRSePG6ohv2DvWzfHBlnPhC1ml+aKnF+rXLKewS7vEf
1mEzt6+v6N7F/2n1BnA9+OYdTsUZVYhZyOVUiCzxc31fHyZEuYtkrHAZgehj6vG8BeEnb7KpTfBc
vjCo2MjU6dmT6++2WLX8ul23qCSvRAHGExY9yZ5SGg24fEMuCL4l5iF8rFzAbN3VkClOHE8QZP+x
Saxekctzd0zNzJNp8KLlP0jy87OM13WEkSEN+Y27yRP587FEc5QrW05sfqZeKe5wY6wfV7vyZgE7
IRdv1E2gXo9KPsgd0ks0pqhAuWNqTyLAZlUY3/1r2lS8Ehz/CMoBugpQhe4FZ1rJA0uZHQdwDN4M
zdf9fCvsBluZu6tNdEI6krptHoKxMpZF1hiQtnht0rlpU2vkmQKVLtaVRlZ4YUIAR2HCwB/24CKH
ieVkJCTczyGlQuU/ghW+Inma70ZkXSUnThL3DkkcsGV454OeAA7y4yAMlQYb75hdUj4PokuxpwQ2
JQfEPsm9rjnwZY55rENEPm42tSQaY7aNSTUcOePasSustCFB3uiQtOVkXE2UwEkX2/1Q6tsldD1p
6DuubfJ7RzCDHhui0hLNHoeZDWlmR5z9uNTcSsYYA3CCn7Ux2Aud+uwZDx/a23xI+qxcTdBPaJAd
Z/4KuWwtMymgnJqGoBbIaWJfej3Ow9zVuWQDNqCeLzgDWNIkPY0hvdo2cgaimSSbQQOP7UZcgwrw
wIqZYyi3MSR+1djcvbnSYtFw/hKYb9uiAFVAHu2Y5/U11IgiMJRKWstkXllOIzR/Ok/e9eulTV2L
lyGuDmV8Ybdf7wLBmVPABARoKMTM0QfphFP95r6myv2MUyRfBJww32tBgXPsy2XZKERjawbux4s1
61OCGYQ7sKd1KAC933CyLgkUgdb0k0R7xZapc+pcAUrXU8hpPsdXRpSlJ7VQpz/evLfPiLSGKcFM
lat/T2bOoLlhc8chZUSOfWWxt3+kEtw8ov74ELnm4MA27kt9PKCIPRwsApdBZTrPtmZjahWGP/0v
qVCN12UF6FN2P48wi7Qre2f6+rn5sDp+YFI5xv3CwciYFmaM39z4QzGmLHYREfAc60m99UGFbpyk
rLhQacHhlY/rSJFHKvtdjDVkPCfHm9TKiXdQPzErqGEGnCUaZnfS9XgG3E5KwGNnZApLwY1auUGC
/ADbOjLD+5WvHhFpOPPWxa0aOYvjYffIrjlrfA/U7fKNrEKmKqq3yVR3RMohaVteKcaCJB+Vwy2J
jIvN77TSkLXdwdxWSvoc9JsVBn+ByCNrraxZx0r2Xf3n1UwYo8aOs+3xobJc0r9uOKIDvCx5BwtT
1v8HZx0zi8zO44UaHrkpzZPMwmnkFnAmdGmbyRF0CsEqcUYy1WoDctj/6G09hL05gZ5SGX7glGSh
zlwlTNrdukovK18ZocTf3Ua+dmqJ4rgbvdOtJWwoBrB5XUCmlxI620iduNnjj/BO6wiESJcYuTM7
o2v/q5pKSh83zc5W/c2jzZ1JLD8zWEsIwXmedhYVR2RrjPoht/yY2Pt/nTXGIN8z8aA0AUY0FnnH
qJSt6f/C5G6ESmFKnXhwZbLlFtKHkQ5Zn9UW0tso6LOeciipGTRx36UTKyr4EKXRj25DcOwaC+vU
2MnbtAQpj7CcKpZSUEtECZskC8YstKvIOqQX4LnwEEknCXWM02y4e10RViD3htBjHkBu4rhO0AYT
NhfnELp+3X7zM7Fdy1F8iT+voiyMnlImSnRpvr1T9K3gm9G6yPrU4TUWkBEvY86dP5Z3/9GHbZGd
fJySAMVxcW8jAjRfih1OgD0xuCm6s8FDBmy5OuAc1mPjtksHBHShfImjaRxVpGdxqY1KgeFCQSw5
uWkujgRPmIEaw5UWu/sP4PugM/0BcYg4bKR4F9lL3Q0QIAPLm1qjiwTlbcvj/aC730zjnmTDJ/dq
OeimGuDKxflSwQCptaGzf3oWYtRRKcrv4M1cRgP4hm0bKQEM2Y0aFCv8e2VEz0vThKtxAxTztnp1
Ox4DI/c7NUdefo0vqHzQrBYe70Dvw668eVgxtAfbNDXJnSYhzRcLku/GiQaKk6dvnuiAmQRLZ4ag
n2WXdU+SxQQa73UzQwtmD2DCp3H2b7Sl5hjWFn5a7GsEnjaSqUXr/gEHKHKWQy8uCpwoSiT9ENVc
f5J+W469uAAZj/EFgOyuVopTaVz/UUv7hj9uVrlQ6a2c6TCksRFwg5BjQO2zpZuqtsaxx1Utb0M9
ERa/GHWG83kTMLj7/V408NIYi8cvGVdNhrkgCT7MmAAwzMj5LovCfJzhydAh6YEv/eJFM3fq3EsO
6K2MORB+GEsRx8Kr7SvuMfFhKMCJLVWiIqCVAsW8hDtjLAEmoNFn4ZH6WZlxc1O0fsIkVGZFs/Pl
LSCft6ePJiNuRhA6LJRbl9yrViIisrEbd6O1DNyWehMar+2zGiR5AK1ukOnRHJPJPGHizvlHi1Yl
6PoDbsaHwQTTE9GPU7fm8S7XK0vlv3gM/TlafYvjM9uJZxiG/ZR1A5aAmjWG8dcrf6xmGEQHXwan
5J2dZlPzFP6nvXKkwAKA+lRQg5s0huXaVvxEbVsCixTOKY0tHuwayEirHKATXojBaY7BMDdsufQy
gWZ06DRfjXNV3Oj3eeJ7Lr2R8qnWRYMr/6XMFwkHqGcqfYMMBp1/DjbW0lHAmc6Ws2UmYNDRjzv/
AVHUzRR5nLkbzPl3jH7+GBB9Jq2DCf0MtMLIRQlwf2DR1Fo9wmymNOvO0XKOViVKT5D2AWxjW3LG
rM//Y0yKwu5P8s6bJm+WHeq319DAgYHcObQxUuVcvQe1FQuc0/XIInuk/xhvEP7nct3TMcucbESk
+MuDHn4eBFaFbhwcABlpwJL/G7EwQgrGKMIZPa/ac9M2vZmpcGUqh+UzHIfbWQa2kV2HKgMDfTKz
RITJyvGh+hqvAFeCaF7JqZJz1ZBeexrAC9h95eUBWPf5vpHwEXeQB+CRIfR9UPVhlwwxQq/Z1yuS
eJBvF7WKAys+TvyjrIDrtdVG/VGJxugKk7W1DUXr70beWZUOXE8yUqMdSvOelgj0MhB1c/hzwtXE
MEzL2U29KX+AAV5m8Pk25lM1y5FHKPOw7/qzpoqDIvT+TMOp9Cuo5qqx03x+1gJxlbf7QV2ymaEJ
//FgQ1qinOdOCKJOnRePxZ+tOGJgmsLo9CyrbBFmhI+0aQJgcr3ug0syytM5DvXJoYcuvTrq/uDz
Yv3DFwhdk9zytCEhvhCWPntEBrgM48S1nv3hbO+wrxHBedvfv1BHvKGUO5/j83OlY3pxh3vnX5jO
MMFg/Oe7lER1vB/J5HfksovMTBhdqQzC+AUPbzbl68q3HwLHYL0dY5VLCg/XIwKTJsidXieEc+CG
gdzQ+Gnn4CBBFkZbRTciHVoqybntEUmDhDvNEGsPCB/kTtHZAeshIOpa6Jiw/rdrcH9j+2GOlhRA
vr4QaB7lSl0PGv/OWMVglabjKxX2QoNKu25rD1l3RY8/mrS43sDDHZLRGINOyYCIOF+817tLxGrp
3wz48Jn5ATypqhrlNuJ5BwoRF36LNngAa+io189hEzNi84U6oM38AGEWaGbXByhD1+xMZb8Wxs48
o79SS9UwxH1Om8N4iooPDzteFkw5vomFnuklpgotAzqaX+ByeO96tTLK68AoGEaJ9GZWewsamyRt
NKbDI/Od388MmgVEf58cJMuKgzBWm0AHnM411VdrBdw7ogCYp7+2HoDX80F46G8dX2Pz3+2CLD+l
dtfoQQk+SvQIorf1q0zjb5FB/lDpBzFB4pzfPtONLB2v+UuYS/XJnNG46PMQ5/2IpFNXZ9Q0TT+/
f9UvrICpSX8zIHFCO9sZRgUtm8TIV6Fk8yDWPhhzKUq7C+6fkrGFgfaDfj/7m2g9SOlULlPzZ+Q4
xbME9Hv4fEAE6TOJZJg80n6XIHzFM15y1jx2ej5IRSVa81fme0+B3YbTho4iDPQhLKsvHDXQlhmq
QlWX7CNBijSfNN6sejBIZH50ctacd6d2AGXiBScFHxBcL/1WbzDOVqjDYOAqK0p9PU5jiUUpod6h
rK6CRaaCbn6PznUsQ8UbToub9rxLdLfgjYZcT1Oz4AM6RQay6SQbGXpJcHoG51iOAGzDl2yJV1UO
l2h87BoqhWFGBGpR4QUb/vgarvVNtKzzgmCEHK1BYalV1YhkuWDnR2nzY2mARJZ+ZATWO4UmawbU
2dS16zNI5le/EsT0+SLXp/MdEX8cxplW8YIl/Bm7/BTXplY9ZIzeU6foAl5O9Ml8C1b8A4QX037D
x94vRgYdylRTKVOUqE7zbi7Czmsb1K2v7LD1B5bUYDSads2vAPSJUgViIbjDDj4JDzIMSK+XUYT7
1XyEvQ+9tWDB45kuS9AgS4ZoPbMlZcRl7k+SNCBzm8PGBvKgkpNaAD/Hq2d1g4h8QeLns04LOsdR
vfOVkO4e8+85nh+izAZ3sqPzq7szs/lKpWYFujE/SnOa8V9tfpxAjqfxYbOeUe5J0FJTkwR0iNOM
DchQO4gwWu0nG9aEaHDziNO735YdGuBhfKKzM1BmfRh0MBfIVksD7ckyqnFTvHJiRX4SYMZvCj3A
t/hiLW0VOjwMW3d2vG2qmBayzn2naQ+t27t/W2553w0J8OY6c+9YWd6oD1wcRU83TMeOZ9IFg2Tg
KgQoxNLOU9GLVP6+3tcrbgQfkCyv816BCNscXhtfIQl+y/CagJti4CwfMVC81lHH9KSQS5FZAV90
HgAO3fHD0qt5zde86w4eLw2JkRRKkWxTXjbmmfQlZR30wtzL65rJm/CwElkGMZQ/CAN27QaIRSJ6
MX4mT+NIPuNu37yycMKMRKIdPoNfjK0IOMSpScnW96UcW9+ZLeWukULNXxHRztaH7O8A9ZWjKbE6
AOL9CSLUJp0kAKQAB6e1YdvjLLwa0YqR+LnUbI6xe8fxE7Gdt+iH3kSkiqagjpaI7rFiuS+Cstsw
zTX2MZGZxKeiu5Hgm6DcZxHJRk8U/wm+2uSJW10uAPIOiW+zMtLSFpDBC1UTMNiq1OtjLI7Rx76N
MQKtl0keuHcKDgetP4M2Rj8Yo7wDLjthnTVJTdxVZ83sVg6j1r0gufZX0Q9Rbu9+HzjWvnz8wK5A
mahLLInI6zLcbqnXdajZXYCXnU2vD6/kUSjRxNuJfO94fOXAGb/WEEHwTAoMXrwR75ZmgIyA5Opj
1j/vaGlWLtCjstbaA1OAR3MLJ3POttS7VB/J7PXBf0AtVrhJxPj0hj51oKrxmfJz8qEoTwKmrxUM
s8lxOeVZViodLkatoXIk98iKSXYCKouxW5Kfp9x/LVWNWgQ21paWUGTrc5l5Jdiew/YRHhDvShuG
gd/iCI4tc4k02FTocHl5S63C75QZGhdCgmBG3C8Ng+OfiiyhNzCZLiE5x3234lnbp8TP9kNMkgqB
gyo6r8lBDoWZYv6zlb8OHksOSoowFgsq9DGdaZ+K8gH6+NY7iHNMbZZ+zvdORibs8LVuw+dXJRa1
bE0AQP7WIbN//N8gxAWbiBxo4Ei3G8LxhPNKQuuIUVlshZ4jmyovbh7xTT4kCpm3ZcFsD+gVY7KD
S12LKh1FjuaPUbSdrUqaHhPJz0OLaU7Fptdmck+R31qRWzNzTuIJaUH4E0x7m+3KOYgqp/VW3JFd
wSjGOqMfSdUlbnQvL0pjy2lqdf9fXEJCoS1Fl7nr5GhkxAXNp/hGDwqcNh/fW1N7dWMYs00dsMSu
4SvkxIf2yTIV1ckh67439sMV98Q8F/ffD9MmxotolB+k4t58+D/5uPluQSLB4xxSCJ0M88n5/hiS
xEebI/C/6tBbAAg2Vb+TIYqgoCY6bjI6MeoOYsExewZUHqp4ag/RG+e2t3UI+JBO7qofKK+VtEVB
YLmd3PZEYC58CJP/fpM3ialqzsQPtSA0xK4RscaDqNu9ItvEshR+OGrFjB5CaOXrI97RKlfgBoWs
FvVx9NWxivL5FUY/1bqE5PP+GEz4Rdz9AQEiTl2LOB3s2alQQg4kA+5ZSa+sCu/dSlfa7Q9rbofi
kyt9sHVQfmehlMNkiKSCaygat5/M3mq6TFAHoFwQOH0Oip07evMLnnbpumplTHgCa3v/4F2OBnGu
5C0PMXYRff00y/tpIrGb0CwkiuesHjf38iNSRjsrkoEd70VULFEMfrWxOiniW7DS6GTNF42jFSQt
e7aI6xS972r7WK0PWxkdn/Z3JB+jUXsnc0uKelhxs20R0dkjtB+LT7qFqCJenlguWRAwJLeUUITh
KwFM1B3qKvjeDQ3BcmhMXQPVFEeGemq766Lr6Of/z061PH8BCAzHD8TqS6lzi5vYWY6LSq5JC+Mu
arjJxsSHU+ODbHcxol66glwaHvx8ZdPFKlGYkDwDxh2z7em6NFU6JcAZysY/gT8LX/+5GuVA4Cne
QpFRGHeDIKW/bymIfeZEltQW3IZA0qXgz/ArRVLozXKbJwq8Wy8L4NJ7c14qoQAxmOyvWh1NcXxl
CPEp09nKIheM/rFoZnRhFT/K/OIqeO9kEJ39Bbwws+J2TInK8kvlW7r4EsqdAnzY6eZbXc9qUkBM
nr6xu1Tw5RL7kFfG61TFicTBnjJt3+eMVb49uGizrv8ghALgEWPg74d6yK6hYUuT4Rkv2q0GFH/w
RwVB/aw7zee7Vd9Kj+EMBCaq1ClTEh0ygLmeRrn/f4F3hiK+4D+gYcYTe9sgdrlTZVKBdq/P6lBT
XwhB0gyIt3USITYJq35ZxL5WuEVI5CT9PgguBeBLB3ohHR/OB6VawFuZdza7aCyZ1Q8Qj9zpXUeI
GRXwBGdtbwlHYuFHNpjJS9LrRKQeG+XJaZ/qFV36ByVsAJ7Q7wn0h6K/zKCmjkHxjABqYLyACzSP
ezwioq4we1/yFP+oZ5u0Y0iCJgPSsQ4zvwwDUMXX0jdKNfBg8XGzd0mOlbenwRKKUpqodmJQfBE6
QYL09JtyXgLnjmXr1gqCt4w3mw9+o0VZxk7ya30cxmMUNZsroq95ct4kpdL35VC//ESFU1UXwa/i
jBSnZRLtRhaI+auNLUyKr4OM1POM92MzESoC+TA1BNZ+YNWCSDEAClV8oSCoKgCwVmOSaCfk1U/t
MnWWqCKdDPw6W9ytxN3fqAY9oV8YI6Twr3BOGM+6I0eOwJXljDdV4DBFDwFwkf1Y6GN7P0D/6gmd
GvPem13gAMqAc21dMOQES4LgHQAcTNpor6Uk8B2RcrO+tpnzND9hw5czudyCA3LaEJw4KiOG5ZQA
f0QgKr0qJS9SJcFlFFtX4rhaaaPtXs2Zgg/MRy4RhJA7Yw0vSYeyP3GJjecW6PANQjRUq1PWWOSk
NqCnPhjtxkRSKcBYH3LUZsUl9rwuVtOvV+AyBQKn9saVS5qmNlWRkaWyKjTHqnV3WHvoX8mbDgdq
f02tRkW/OoyGCXbqJEEjKPLmsT1xXN9tjTgmRq3TZe+J/fK28ImDjs3XLThJdJ/Mf9uDVZ81PQw8
aLigSYQjGQG/cBgHva/01d7igIM59BZQZxcICf/mM1FnCmLK+bgaVbtOPIN9J15l+Ag/UBoCw/hf
fIODUqv3DF+/iufDH9L+FiTlV2wIBaXNvWd3IB7f2lunFZ2T+FssG/Wg6APFmTeWxeRQo1i/QU5b
Hvf13KH6lRvrjnCMezTxrvv+rXbSw5SQvbDvdvtZgkcJI8DCkEdqk/ne8erUm8apSefkj/ipeJ5/
Opwe9hIPifx1awyBXcwJRlYwlgPfuLmhx59sQblR0hIkd9h9QAXaGwK589T+a5au9U98AUq9ZAFf
dDWow5LWTQL2T/60aJ/SAr4pZ8PB1jbkppxrQ/BGGSeN5HSKVVJNtRfXrAgGVoT4n6DCvcTblDUD
+mMbwgwIXW4wLVm0vztN2MY6QMvYWDe9PP//OrQO4TKZ8PjUZRBlhPgWJImPyKRscGMLhweQl6QP
JNZKVVp83+bk1T0KRff1+IiA+HaMtxIrPdmPgUQ3MB9Fh+mmbzGKPGY2fZHiUU3g96CoQSVkll3p
SO9aLQGeF19xI0/NwzoqURL5HdmJr0ym1o2yFBH1osHaMOIucrGsLCwBLMQD58RI3bdQ1K6Yve1B
SwaqBHHvHMYEdNr2YPb02kdBF/1/OUW5hUwfMK++BWdwFty0D8kZ/tYooHZeMbEgiCtyG28bLCNc
iDh4y6rkY1sOH4VM8acSEZ6rI5otIud/PO2LS0D6uuiRVvkTSXZjNxZGMraXgQ2vtbycsUmx4WSz
jokYTaR1lE0z6AnqfsyHv1z6WQsvtqWXmdew0c4vi/7A5d+5GswZSj765rpGEgQBeBQRTG4Rvx1s
Umb+3XWnbT51NyHZUkjnN0nAmA9rjBwGpXTcFJxCV/QP8Uk9tzmE5SWZxpM5+bRQOI26M84/mazP
xWIwpu3C0WhJZDGtlZU5bLJF8vc19wRQNaAjRXue5RQXKCyv5hNB98cdF+cTfDjSm63bx+o4iu9j
8xd3Yyo3EnpK5xoZ7HuUduFD1oOjkS6In8kPLNhpQss893uB/9mKsLDsa8mr5D0nW/CaEW4Uv+OF
Cd+WCpGaNcRaFjMmQfC8MSW2e0bjpth4/PWu3W8r+Pnt/1e78fCMhp4LSSy9imyZgBbWh9xwl2F2
SQpEf1FQXypdMqAXw89OKC32E3OOLVHKMUVZURBaG8I3n68uVhxMaaVmPJY/mubaaB/n0xMIOEe8
58/tSdWB8X3Wa8n3/Y69CQuDrO4o4tPD5wyQjy/jU27jdD+Y4PkU5HJCjYMkeBEHNpexmw4HzL+7
gqdo+tmSWszFmY4tOOk28TFE2f/K/1lwTarI33sgmfIXx1AH8DcxJP9Kv1WdD08kOX7N2n8Dpw4I
+HagCBexynNoqHEYTG36Foo7V6rrQqtfTTjrqkj9lUniPMbp3ZBMQEZDTeqpOc1aWFA78rl/O2K9
pNHex+FFD7zUc4jttCnJckIALEBCxFkB5u4KiLYMrSjOoYcVx01RoYgekomGgLp6ruSpGqJEXZ1I
b1zpV7GXH/c9+/7MLwsJ/4djo3q5O02UT6s3AOsQpfEW685F/kqikF3VyFW9iBgK8yF24WR/wMol
GkMDxN91vu1N4meR4bFC7Nwn7QZ6TV4xJeDGRM22hmMNZnYygxp3P2+Eds3eLQsaBfitnc8+0y4p
L234v/JRgAquZ1kOQ0nK5YpVCYytW83CPjT/GObIcSamRuOs49jgStbskcXc6dVMVuQmFBYwjgA1
aoBft82LnkuGAaFgJvRnyv8Ufej3pcOGWGIO4fll4CrsygWLyIQm6kfAYeHTXrEhV9RGbsRoVybh
ArLjl4Xy+rt6JsWOprBd/6ZQ/H15PZqvO1Aw/YQ6mpF6d2iaZNedJEuSI628VyEP+CIMpM6En+Ik
liXSUI9uJFaOWo/dFgABb/s1yxGL3JTuJb7lipUW1iPDoKP+rZnjdagOPhL3FO7ADhaSarspZ4JT
GA8+iQiPAgFGe5vU2sCndGLM2tiz0Y6L0nIclSS0LufdAyiIenPXI8Yn6VrbGEFRuHpQd/qROazs
hyd9IYV7u3VKKKUQo+IrgPW1ZK16qYFRPcfxne/65qmT3qDdvec/fj1M2oB6ACnddy8+PsaQVZdM
eWGVhAU0Yg0P3DTtmh4pBHED6YGdtwMkKziOZbMOuIeaupYXgQw3Vl+WmbFK8X3yUVbYjmgQiBKu
HlHum9NmA6GEflw+ltepZIuSTrLMPwLaD8QFttqPhO+YUJMxSnC64p6Qs++ABffjdLAAUZUZKvK5
fQcyXlNhj1PLGry/C8O8ygtICZRiCN8Mlj6qjKsmMNpiRYhe33DzXCPyfgqTpF9V+H+6aRGah0Uu
FIwgqiV0JOnFiVBlAo7KsctcDMOraMQ6L4UMTRS8MsXrKzerRwDUgBn3iRJpS6SPK2+uD+F6CCmw
DDs8xbpGFQhTyJaps9FvBZ+MjtJZ7c/TmpMGZSrVdsbuqNQOGhHYrekoyZ5JfN61gXwyn68JWBIu
ODEJWRXoS9PpUCVE0VbrE9dwNLc2WE1VRbgC8H3ULEyEAv97HHMji8hlLNRE1f9M+NCuv2f5QTks
F6B6qPW4+SSjSG/IKu0c0kflp1WuutG9nZM6ZPn9gU2lrIdKClPttwd6qzZrUEi0BkG0iW5brzXq
SWJZcF/AQE664sevXTXTzU25IjyGukD0y0ryXNRA2O/k3foK7VsFZ2fMglhLfHaui+S7peT2soc0
6Q1KW6iKiTjYGFwpEbTMUppBOlAVV/rKZ1lTubZ1ulNdyy4QSlmnck5gENRYDxSOdOGIgxALGln8
4XYGGAYypyWrU+tQAeTSY3u95MHPM3fOvDea2VESt0Ko2GrUZvaeQ/BfcD6MTjzOel3iYeDlgkbb
RPB3z4VGIPhMWn6+xlQjdVflGYP97AziX67K5VALVAQeUKTUbpe4Dj81ygunDpqKkvSqGYycvZCM
Owqv8tN5SmL8cEgxGAv4RSfD7Z9w5O0eNK10m6W8VJ+dhyDCukjTI+aQCgsmmoHQB1utuXUgyxuF
lMxjl7ktEgG9JinSoAyxJViCAW3JTNtlKhvfUi7WNMgnDZpGSPYjPlKmsZoUlCL92SU2T69HeNth
i02QWWlMiCI0lXIx3XI4Hocdl8uG9IH9pVD2BbVDDuR5z+p36Z3hZwfX8Vq/wS11wSGsLhbcTpcM
NI3A6luasRsjiJkvs+RnPtcw54DqF8J3LmukTxajJ93cAyBu7rJv/bf4SpckGuam+76Kjf1Kw5+3
WVlmDdcP+LIdYIreXBoUDf1+yDweWkEn3CkW/Zh7C8oijAfkUg06CXY+4trt4j94OXDDxfJyPoEG
cPwRAleLS6VZ5Gv62OdiJYxjRJukFRtbVAK3AASbS1yMBCU2kjr1EecdajhmIquhOMz5NcQJmedl
AcRzr0fwKOHZf8altjK3k58EC8Qj/PS+h6wfjAw7cu863W5k/pDz+xxxU+LVhxThdYv8a9tgVqUe
LVcFzJUL38GDGEXgdYtYpXAvyNR7knPlpgVgjaLn19tJFtv4DE0TzxlbFDgkXo5kPbmM/sEfMZRf
F9jRDLM3K3fN+otOz/QGZGAQrAKioV04qBA9kjsYD4rLfHl2bS05Klt8VuaI5C1vvrn14uwtOl8r
30UsxAbKVDEDeL0ikxQT1VJD/ONcAsTrcPJtBVCM3WrFNEWU7EHiAS/7qpZKtBIeFFQxRslp6F7L
tXRsUvmbiQKvuU1PLXQyW/ec461KY6rfTfIPV2kFArURSTrSbKfnXWs4rRw4IJs2vArFDvWMwSmr
qGOFD20KisaLY+YDnAC+j2mxs2mkDAg3ySmd46OPXoUy7FjQVi8uFji4JwKjswOobNe8rEpf47Zr
M8y5iuFInbLlYaVbqyWpYptb7hj131OFAymP3SuxbCpi8V75Vj5b/w9F6H+QrFMw7O1tNUWtNjuY
TyyMHl0D0hMa9jD7sDU+b/qBwPdvyR1LnyXopo092hwboePvdNMiL9MPsLTo0VYJ6KLUa9sd43gL
uKNADVX7KNK5l+Gnw8gnKCp4+Xq72lNKBrW/juh73+o93XBJUOMyL8/4oSW5xCbgq59TSWPmRcRV
P5r/MeVm53EIJ2uYu8IHGlY/gbqQv/tuil6+9tKzXqVFCoQYjBlF8FQKSEFUkCbuKvqb4CRacy/d
vYR8gGR9v2y1RArDygQL1mXwES3RE8JoKTfqWVdU7pHN0Y5kDbjCcg/E+tlAhFJVxI1is0+//2TD
aSRmkFIIb4nN+F1VOe+auB18uOWcMsBSHw5RHduUJ9NAUCVmILOkb+kmagiAL8jWqNpIsMQy8goG
WqIjf1rjioiunqFhWk/LlbTMSoz8VpzAUUu6G00FOlvz+oSQ3kEloJK6q9PnxHN2jpdEVae0Sw6N
aqdTefzmIa3f7tisUrw0c8Xgq5SXcpagZCiBdCy0Ux3czaWdLA/rU7kwLtkKVC4ZV67A+ZvnPTRN
o6+9tgK20AmCqGfvHRXlfUAbszS3HHkIyKsDol43s86dg2VD/DchxWMTgfVXX2s4cpKeBPRg7R2+
jK8/IcZD7/dfSgpVgfsIUJCckxOO8qyOUOH431GwinqK3+DU22FuugTJTtcLnx/BgEHc4RmK0jje
YUkDiRbarQa+zEGRhzet/bk69tVfzzhEvxKvipnxJ/Ue84Sch4jO8qF1SwhGjQW664D8rtjig4yN
4sleTeZ/63+NQhPSKC6F27IHD/fR6Jmui/6xt9GznhUHPVwJaMIpf77e+8aWaqSmDZ5pwtkj/77D
kuN3MKu9bbGQaiuDm3QlLvlyPAaknjjv+zLeJW5PQBW7vB1IC5WBoyfmwV9D3CewdALi4amojNfw
C+/oR4SlrLyWYA+JUZVKfmfRF11TXNPofjV5DcG+jIBin9YxCndcDO7xxwA+0/AKR3k7+L6I8oXR
m1vpIig7yj5vF5cVCKKPg3ZyeEd06A131RFCF2lso8pFIzF8/Gv94HmIBJ95iMaYArp1L6K+Tne3
0cAAe94jQ7FD2sQJGFXF/3DCKmuLfoKoHyNX/9cYuoFlhJjuX842Rlc7ycA8PPOgmcGadUbkljTL
x9sZvTzUtoUxyVAiuQWxoh7EJrawR4PcqaloTIs/rk6zK8XUGz0ROgPohIFt0pPnG0DWzDEb8PYa
pbVOkIOU+a6sAshM2hNm5LQSRdbi3PVZWDUewzwjxqA84CqBzQ6fMi/RxJsmPBPpCKteotSwuk3d
zNvvenLY/+Vja9vnnxKU/d9dFBp05gEGslH44WRnBnD0+BWObNdePRxbQ4al2UY1t6yCBef8/t7E
N4msEM4cYDqOIfNAKSOwz28QoP7x1D7H9DwPXaIuM7uzS1CvMUYNHUKs7sHzCcWZXvibVS/I6JX8
SYJbvftQPsMI+evOXfxrhzcWGY/Jnp5RgNcTDr/806hwJnnMZ/AnDtYl716ZzuyEzO0K2gXRzyNk
7kbJ2KS4QmZr9g2Wp8XI1flQR6P5BAU4a/ydcALSOq/csUMmGY4wJHTGwcynTXeFuX7ihu98ysfJ
5fm1IDXhTzCAh2qzRoJ9+ocxW1RWd0Cy52c0fGKY2OiyQ00PR0iwG0u3sbZIiv6CWeTfMvMl6Y5o
lyqx2QflZxVjaF8Mfl2N7rdIS8nFF/W/N6Wj4sChTmX21MbNaOMqOlKMsVJtEHqV0olncbkqcKix
uOKTWnVA1Oed7I8GRDszR5K51fYzZpgy5bgUlWh99HiHvsWUWIDVVMAhEIeTZWJuJaJPk4wDJ0dS
xpB9WjAP3N9Tl1Sol6Zshfc4xdanIUd5orca40HH2WQqkSvCQJPYsjm5G7h6Jt1MbkpnSnIXppXN
DmzhZCRSei/WIJOTqPZvqR4f5vsS/MG1vHs2UeCSaqjiyZhgu4i2hUgC+uRIwNKjClq/CEx5ErGQ
rvQt0fpS+CZ98kKTA1o8RFuwqwbi3UWceif6oqjqQfYSgQFJDHPYn3WjsGzP0IXmNZmdpqBPolQJ
C/nwIhHsWS6lknNIkUqPR8Vo9DlOc5QzXJGRQ14lqVNVeM7H0B88E/2rEyoj5JKDXyPbeuVrPB1Y
e+7TPHVMW5TevkQBVD2Jg7GL/pg8wIiIoOnLGGpZrNKRiep/FnKVJ+EH4i/kgPmnzzACDXJeczOt
YAe4JHHsI28cYADJTsKxwT71UlQKhd8t66dohukLq16v3f+g+yMFjMWGOGl1C03cYFKawOJ8vkCU
r8tXzHYP5p8wFXZT7xo1r+Y7zHq1G4qAqAA0XKRgj/OyQ+ygoxMr+jIRCPMoHf4zFpHvw9GDsNiI
2eDIYeV6mfWMUYPAn0jYMgET6bSXNher4eJVDVRrXf7YEgN0a1MEC4Lnunnl1M4rPwtflNTrv0tF
wa8I1oBUSgFBoDhiCpSFMs3IPhPx5ueXH2qGRamseb+xYM9aso9VPcw/qDLGSFaqNe+NRs5vFKv0
EvxodGeehrq0LR9BFCmv/Mew2BnVvO4oQ22wpRKLoMLOmJrO7YurWQ8JvOR1BG3ECdzDdh8MSCCT
podZk5z253eBvVHtzGs0zqYt1QDaCuXNuQh9QKh4JexG4int/Sx09CDu89/prNaaGj3PeLnDhrzp
n17WgKeTHL25tWj74Rhjo6d0IJllBPpRnAhfzagLalEcEStT5IiwHBtmhsAbjqXrc6xm3eTDhszt
6e6vkzVPaISR7JQE7gSa3cOU1XDvInLL9ICgk/b39F5ywhj397UEZa6Pmn7bLk19dpAZdwfAfLvq
UmwrLD/spv4OCJHXDBmLlrHAIqdh2deL9l1T6DcOahyJfofLskOBSHdJAtCz8T3yJK556H3G/btg
edQQDKb0ublKd40MbKYm5SoBYda8bjjZw8eaglysU+5zwbBKfYJSS9sk3Xlh+irpN+YHoYGAB1PF
JS86VoiAvoqNf82Fa95D9BW56bD7w4WiYbSD40GRKsxQLUC3+ihGhzbCUo8I++N7obT+fz1YuKiy
t5qvUD0AVEUZqxMZEuXwVl2ztkEEr1sReCJFAawrJfDbuJe4jWjTPt3LoCwY2UnCqhKcYaJhXs7d
sUJlCYrGuxZJiuQ5c3BS8i/O4xRneKePLTpGMi0BZQSvgyW0z3D2PDQfF2UX4a8/vZH0uuI3jXyM
Jv1UDEfkHBDwoHWTpykM5acRs2JbO2+GyjOzb/bzXQ0hmY8QgZYTU+pntM1lS9LTFOBgRPfOQSDz
D8KWZIbmA3Z6HVZygevIT5WyAWTPXPuTs27jIkw/+hjd8GHXxkodLmvbCuaLCoR0+hbfvlaZmIZo
3PNE9/Idm8uhR0FjWywVJcGvO7MrZkIAqQshDq0zQ3SbnAZ5G9TFdpCqfeBwBWcnf2xnvMFtpu8y
ERCxOhB4lbzocKmUNp6BWT08R6l27c+vlahhMFPbnxiJrst7iI4sHAq3j+B70Iwab0vM/J9Wzolv
qY86z816Kp8MHteTSVCIuiuYf/S0xrE7yWKD3u3f1DPOuuzLm4N3LQngHgb4e0EFu3aP+t6KtJPN
oA2TrA/7cbSQ4gbORexTGasIFlkyyRwIwJV47EVthRg/tKO4oX+KLfd7xdbKl3wyq+kANoeEmQPY
B+460cUIR7EC6wr7Uz+4OQ+vfociq4GILKyPuKiMdnRRzoY0gAUttfWaPJyLhEa2tn1opt3YRcOC
l5oQre0Lh9KR6jESV05453tm3QE9V68dT960OIhFivUXShVCIHigO6PIIGMX/9XXZPB21w32ykUb
MFR26VXhVd+z0cUPZpDNGk6Z+DkTebkebFO8PeVT/AC4JdF8/mtBjWWWjYRzgbssXpeyce5uFlJ+
b6yFKN+dHulbGh+158ejRM004yB7jH+oriLHEH4Wj9Xx+mg7ZZS+4ZPJvCfgHV5/IeNzOljCBaQC
3Z+7Q6RSpdJPQefpw5ce3qAzllwcgpUelQ6vd2y3+kNaeaTyD7Q1zKfNxS/1PsbbgVIgC4S40D8i
maj8yIYQSfkWeIB8zMJMwyfdQ/k+E9TL8yjfL4+WBIi8phAJ3C+l5gYaM6igMpqcx2zn+HG8J+x8
+BeXG1bkuLBhnqayAErz1X8KYkkzYbzohPBAVKabYmS+a7rVySj34Xn6gkvHYuf21rWcwkg9acxp
U0Auk7B24igYFF8FfaIpLigCxxk21M4aOWhyfFb6rpJRhfQ5SIKHlQDC48v6zJQU0vIUa28rjucI
JguTN+lagQpq10NBAlMIOZ9BXzaDfPlKnRnDAFxFRCqxDm1795/Q6zCeKTx+n1a60B/C2tqWBaQV
E4eZgYNBIS/2B7/cfgW4BvO2EKScrFB4DgRNTQZSEnYhmBjJbjCTN5hpz5AZN70O0xop+Nz2WkuX
/Pg46ENx7+/PY4OxDHUttx+y2RjYpFVaih9wkIDSHMHZYomwThGa8KbPeqIMGbs7Uw3U6gX+b22Q
wVkmkLJiWch1ZMkaki5BD8k/dxp4YFnv8Xo8MC6a8Em3bz9JUzhRo6f3H1fii7HulVM7clwoHHT5
jfumxde8xeimkyqTWkLhdr8Yyst8x1pTKX4TOWElOgOtk/iDs/85JifL7sCOjt5TQMkI68Kfq13l
KcloxPDD9e7l29pib72Qbl65xcNEVsYdEeIU4LJLi5oH6pDogdytvau3E/ndY7IeQnJtkN1KQ5Pm
ixl31GzGS5mJqscq+VSmPGYwz9YBX8y3leivgPmnu5DmxHIw36dUJvH34/1c8B1GXstBsnrKqkyh
R5gHeZXSYjYWOhAp3mrT/CaKEUW6zm6c9+2xN1xz+3f64stnQkxaX82AR82mUhsqRR4dnVSq8T5A
HJY32ThkJ2iel6VF3Qm4NErILS1YddH5R6TVEzc3Geg92k3TtXzNJFuMtIB565YTzn7owxl3SMsn
Hb7XEUMCPcV0ps3+SwQDJgS/lWF9VrQODu6EqGBFHyY6huLgQw+1HSqtY0yBYMqe1ViDKhvkn0Z5
B22P8NKFEQoZJzwCEoipjmneLtMRtaMWVnjl4d/XgXhE7Zlg++55H/3DAe4fVtRe0HamPTBOzVxW
6UrAO+k9XF8/MhrISOJR+kMsJjwc/nDRtw13oLMaDsTpnFbeqZeDIlWoJQPqEC4iaZ92+MLkWVKM
VUT21u9C7KjQFGHWyqhpo3sQgFHiK2d4PDE3a1h5wz4LC7g9p+V5qiV1mY+24IBd0QueBtiiBIaY
A0k8jIdIoP4VedDCuqqpGBBp73/mrQrrKmYXb99vusoAsKWMH8kt5TLSg9VYzcwSaes51Ye/aP5a
Lx7zpSlvgh8kunUDvMe40ZD2/6DwBkDwFunsOZwHldywNO/gczrm+flLTRLG1MA9rRprPdAk1un4
s56Hc6qtLF2CazG57vJcYeQyJjrs15u9PpC/bUMrN3gX6e4fNukkyEBL1jxhtowPOxMUWD+4d4bX
7mPcQ/VpQbUgMtPpUwo/MEvNgJH9iew+8e1zMqsMhkq1uQg8AvrVfZljzX+Z8NDuNGyQaLBMWMUy
Ri1/l6WrcF2pdjjtZGYhw4/oaudn+Z1qf50LB3//qC4vCEpc70HHKmlCkuszDDz+AQpoWy0cB6iX
me394Xu/R7RRUZPGduQZGkVawMhbkLnP1V99rX9mIs21Hg09eG5estffXuoka+6ZzW9DGdZdyB8A
c6YRzH+gCt3gqP8FFPD+S8WWmMhN44dnnNCNvZ+bJeTDprGWXzDc2mugjAZ/gPWaanfTi38B349o
81SSeFBYIB5YNtn00TwTn80sjBokqXJJWAeZqRI3+TKgPjeg9Y5F2h1YTotqWpNuVxe0Gi+KBrQ9
TNrAN/DiZzFLeDKMkWe2m+7QpgBffk5mzbK+4CIDqxkvflHYYf7U0/1se43pK3iYWIUZ1R9r9kAS
jlCBYGPQbcLW3CW1iYcURn8T+9Q0KZjvoLIu++3f3GMUyUorMzkjFtEqLJ2AJ8UUN3mK2mYV0fU1
XwyA3E0UpP2gTKpGSydfrsBa/r517tV8nIxQcUNvPUbh3m0jvp1lEDCY/hfG3TOTpRBKwgz3/5oB
h7TDiC4LibZ+FO3lX5/N164oubPu7uFmsoyNtc99uzyT4zohZ/xbzTnldq+aU8JKYZk0ZaOZ/6BW
/Qjeu+qrbodJ2uP3qyM3HIxFPoHLWtfEfIjt8O0RUKwAaUM5C7WS1K0qe01W3uoQZnmIyUrGSeYR
e+r3clpuwwhWELWrFJR9bmGu9IMg6grYt/76V+c36wjnAcYvS4pCZp8tTnjqMl0cVu8hepZ/iDyL
d1cj9chS6UscAFer1Ke2kZWh2w9ex1qAWYo0j63R3LJZehXWKj6ELMAXCzQJPkIJHwautjxe3+4V
ABIZRugFIz35voIPGuDoa5ha5Kj7CfoZTZWia53x6Z+RjF/2jfkgnITT5fBlQzQg6GyNF4YbF2RT
qu1jlXzxxQO6f8bH6lgujrkixRem57RKu9hWKnlPL4FpOVMMIYp5BzfbJeOsIfWNo1Q4IMuGSXJh
brqRbzBuYEVDRwJDf9OeaflatLxYv+ypQoQnB3Ft9J0aNUmqm6eID6o2kPA5QwBm/iD0TtBKuTUg
IA8K31CWljecD8Kh72teoaH6BIQHr1qzYN3LxcvISgtFwF0I17oSU7cCGMHNMTnGx4UcVS5x6ptZ
SsXTr2pIiO+FHm57F1O21OW1ACBTVpcIFUFwXOWY46pNk4mxRR7fXPuHULwv+tQUyi1TDS3MHBxI
U4XCK0yjj46TUUnFvtacJ/IWJl/SkOjAfZATdPY20IItcGtsVu8r59CL/Zh1cztRWFG73FAUtOrH
XQE0xdXqmQbs2NUADOSKG5EO2LWIGDLsy15Lpyc2OrNVxslS62wLlngBZ8pwBNE4R/9RtY5TlVlW
dEYytSjenZY0UwpgKbc02cg0yFGVOqvIhvtLH2oEu7BVe9bcorQ/6u/osPUSdWATwGWi5AWMtAMP
h4lobKhkxnxpMZf+9V/wTRumIacGfQ6JupqxF31vbAT+ibcsqO9EjTaCs6Mxrrph00+b/O3U0QcM
j5ixbbjZCUDMNQwWR3AG36sNJoc2QaHleBZmG+aZe1GZhsv767ta8wUEyqegqYgFsRxrRRtkPpwC
Lc+jpc+UAiYG91AWdk/d7+bvVrZxj7Co20kvQz5lCMxXDZ6I0wBmgvkvjn3DQxkfwCxF9s+8gUCI
65uOnbysTZz7Kz4g8ESkYtf3q8Lhf2aTR38/dsC/xCG3HD6cMSA2kaqtXGheDu+BXcUMJ+iove96
qf0cn0x2N7me7FXDLn1TcphmQ6BzdWhjuazrf7ri/Kt7zKWuNbwgxVCNnCh1sVNo4QXjLcgAqQS+
PFRuVX0GscTuIO4q/VLLokEh+FdjyxndL9JfvioySesx56FnenIBY1BpGsbM7IVc6blVqr7OmCkh
Wp1AdwxQyO9SuxY+KjpI8r3M6jdYBBEWG/S3S/qajMA8mv34JjInCS4bH9iPuVkb9DxY5B2cNHuD
psA2Lf/P/ARkASyLf9Ld73M3mgI8qijwGyWyYak3MJg00QuLmonUepJWA3GvUaGmTvlZ+cL7tKaD
EbG9aMmXCy1qOVwZrZF1AhIr24ZkhklWIi0Nc9tsXd5qU9ihTMbyo9MG+pC67fBFLmiJL2lVg0Lq
jKZ6Pw+49F3YjlrnzbWViWEdFgTs7f4FAvcOxtIHtJvp11GFUQiWGvkm44BkDxKgOr6U4U4aVQ0s
OxpGiGhXxYAR7JZv5Rf5beEsyRyTI6NMbLiBT+GqBQDGaOs2MH/Huo/CirvjsoPO8Jh2XXyQ4dhI
DK2Cig8iJBgODPJBjY/jDSsMV0T5uUOGUAeAFhb1fhNdTqlC7K1Pjvm/LvxeHepqlkInS9qyiS+e
pc8KY44V1OOOSGTCCdSvaxAgdEGlCnUHPV9beC8XddGmSNHvzyIGgp3NB3A2Ndn5MMu666+I4QwU
5Q0EB4NzWiAGR7piiR5oMekiiv52CHCrZ451pDl0zg1KpiG4fko1iTSH1nL9UKkrcMxN2KqECR0V
EuuPH/3pAe40HwQlFKtrlz+KNiBA7w0ntll9j2vrNuLv+9lpCdwfBxCUXF7HUWFtHKiBtzYCUb4/
eARjvDdrXFUjWls3zLDWNlHINT1DBhKOd14zAR8tG/wr3Pq/VQHvlOsuUWm6+cpiBrkt2CTtN82+
WAa7mj7vUZT7A5wtGegpQBD1noAV4b5Sj0aHMOffiZqlOgjx69zpQ9i2sEc1VhLvB9oeWL3kwZiW
hM+NK1gHx70t7RNCQm8e1kwI8U1zUyx1EhRL8P/FD/GM5FmXNLb2nMuIGsgDx+E/DDgzoHyrKvO5
dYpGUPf8Iaawb+UYnzDbr2r9HqrdEblfZCRKsx3vRohqzy3I7l5ql2XmNrsExc88Juh5KM9L61Ju
2gjr84zUWqOi3dR+MvMquxpasDZZf+jrW0C/x4I3al6Yc/Lc8Iqw9J+4kYTi+iUk3Pb+rKqBv65k
jbrTjQk1nHjiPHzTmkZh4y9RuPUbno22nW5uThHLMa+/eNn4sKkN3/jgEgchd41rHM+VWPro8Zg7
pQDmmp5E2JQQvGufaO5ZQwNo5psC4PyQ1ccp7OSlgIp+hBeB/e87CAii1H2bPi0caUouTOVvewB8
EWmzM7EIe7j7vChKZZRV9Ft4JzCxKfd4o54MafjE4ptLNKs40fwhfl96z1cj0pSvFfzf5bkQ3HW7
booMHPjD3SO9rgdB2CUDrnsLytD+VW1TyvJCToTQYgXONqOWZxlD9uOb8wu1qZHEjjqxjWiL9gog
11UHzoJKa8YurB+Ekv/v2A9kr8Jc0SaE739QJ/UP/C+VpkMLoVjI7L37N7NuRX86s761YUvUJifr
PuCIFDDKAw7FKubFaoTGP2PYlVdhbEH4DSfOEC3KlKCdi2Dzm5DxFKAuRADRbnwjF6y9wfy03pIS
W9Y0kp16PvZ2Xs3nrguM+OiYOKJfVRooFGS0rvnvXtT21jzPTagioCK43iBQhtldH/h7Acz5o7j/
GapYRJYDyq9D9TwcuaQtXB6bD3+jNGcgJ42wL7CDM/giu805v04sXFFBKJ3IXACzfnC1Pb31/YD/
ESoOPxAjOIjsvZ5CirNknlXeT/J6GB8oPy2Tm8AbXUODopuC0X1w5YgYENvZN5DlQx2QbyWjlp1n
jO9uxAw0qoksyznzOJBPEnJwbqCoJfXH1GFiHFvs6z8PH1cKaUjzTsphNSOzpPIfzAmphzY+rbdt
nMB6Mnnlf9qy/6w53JhCFGEaWQlcC5zfG4IM5wqWVatsmLao/Kk4SZW/0WXtdI/O7teMkujBLGc6
N9QQdaGU+KI3iTYb3IJvnpY9qsNIPF4lv92jovuN+MSsJkHc6Uh9wk5O8ODGTG8tyiI4aZqYdDRN
ABnh1wgYcVuK3/GWYeTfzONFoRvvdGgt3Y7/wsq1Fxb1SMk4HO2Me+YDByKq3Hf2IBztu1DVrxWo
kgJZFCqSyGKmtnlYYq82weoeB51hMczL+tBQVMN38aAhwcvTVcNz6XYljBg7hE9sJYLUGPtMchkh
2ktQOsZ8CqnBFOUFjInerUCTGJ/S0rip+/4BdT9SqaV0qEgAd2m5aXiOYgdbDAUNufhBwnfXPhVb
gVemk7nLqzgR8mN6ATkUDoa4aPQHwConrG7IXTZ0WXsq39jPk6s9YHZLCgGwTXXcsq3/DQExYU9S
3tCTqeSA1XSaqgW7AzKqumaTo4yryPOK6QNURHaA5baBwdfmjtOkYeTvUlELzCBDyRqX5Tg46O+j
5nRPk6LY+g8xXK8O/OyGQW/SajPIKjDnUWrXUvHW68eKCcirrU967dgl65mbJfFbIAGlzplWqiPA
ETwMVN0FSZYstq/FqwA2L+ILLLMPiw6WPQRUPuG1BjDajujN+V3PwXJ3ys208H0Jys7cdeFtsBzx
X9JmMLKrfFWxBXJwhnA804+YqO1Cx0f1G94C9fZyaRAXhh6KpMeyhlhzkgdrr3HqU72uX/Gxkb67
HiU/IS6OeI63Q4oiErJr0oOo/7FcIulnYcBSuiKwKWj1mlVzIN2yY2fPtfMfEEGIl/lHR1wce9bp
mOMC5K+B9RQYYWG690qpLAm+KgYWPU+wy+BTviqJGWSiuYUEkpH30QoFkE665SYr9OunhXfWatmH
j+/L2jOX09YPThtGaM2Zaz5QUqwneXcYLp7q3Q96usZ6PdEQXiY6RqeJR/sHtGrWOTMIILXDD37Z
s1QtUOY3KnOpq4ZH0iy7W6scLth7hZcyMgqhwkmHQQmgukwdyYvF/6Y7FAGcX4BEa/gNbSpDOQGQ
W3E9BoevHloUzwHadyUww0LfH2UVJzHVxdW24AwSFFnogFKrq7TI8z7kolsGw4N3/3DLemuahfaQ
tpaxp8Bxgk/mUw4RXE8mtnwwLuIrLpbMJY9eDl1aXc6c8jtSLmcad6mrj2jQMu3Kh3BBaHy6E+1X
GT9DRY5w5922lLLG0mmh1GDMz17WjJQC8V/3iwW16wfnxwnAotMHPpmf9yjmxvTeC6cyEFRHpAra
tYFQ1lhHJbLwPAEfllHVVyeDr7Ns2T9+MZ2H6fYUpWR7X3vtqjVrl/9uARjJEvyR4B9mGxDDcZhB
uqg3uu8U6JYBjuOCIVhl595hp7tyZI2Oyaz+RVm8RPrOkbNHuilQtEIDkeMlhg+tjEn1yJu18RCT
rE2LYzw20tJnB6nWrZDo83h1PpMBCs4AL2HSjbak1yGsZ1ujO7hwxaR6i7veqYyv9w9UNUjnVqRT
uuBCklobKvk4d/AsjxaohibXcUur9CsX87M3O49lbwzuuJVIZyetT/UxBQJOOHHCuhOlS4hM5Udr
IsEC5Nns3gs39Ra+C0ngX8xH8lTkASY7UWTO8KX2Y0wGZnEP3uWbVcg+o1bgv29gylnz1vjW2leX
1KuGq6aBisZMkkFAS9r0iA00/vC3MmdjVk6n1cD98uo40RRMJl9F3xdy4uItcOYE//gHBsffsAMh
FHhSNZ7ZFjCtpWJPVwljQuwtu6+CFDlFZiTNLIyb3c4HJimmpbz06IeA33l/qfUzibkSMZ7FqPnN
2qpXKwPYSVTQN1WF/YPR6tahy0B2d1S0V8clytbzdVPmQFlD/5Pg61apoQ5JaLlgduWslSXNI70w
kbihGCUc33R8ouat1ISo7jpIty9meTSKyBUQJI+Qdmod1GqLGZhsHQCyYL0U0i/pKq3//YVj6nrk
tLhxWd9+b1dkkg7BzL/mfwTpBh0kOw/vCmGNZ0yCkQ184w3pJ/hBJmiKsEYZOY1xB14HWJchfz+c
cJNSBtzuLCA+2F4RkuhvQs0kHWC/O54coFjbfN4YaK9kC6baxOU5a9F0jBqWqRy2vx5qQxPa8FZ0
oFNpZULUyFV5+7aPpxz5o3FCSTrSpug3EvA3zWxzaKDvOcxqUxSdSDd+Q67ytsoYTPiPlNpBaSrV
NKpzb0Yl8hkzp/bMiOBDBaKr2XgjcIOf1RUye1ZAvjrP9TQr9lxYrwDTobSH6GJS4pjMNlZGbnHy
XVupScI/kauQ/glpIL2GXFa4RyY5PSL5rfvqMW4AdejRahGFRWbQQQRiwDn31FGi11tF+bxNetUq
Dm9SucfxWIsB+2Rx0QF9XklY281L2TQIytIkt25qeuAeVb9oEN3XjamBoTDppSRL082yphYQAyOf
MhZJ4Go+fHvSqT6DddBEd8vzNTOJxHh+CbEXEWR/ya1x0d6WbV72Fh65tTWoH7PmY7fBSu7jQYzY
G2hJwcsDVPBxs3qtO/oLS7otFvLaI9Y8mjnalkdWzlYvO1bd9a+ErjbUoXMqAQlEqcArPlCZGAyM
CnO2og18SPPvz4E8MTVxBPKxKEvI4MHI8kChJ6tdMRxc3xXh0Iy0ZtQQ2R4cHT0RiQiVv7gwKM8x
+aBQjFMWfdMq5bGDoIyt618FA/0QG2ScudKwtMNezCajMjAD1VqozRZpPQ/iagIBOGkSGE+L9qk9
a69wKVHZq7GwrLfcRqA1riOWVCLXZTIfPptHbv304ZmSXzjIiYf6WLMRPT4mK2es28FJNcfu0zpI
rq/XHE95l2C+F6BqQFv41V6n7BE1k4VHyDAU+nPiGC+zPXOEyWLO/H8avmPfmFeOTBc16txz5Ppm
YtfiLvbx0zT81X8Vg33fcoAEaU57YQecivYXaYRyfI6sRdEyG+c6QC0QkYVJEN3uCMYTRlsPx4Y2
EUt6W3WGW+SXDzQO/HDVytcASCFnWd13k9zNhSVyRRrxZhAymbrLemj4dE7ahrDuJBuC9hrxOTZn
4t966/I0ulm0QzEJly7KXs46N8jHhrCuS3s0ba9CgG1l3cuxTLiVlf9RPDnPIptnGLvqzI+pmYpx
NWVTANr384EsVccvj2nQ5X+EFKsJ2k0GNbOCQJ786kU7T8GE03aw59b18uiXwk+7nlfbEMZBMejc
0s2FTTjJP5SgtERuO8UblPkQT2KYOheUt6GbgidpPrCx9tZi5G+TzAza1gQBXe5yCgeTUH5Cx9v6
4Pz9HesyCyIBnDunQ/AVwQgKyFKKjI0O5Q4gPIxVh2fgtfqsR3gi/JNAch0R1WO3RNNAmufjkQfh
sCgijxHCS4CR7UyA3ZttrRrAO99seS2zTJ19CVWz3+aL15vF8BPCNBqALM7cVdoMir/lNTVYMLht
32BpXsXxTKqGvd3xZNsoNFTD9+rowQJuaHhpyvVAbxnif7oA4Kt83J1BjMUGSj89cCnf7W2wn/xj
1haUfoOYiz1kmlSmYbCPVM39XMPwy3nfyQZJ9CCEjMY3Sit2egI1nhOzCOuAE+ImdERgt5AFjny5
/XSZPmsyHaxvKUCUlrI6vVcair2X7QZel5vcwXF3DDSFFzWG7nXQV5S3HMM7OfBQToHlmzfa2Zu3
m3u1bmH6BSWPs/QsTZZJuRlgucaKlBLZFzpQrrFcv2+aRog3nFVYGVFqtuTSI7aNuDRGVa7255qt
P+DRLOcOcH8dQ/qK8V0uC2UZeXVImAULazpscJUvvnYqXuOre4llq1hgpgvbppf7ynEPCJKMk+wk
c8dL5tEDCVoDmxOOewemWEg6vmkElZHrK//nfrllFt9FibSBTni7wIMDrBPU3l3ZKYXC0daNm2RM
4Y+cmrOs8JqZuSDwPjDGPmByIFiFEHBJ3JFEwz8UC7Jwyv8sE09bABbi0XrZvdSlU1GvwznwN14A
gCKfSzIwuj4yZ30fYfTJWauwKhmetz4yqXUoogQ7aH6dAg9XqYWbV1OM/WBkmIilmP5dLkfwc1m8
Ia9n3XnN/MAySVvOqfUb5GJyTgnSlgVctr4dBrxs6l2ltb09pftIdFWP0m8DGjq4d3OPhgngdENf
ZoQgI3+KA3oSi4iZtPBPQDDqYu9lgmidPL/WEHx+M3dwwxJlgzMqhbTS4VPqxzF7FeKPqBnZ16OW
CFua+0zXf6m+YxbUBuAqORKqA0JduCloPOuRD/w10S4bVbCYAwXUjqjiJl2OsHaZm42u+cODR47l
rInb4nftdsYqp0a2o2rPrpEX+urY1SANRT9FBJzpUGNiuGmLpiT7KHleGzPO78BI1bPlk8xfZ2Ui
oQU3SRYfss0k+8IxYdHWn1CeJVbOXkx4m/LZ7quRdVHcOnqJwXV8GVuIS/I/s0NItha1Ll7x9Iyq
REvrfMj1N47TBU7GUUVUA1yksnFms+b3xx2rxmz0lszv4oP0uhiSgS0PIJmVmb1YbVvTfKhaCbkQ
HVeLi5QiGQtrpzJ2/jVDvsG5d1EU9FYQUJjfLcJsJI0cVEej5zn5vEjEmprA1EQw7CiZ3ukvVrZH
PVS2rbfj13tBEokrgHO+IrvIJnrVqETKDUmRD7myeorm/z79/+hGGX6+9Wp8e4V3F22KFhIfRCo5
5iXaXG6MbXpMUMOigTpnUkVw9RLho9TNncLPantZGpSMLaXTnFqI/quYzz5Y7FgiqvP9So1/cbzT
jrIWSCCH1ub8dXhtTiSEoMnUPKNVlksnnSPSbHFziTaSkFVbXqS/UhmmQg4w886JHUNGF8H3lv7p
5cDwpdn/subwmuXMtY6lkPYmb18LuAm6vPxj0j4Tg6KlkiuQPq89CRrXp8YgweIitcyrbEpnwl7/
obtwHstmi8erOo7JE+JTan6L79w9xaJeKurS9BE7ykg07kF9Evz4uG9tHmmfdZoGjTU5SnIKZNBC
yTdxcZr5OEDxOvi8kdIV3Cs5st/Umq/KqsJ64orSX8JETiLxNGP8qYTKnKB0T+L5GgPJJfP7IZFf
684Q3khQH+D5+DchjlLgNefrKvgSvXK5vmmWZoKZ1E7dtG3h17VPvOVb1ENpo83qKPCDBLg2X1F3
FfOVHviMCjZaUwaGY4xUcxC1dj3Axu9JdD9JG/e5Z62tiY/CcUi9oRQe692nzp0GGKjwOFd9AVUw
ZUQC14LddHYSjrFsq7HfJVpBItsF5NUtyBH7yhjhghMGUnp3/SGKQuTWu3CTSTaDFXYuMC7F483X
Uk25qgML2M/VDomHrjM72wLcsd10H47lf1VLtKVd9WCWOXGuheejsuJmKkBL8WcyKj/tdaBTLwYr
YwZagd27maGu0bvGAto93GvXxOg4d39+W3dmJNrrNN4MNe0ImzbZOLRNEmQoOq5LH0hE1YXFRM6b
cfHGlV2wiH1W5VbR17xltPQae4XhEAC9SFivvasuc8eVJZ6OINxzm2ciGER60o9JZ+n1ej9XQdUS
/uXoPUFLrEgBF/DPoFY4XQP4rX2jjOlgF62yohFOna5ABhjZwcBv2XTxSmOwnKDVQmA9T7S+Gpwm
mnUUCYebCEL1p56pC1b3vX2Ao5zgXp3G/JC9yeUsEb5a43K6XMH91A5fD8eqBdtvWFxAk8bhuCYm
RGqfGHNEZUAp+JNNWNvYTiY1gsb+zhFrgZrDbjtbuvCciNaPutu24NXAo0uP+dvFj6n79HaTlvlN
5Ok8z3iCT/nA+IJt5OI1obkqqsAvXabYb9yZRO+xI3+42IRcEnFpdjMDwRLVcVWQWLQ31LAp/Eqf
9y0ck84gdYtpFf+2UZLRattMX+eAkL9sVwk6g8wWhZudYoBY/nPtyh0w8fdo9T8Isf0QZc5hGcZH
z+jbxnqqx1KIq8DKc0rz7tpJnWkwwLHIW0lWj/jvp1KIgAkGh/iRoJ68gEnjMpygxY38KR13qM5N
Zcw++8j7Fju0X1C3ZR28QpAuJirNtX5E0sHMJ7uEbI9PtMqGHpXILYOarnT0RWHw1qcfv/HU4Yct
+XQ0NRtQOF+2YVUZBcKY+EOSgrP/gs/f+UcALqJf/Hgw7NSFWIuwS21wcLdizhuSH/iR9kOx77/9
NBq/KnOlyMkJBuVDoPX6hHrcf60gJln15ZrznOIVkOMI9OsaSmdx3uXp0zU3fkSxHku9wwnofxh/
/lTaofbCSWT1AQOwkGyQdkRl4NvQuTGvuzjEkNMOmlJS9L7hCw7e8BJQ2+Msi/Uso4DtvuHhxMyf
IWjJKwkZVoGCkgDD9ZbKmhDSDPhp+RifyY/I4A0Tsc9TmtYppdBDS5Yo4YLmu79ri8iYX6mbzrNY
/fu8UjlUixiGlkOm6IMCaoPeN6GjgvxJE67u5AALsbd5xj/Q8YWpJ/IdpaBLWez1+n2s6EzdTMy7
UQwP0v8U4fhtMP+mlm2CcdojokwPIjkJBkKl/ezYHaayCMuxPrMSe6Eac9ADjOaWUZuNXFWY8ixn
BucQNFoBosyeN4DXYxRIIPXcMphFww7GO1lplj2xmCBkbT5H1LqkGpmJIai0AiXZmIE0neSf9t9N
zqtuhGAvoyGXSaETrCn70/k8dMrd5cS8f4IL6l6xXzSiu2aWJl5LUBHWrVy3g1Gnr6AazoOHF6LT
ZjX2jDX4QzqSSzXqGUobur4cYIm2V6gw20No4Hvob4HIUIrarIc7OC9B9rBQJotSyiIy0Srx8weM
YXWoHPwNbG0uCeMJhlBOQKANVMnFKfy5G87ZdT0Oiu7Q78Z8XuCnjLwr53cLBj+DuuGWgQon5FBF
gM64m1SOIHu+6aLDcgCcFUQj0j6daU+23A/UkupI0uruR0krzfwNQIX7Gm7mDLP06mxNvbDbms/0
5h1diAZsAqII86GSCcWuPdV7uSHrWEZwK82aiM/P/h6jvHibBCY+nF+5Dw7n5MZN8f3pvoTvZGcl
Iq0uXHXKFaJapHrCldGVAzDg4CcQ8NyV4CcDTOyoNj6FX1qmKO8vbzQWcoHo6cPDOD1Zj6x6NB7P
Nx+L+hmGQKlu5nnSHfwU1bzVIp/n8ql9Y8/HRmPh0WDybGp3fU9h+eMIKW4oniuEWMxgyqAjKSxb
eYi0+2a4AM8YyArkWdEAApWfuXGS+YZJ+6mwJNGksSvnA2FjBKVarB2Z5BYGsaj58sjlsGpUYII8
OMD8zDULLeSU5bgIQPso4XLSaU9qulI/ak9A4b8DPdYxOFSB1vc3raCD6zw62JsIYYp2xJFEvdaR
sfMd2t3zjW7KLZinEndsFFTL6633/haiasARhPEZppjIbBK8i691UxS+41o0Iv0up2Y/qfiKUMJa
OWQEsSPmLnXyh9E8zaYtZr6NK2WBne/yWpzcgj1ZGWywMbVYxoI86RTfYXdUkbIk38kGhfMV3urO
SF3petqlbDiLIyj4ZOgqsFOLwymmWm/CUQllYdvpp40sTHTPHM6BBpfHTK23i101iBVjE+urxGm4
0636GQSZIT/ocdVThrpizrj10//QZyRzMAtkr4DEsVTLW3fYCTY+0nIiTARqvHJcWq9mHHO9tA9J
vmx+s3ts6UfhzJipMK3FqHiquQtjYzTj8/RVB6e4Uz4NFNUSTmBOCHj5TuBbFaQN7PAcVuaBqYKj
YBGQcmJAJDHZOIJCb1BwImfqIDJoVmw2RCaBg3pARPf5dXcgeYfrcuHyAqaGE89w4wocL5gCnvTt
uRrHIZZI4i+RUsoANvyiWiWc0i224c7h85Pay5Wq/MmVuP1OYWnnoYx+XVm8GgXirac+PzIBGS8y
xCdiYKHYIKF2+pWFmxx0VHwL941iU8QLjjPl4UN6pwUxq2ie8wiCDvEqCX9LkByM5onIaYCT+iZZ
j/4RF416P+fyB/9UEuw0JRQlNoxLpKyidOe8ymsxOM+GIN/bDuZSW742yO5ppoWkWqIVz5UGTlW1
LveWats707NT/x1/rW5SpS/IA/F5klw61wM6kDmHIutFGW8VgcPD2A0XVoGDlAVdTZUlR27AfFRT
zd6jzi4sZ6V42s8wVpm/lJ/JahnWTZXVsm9U8yDm/nfow5qD7939ynGawCRpRB1vu7pw7Jt3K2Rh
Hx1x2o1cVZM8sGJdWdclQ9vNRDve+CR3Nyu2fo5BlxsW2P4vvw//jwbSumV9o/gSKVDw4mAG8+Ln
ypt7hRKAc6W0BUK63ro5Ewg7TtzCgY9LLHgCOk/n+DQ3kAXVqbHhJ39mJZ7cmdmoKRoTIGPy/M27
YA/70vJGJk5r0roEnswZjFZXywrI0rBFWn5L0IBsLEhn48aTdlu71FtHla72zwxyKDfJjH698wXR
2eROtXqj7zZlpWlQ8h7bGORnCUm7CdoRIx/Buhj242xO+/O11njRtKCnNbzuJkya+IzaKONhvzVa
k2f5uaul3kjC3Kf/2mOIuvyAyhJwOunaQqwGhR1ItxBIEwPLckLtTyjSJgy/Q4FNKuD8GXD6nnbp
l91MVXdO7SsmNzZ54/GnkR3mJhGjL0Gf+8bNqcC8yttYyOIoYWR3N3oV5ZQitePuCBwsInDGNdOP
4Oh4KBK5+fU1I5WQesDkpXzbEqngQF1VnCYELRg/XCeM5zgPzVfc1esddKxHNRCSmlckyUD7ypCo
mSbCDSYwej4QtNqTYcvMIaMtq+jrglWi2/OsEn3O75bvYh/nR+oymhhnKtDspxg5CX3i0ht5dkl7
p1Vz32gMBDaN0gkLWUDGYR5wUtxcrrvTBQ0lBUPLueSDtcymBoy5AaNh3dGa3HqWRIRJJdn3DxXM
MACdlBXyzv7dCYMAQetrhLzCiLeD2MW7eU6gqCtVEKe0SwSSbb6ngIoGjmkA3VDs26dAjVYxC2G2
xVDtQgRpPOy/W+61S9okAJL/5XtHYYsjXDIkKDOPeasS6yaogvfaj7aAmNwSNycsez818VZGna3+
wr3BF23nbMlJu+SmvwMtl6UIPQamzL5oss63SEi163seSnd7L0Vkc5sI+h/tjvr/7fQVrbfkLNQT
76qJStMZ7NJ2bUx/bjwsS34SN12leLXFVppDSCcClmtqWgr+fMe8x/uF3O1e9Xp449WU1TfvCHbN
poH8xHEShLAtwri1rtndkdl00C1oO5hpY2lrg8YqUT0Orvve7NTEfv17HeMTLNgRoqEz5E8KrEbE
VYXhY6xbv8H6qLhr1DIO/GsC7zIwCfm4Iw7uPMrpTwLlLX8kAuWe/aRf2EZEFHCqW1Y+SBuQqJnx
EuH/kLQ8jDhR+TJPuHCJdx5c7owzpRTajrmGqq2kHsFphWKCWQ/GaAajiJiIfHPwNdZjAgbrF44f
2JQ3nYaZtTlPO/orQ9oNxUq9M+lSpVqHc8CVv/MrY8anPVxKahCj1/TCOVul8Qt8Mufr2dxyOppZ
aCum6k1GD84PVaEiZmLFuu2SqgH/0aJseMrFWHXMZAHZL9QAJi7YzDwI2Mkt+sPtPh60OJJAmUUH
zwDh8xgmDfOvhevqfq5HhiqVJXTnl97kkMrZwL81V2HcOcWpO5AMEI0ZEhNnF3q2bE9TQ+1iHIlP
iw51LekfSrXnlt9wJuEGyRRIwaD6sMT/JBKwew5vgT7bMasZI3tVH4XAAScKava9V8AIi3s4ip1l
aOWhZgpb0gwKzFOn9zDXivRnDTjBXnzWtaBalcDbI2AyTjMWHbutFHIfeHKrRmSHJ+kUJRcDmHgh
V48gNNvTkGjrc/nTE30akPvCWUZWaASTxvDy0XGOznMDM0l/JLkk9ROhSh71h6fISxDkQzXlW7zl
BLBoRx1FGL8E1LAKRwWnLAzFLj5gJ8r7n5IZl6yn/5vjWqmILwQdm39jXlG91CqhaYHfBWaA0KzD
D4QUXFdbYkpzO8C7A719s4UkGl4dYgHPXSjHpTOojO08k93Xun1kQToB61toT3pCCDl9jSC2J4hM
uU3JdG0DN0vbsZuE4G/3QyT9l16ENhUv+wZXp8Qr9r4i8sQ4dCrPouHjNbHtVXtttT2vMdpqhQhY
pg27ZoaPeT7Xqad+QZkvvKV00eBG0K6LUgAHWX6TQCyHCCViZuxNR2b2VPVXFCNViwrHDVA73U/L
J5OX/uri+2tqAwviw294zIrL18xjTOZ90k4TmrYE3amy9t02n1tZUcSJlSCzYj1KDVXRJfTrVDAj
QjJ6E3DNy3r2GGbwHUhi6ijjfuGt55KA7IeNYadnx0HJW1JrmrKGXBBiPUndE0xSwe3Y25PobQuZ
LT6g1NGNgYuXiksgLfJbNU6qgEe7xuSk2RHYY4DYfphsbjw22eK2lYGBBoFLOxGjgSFR6/jBayKc
/auk+TzQVlupAJ5HbjTaqx7wLgfntVBfzyLek3Qw2Pv9rG9f/aA6kNEVA0uKqrwkc4dPiMhD7PHr
wONWQB+bSmwUJF1zqZJ99GeOyFEsdhs5Uwm7p1rFZarwUkyd4+5yufFlekXSxPROEzEGEGTxweAP
hJProQUHa1nBA85phMuTwuVmE0KBiAsZD/MjUgQVDuZzHHdky78+PkR7lH24og0ipYoMhAGn+TCX
NqbEZYxcscIdlEjZfMv4QI7/5vPXlKFnmyVK5pkBIztg1ewcCNGiLCnXzgovzGWYmLrGRJSi7UYB
Zj/WZCwoC2iwJTfy0QBAkPP1X5TFXD0BSU3zUOeGu78/LrHLKt2Q8rLpxePRPi7uDJZwMyxFpid/
l2vcRGjN/sjbkejoI/VCYwQV4QBhcTiPBH1q3jkWNYiPIBVvjPs/00OoAVAcmJ1+MyzXx8Um/dci
9imNhr4f0QvqTOzdiJ0yTnBUgsdsitZLURoYZTEnzPatsGpGx/9Rs0M6mvXSPTl+FGQQ3xsQYG1L
/C+/doozfRSBdzwGJ4DzEuJYZ6RDTdT9INMXPjXyl41HxhP5nRzkp2dEhCvoRgKxW4gv/hhMS2c3
vvLNZLmaJPSZjAZsUkMif5L/UaO5OEgeITEKmRlQMXjxidquBCRcyUnlDxFyle7iVZ21grhDLS7l
63ZJtQgxzy+vsT5kpqtCaanW1TFOKenheROf2aiVpnptDuHCJQHAEPVZFw/5XMDKjPANv9d0u7Xw
Ss3bl86X6ed17xr1dBSmj2kVlgIHArehbkd3BJgvotZ6rv/2nmp95RCKC5o63mnhcRA91udi1lpd
I/VySJdwHSOPm8H9EReXigEukizWocEjIlasEYa0aS9iDWddp2b4pQa3kQEAV4EqmYaiQLUFH/Tb
MBtMLAhdGZgLLX6QNXlQXrgY3OxmswFxLXU0ANGMIz3n2d8VapdLySKX0xOf5ZF1Q0nFr1CmxLU1
RULYlzmzLXnkNvqVBNOZICyocULLqxBT3A8AxfTe3l1+Tw2FivdvCNG73xQNO3n43cKhjgY9Lafu
cSZRjsQLO3JAYUXxGivQ+9PahzdbZHf9teW5u7Lz1FIxJiv3yDisPdExC4XpDXGX7sZhxx28FIGk
KXxhDx0eavvQe2hwRoKU5py3sUHkx3XcomYwZLgu2lW/uhxt5JFO0z8gwGpV6z9NhGylGrr9jzPu
tIqy8hRW8e8Tput8zQS0wUrkK0h1HiKg2BCJyzckCMajjfw4ZYMHRwdydyzWRrX0WIiSlAclEc0J
tcmCuWovF+5FsqkpDyF6KwIUb+kCCztk8dEOTjtRvMCbOBdllImiW7i+OFvsDuHuX0RVlYf7q/86
T9Nvkt4EFlD2KSOCjs5sYPcSL8IggrlisKKtWqLCPxO5pInMM8T0KnyXvaBIQqTc1WeZ4m8ngEXU
AKwEpa1NnlF/tzW4Ynt3/2PK8c2o00g9tAMEddHV7IUekPwPnR/z+JDW22BBMZ53xg+qplzRaQIh
+K5+cXFj2gcC3Shs1TZ/1xaN8P7qmSDoL7rfY4kcyPibsW+MsuRsEbiA+8kecuiqRNhPjm9MaYNP
djziCgxW/NB2LphcKEcqgj79xSoGTstdn498/wPWrq3xxZ5YqZwQn4xdluLEnluOh4+6YoYQO+Wl
RAG/taXPd/CveCq1aeeo0ESCkgwKLZXxz8GHeK11AyV8RbJnEKVQxyfl7WpxYDcSF20E5KycRvgZ
GUzRG9MU3NjjgmqDvlkg7noe2OlBDkhd07JxsQHW6FTwRqOrjQ2Pf/2QyoYVVMF/SlzDYZDRQZJe
s8xQXpY4jXfZbY+s4GfubFpVeaDsBh4d+qLIE/LCBr6Vp2DRAgcLfyu+ip6z4gno4r0WNNuw4PQw
oiFk1VMs5RlZ46f2vplJvAcp7chhY4x8GvXxfyh8m/7jcyHbMJ8zgax/DMsDwoIsJaHcba9GAAtp
+yZ1dQu2B/Z4KmfqoO4qYzsFoax1AF4omy3nzsqMuqZ3pC8iA8r+R/X5HLSl7jc5RKZyM2gEN+53
/M9fh5P+i9IHOpqufDDy6K94Du7Qrr5LR0lC3Nh3uTAg2TTKSOJXx3o/GhMBGrXY8ml3GRipb9G9
x4LmKSMlvkX3M4sDMCqX5DUFKLOqB8gsu3LXgLE10MpKnl+2tirDujzqym7BOAxtd+fKH7gvTDP6
KSnK144t4Aunf/LO5eQjnIM6zmOYdTFNt6qT5y0TJ5oLAFtTEeVK5txG/N7kPhFQzpBDOxUBnBUW
l1Ng3BBqqDCAc3+0zg18DkpwgCKrE8uuM/zQO8wTC3SvxrHg+KNw/pVSFDnApEvL3sFUBD0XRyJm
6b0kRDDYoeDLeJ0BrlPvyq2NGrXJGwRUkJRjQxiHwkYMmq4HaYxdWtcHPBYP0PWjTjIfSYtdLa2S
OWWpukP64ZERXSeAvNqqDkyw6rYbYRFEvkcrmCk/Weo7Fs/rJcD2/Q/TajxMOjWA4liQTeZtV41G
/DvXQIkXRC0KSQWmgjSvwTA3538yumMCWPMT7mpSu+T27n5n3Z5kR/8w091s8TubRnXtK1uDrwK3
dog23a9qCc/T8X1tadmTTGGp8ZaWNcgHrWecgUydgcvYbm7NdIfum/fFgpeWkCKIYIxArk6srBnW
dNSprKychWOYgzXLo3qAkVB2cwnOiFeo4KRRjDSFQ68i7xXd4X4eV13MHW9s99PMgfMPLNXa599D
3EfGsKO8dnFz73v7X/FVgL2DmAlXg/FaVFONiOsHn5slVP/vG6gYLJb4ni4kdFKS3t9sqF5NiuVE
8t2KBTgm1X/1Ucqjm1UXAcF5ke51PzCQE0LsPRw3kKI6aaxkmmsd9t7YLureybNqYn7deZn5lZxk
TEwoIz8ZK2a9bKZoZYqX+8fKDzAF8I56lxvOicfRbdyiNEAG1FG1tvo64kDTG92xI44vmJKZeUFP
O16DoZ8OFMv6bnbo/aRQNSXcsmAnfrn8ckVC0pJ0eeYWihudg7u07wDtlTi+YyVUvccnoezblEV9
qt9F49zhhJ2v1QQAiFb2kZ27eJ9jxmgEP+ZZCZxPwazpekP86eVYx2ARQo8QPXcsJOwPRZySlg1p
tv5ewLfQD3Md2pmZBuG+efEuBXk1geCKt0j0zQxQyiHYXPCK6kZUwM4EdUeWNiOytG0FEKy2ARNR
NjNzJ8Ce44z5unQ73vm2nBiwS+6YyhDkS58ZVerWyTvTnosEz/rZespqf+Iu3QAx8Jq5wtmZesf1
574zTMp9HL8ko++I0+7BP9Ll4ORn+V9dzjec7wT+H+qedXVd596mcROPCs7wJNOtb6wn/yGqXsFc
o0dDJ9A73YE//v3eyRvp3yWJg4FiML0JycLxWPw2FYBIrkPzMgQc7iGcpyhud7aTPY08KMgchU7n
2hr0jatnih7w+JfuN24HtX4TsV4fxQLxH5Vzjig/dD4eTd+/1IVPBzrwPrbPSvDeBGDwaFIrXDd8
JtORW2PnbWgUZvqxcI+AH4jY4pXcKpUkKZ6VpQK7rA/V/bAlkk/NdOPnazox8q8qV9eZC9AHIbnx
zfxAsHJunLlLTyOnCjPjr1KN3DDKir4Po+WiaBIh3V1+d4741RCX8MLPBzES02qbCEfsSU+P4m67
y+d3D/7vEw9/1iisFf6Bf5cHou+7VbXziCNIePD10/GUCCtFvD4H5cVTuv2uXpcwLU+3SFuP9EU+
U9OlabHYjE4eJ0yhma89r7EPZgnKdNHHjGtWUPc4eY8yyg8mFoRb8yo40mqcApkNbYQo919MqMnD
X7dtyLwG7CLJKj5TMy0QLTZc0dFd46Yr4CRjdmjAjBcKx/zX5UnSOJ/q/Ts1Vr95dQr9y+PUdoaz
lZJu0KuZHRNw/yY8O9+/HfsHzEWg056YLtq5FKHhH6E3KEYWxCTQIDdZLY+eEdrenEWZKDdwGRmD
UCIyvbcr6pO4zj04/aS7qoEga4kdGDjfI+2XIqrG8IbA8wHVOtaCIgBQHh7UqR4wxchmh3Qz7VG1
+FELouy8Z006d/HjAYDVgc93LzvBCvY/TLCuC8hjnIqfYDRHkW92AXPsrBGpwwLE0FL2u2yKgm3K
ttX7WNTKWTe+pY9hFaCZHk4d+s5ZsA/0nVDRu3RyvrTaokgBw6q5OYGN6cwBK5WJ/RkzC/dXdSxC
PyxeN+0dXreASkyUvtPufdwV86vHLAE0G1OM4OEeXp+1vHiQ8uXrgsNowTJLoAES+TA3eZs+7Srk
cId4x2e6sKDyHuWH/TVddKMCDO55fsypxnGGcbE4KE8JnvwFGEFPxc1ZoFc8JCap6NXyIRouA475
Tw47kBviwUYELUopbth0mRwQ2UvZBOVaOqDKTFkpepcIpggVqSuU7eWU32GwdnojoEKjyHfb7N7L
0R4LrsjLc1gRBIcoNle3Q4SwVxc1lAeDZAm9YPK72TUn6MLpU3jwW/wHgvZ8IpW1yqH93mkRbYMp
uP7ltIZVatdj5+C60W62hBLMmMce4hjK9HwSvfGI0DaAjVZBK4YRh04ki+b0CbDb0lQ/nBhb4RGY
rOAILMV3iEDZPgChz4cptEpbtZtbLVK6Vne9nZZxSY+VeN3O+2dNo5lUYCaxrFkTdsh9XuDMbBEe
0DIlDYW4ntXvMT36Wc3UJFaehx+QT4MpOKzBwthtlzW1k7391CbNs3QMQ32iZKMu75+ffA0kdwhJ
LgPL2pprzzctVs/cKnIMxHYQv2DBoaK/p3+bhjGXERjexx9xu3skIPYJ+SlViRDy+K+AYtJYEI2y
SXIQ1orFGkexaMpJhNg3Q0tydsWwLoUGYSCQM+cGwh6aWebW5Fg63TgUULfOrizxa95nKDzpkG61
93HMF/X60zXhKj3oNDo+c4MjlYAWhsEIMeg60ExPWHQH+niJC+VAWSC0yryPsBMjoRlo2HW4mwOX
0kGZTjV5mVL4yYCNHincCUgnLU/8WOjK0sN8730yKOWdOcbTk6UxycBib2aWvrPjiALVVD8LOcJi
vfEi++xJQjNNFLChLkVxyoDmV5Udnx9cpRh0/mHkNO5Aq+w6LbzwVfB8BzChhzXXPnrm3qUzS4jj
JnxHnTzzLOzUdKFyeQjP3WvEox5RUbMODdJiDNdbtUn5vJvmP8/nrbBzJOYpXWK0ydVCnMnWWHdq
MlGpmenu+2H6M+z8fsay7hwEHrsYqEDxt82XZ8cX9w1FiQDrc4wepz/qTckZSFlA0FxeUy1gOWki
6LDV8PCuAzAgb0QirV4P3XXglinPZClqLnzSzg/jKT0kd2upf4kG+8CRROMbFmGrsDEvZHpoZozC
z4yLLel8DbtPwWXIfGHKur6+2saPvomQ7vZ9LkYqT4Ac6coHCtJz1y3y2dfPNlhRZoB02XFFO2Bo
qlrV1Qvr/rJauA/ZdRAbOoaZB3YPHxaCwePuuzVuySns+xPQ9Bey6fovgOjbecUJ21CzI3NR9RXS
aGZKeoPv+k82lezgRkM5NlbT7H4zTT6GocLXS2/VQjcpHQDCiz2ibdJeG/hgONupXmyH0u8lY7UC
bSxTEheRw8wUuJl2I6ut1236jsfLkjcPB7Af9xAbXanSqvYDYkOSGkQtwyMJ5LIHts1+LC/5kFca
LehNKYVPyPNU4ApGw+SeOHoX6wwvyu/WZcUpjphciVOVmgfri62exIZZEDawx3Om9yfo15nuOtMM
EpyXxRU4HibTBnw8AWR7NKInKpKsnjFG1Hhx43qiuhqLIHD3gWWl4SmxIkExdcGNsk5zsmd+F2R0
6hTyeBYobdeUL0UxDVGyscRNyPGMkV7v5VFWyIkA8JIJ5H5x/r6w5BN1/15/cYikb7+MBn9sTkB1
X2lX419njtQAyXMhRnGUUbNkQ2h+bkaQxhnlDqobpoqgOLHFrl4t5TlU7cxd/ojydnUFfvvn5qpS
QsuNVGMyNlNcoY+j7pJNe6dNdVhFVmAFSMAGB8Efywm/r/e3xki4BF8pRkh4arryoawPr1IkgpZI
Jj3SDtdKkMZWyuWPEEjMBc5CrTn8sL0NoiRW/h8AXztvWeajt81ympQFsx3xM1r4fJjB5YIJKCay
1MXj1TmN2mhXtFYUIXpHXgemHdRUHWQcRhHTwV35Oag8yhysec7ORzqnJ2Xwi7nDyKF7mZWthmfM
9e89J85nDCek9Wda1i0mx+YdrmfuLyd1YOkCLshrWx0+bDGt2gNkeAu0dFWEdHIzPZ1qYp/o7myE
iUKl76LGfWPIjsmbmFDtcKzu6DY3mbWC3I+y49jTNlnuWqlsm99FC5pxkI+U38/qvYuYQ4Lt0Y0k
h27h0tA039cH9bOGY7Y+olOg76He2Od1bNZJTkR2SUtmtCu+Ct8Xw7aDKK9HmKm10OGecdYAm6W2
dUrjjzHs/IPPkKdJtVmLt1u1kVzZhllwkb2RVMorJ0LdAG6gKUHnDLo+3gJgiFCwxDUIJ+4U4aMR
lfH6vBiFF69A74PMoQRmnVTpkJNyxNTYZaHd2LZ0cb1WbgEiCIINTrwMwku7IHQ4iSGImBOg3sJq
C+oEw5V+AKz6mYS76hGsVfxZqrqUGUfL/jCld1s6dV2nJbrJix6uhMt6tEDg6cNLAdiNUFZskGm8
7lU6kTKOgXsZOq5rLSU5/hzDS6+K1OiFEqolUu8YguAKnVuxny+WGNy/WoYYrmSpe5GnF0pHpFn4
+R7jlBQupyqKHLzobCQ5sjpuF3X8mC5jBU7lzHFC1LNCKZuTkROcxHQBH6XaJ2qAgp2u37eaPuVz
59MXOTeOS92rVPX61dNXn/JYapqxHr1XtPO+RdTyeHJ42/MgCf8s5JnsV8birWB8NaoZrsrMp4PN
4E+Pl0nMBTnR+ZTXum0yjar3S6SytsaCHzso8rc++wTqUvX63nw2/KC+6PTUSk8aLbKa6xgxm6Rw
F4ik3gkZG7SSYJOxV3qnhrxspIn3gnzkKyEEU6Y4iFPePFoVrbbKn1tRfkQb+Pr0yijfeUM4dAMk
ko5Oy/PvgHMZpePjkvS6UwCWQr9Kh/xZPqkTo/kG7cygtCDKqv9xJyI4o7Dek1lrUKhnMusNrZBu
DFQmQ5lAnGPNjsVuLHahnKnG46XtGizNxNmG7p8h7qyy/uarzkp1CM9768LurmhYMrEn7TVSZL+o
nV8Q9/juPZCjX+Y+0hV4jBPqwAFOfC5/mpJboqJKTjOwweN+mDXIOz29tjHsk8D9UF8/o2zbDhRd
tV/VeKaGYkrkQdpOJzzEJvl37rhhpmuNFpPu2GENapf8mWp80FJsmlBXNwRI0+2I4fBcoFpe+hzT
7He5GSFNn8WSPWdcpDzc+APviMCJJHfbCO4qc8XvIun2+/N8u3Mg89eXNckeIFTM+qpWoLB+MmHN
WZGPMrkiSR40HmxtkHGAc230xIQesyGRJVHqQyy5t7diu9FkKscMr7r924AUT+ktJEuPCbV5CzDE
PYYXV5cu/rTqtBIAwUlEK/zs2dgRG61iiW4glWD9BFl5MtjD+wQ8TfSsNhjMYXAtlSE6yXmWfWpu
Jo2bbJUr7Qb7dN217zxahRBjI0ofwHN+PuSa9PXRfOxpwTx0Kl1j8aD3NSxGXf4I2Or9eRbfcv5W
4QIJQLBZQCm2z8mV3cuPR7olheS6GFzXxKE+eEV2SjavXxT6w82FpjLrvBor4X7lGgUvrQshcdX3
/CYw3OmuqM1OIbiZvv2XsOVbrWsEB0v+z4FcjklNL/3YeTFUR0vIIqhCoa8OsmgLt4oNR+JjIjto
/MBV+u7jb59PrSvxmBmAyt8FU2D6QMgC69wF9+jhdf8Vz2uCJKu/FoLY+zkiVhHIWhGgm8JT+ekc
FNfaWFGfWQgx1vH/2pMlptR8coQ2vYkAC8aAkvrAg9nab98KfV+0oLMsipzbfr3PkpBv3y95vFZm
RpdPeY1jmFFSHIz1Wy0g/zR4BxTx0I6yHHQh3uy0NdoaIB4F8SGVowzTjqVmOF+QUMHT45ajLk8F
eeimvqWztNOMh1Wsq51TLMyH98PKJtGeIqCsS6NTQhEQkJKRPnVMiPYBlYxQsWMN0VsgEhHEtUTR
akUltSAPNRI0w6SR/q9rACGbQ1JZWznAJ4si6kA/H+Pe8ezATHI6uxI4qVSnUhiS32sC6WiVWL39
mlDUNsDiFX4GGk8zzn74AMyKCxueA8lzcOvcgqxmmGgEM4jH20A0h3mYk3vf1qKK6Hj3XdzGJJ5v
avlh6x1eOgOLffhd/qcFBmIL0qfyFWWXmAlsz+Z6oZ/0OAPfo8SA7eDFB0Ax8EOilIlotYChh0St
xXSttgq7YlP5apXg4gcpy9Lp2B5A6JlVpiAJdjit5EECqsCSlDBoIZXE2anHrDYQJiaYctX3ekzz
NRdL2J0ziFMqePR47/WQbLZA0s+L6tuzMZd9o0pEsJbkPLXiTI6PU96eqjGOH8VC86XlDt8aZN3m
tA71tRKQyFLazjofyM4vB2HWacT/5zfzgxPAEL7MYFCyfATJdW5sX+OdCuxm+OTdN4J07Dbq40TR
r8yUMrPnCfGMylu686DdAhfFevcHyiN3zZ3wa3cemj+6B02LKEI9euf/L27Q/3DRFTKn3h6Nk0la
MIwTS4auIx5JeaWyGbt4+rEatdV9yuHB51ZgsvnDESbD09HZMCZ2rq/EsZn5fcf7K7sYsudlgY/w
geCuuXo5gmpvaJwV/lQRoSKMin7r2ymZr7qF7wKSDe8CCPCq0qzkaJDuI7hs/WC2pI+C2Do03vDn
ls8dgqJSbFPxv9FOba0DbI91YJ4+lQ3wNqDhCxkbpZI4/FvZN4K592flVdAa1BWVtGImxz1doTPW
FzioS+ebak6GeQ8/O9/nnhC8B4QkPPErczyQkbSAAOsdiQxutreDepXDtB5IjkfCqw26KJtU72su
UXbA6kosrttQKD6zaJMZEiRxqrFbHYMKssUnMnj4UUy3MRF4wXgBaNnQ75VmEg0jtIKbZnczNlK5
0Rs2nw2VL4kOPUrVV9gosMG+WlQzNcZS+U524Ypv6DMedHRzXvyn7a32TKjtxDGKho38xbkQQytP
CRh2fHWMMGDDtW8yPQMyTD9LrkuBfirFkJ6sQnKiIiBgi0MK7aEc6gJtapJxLzihhxFlfDDZrAVp
g1nkoWuE8k2bvQtue6fO1M7AKZF9Bw8nzh1VLRpBlhtlAjtkS7R5nYPwscTBehcGeS3u5iRuY+am
TogMrK4iw0qD5ArmrOkmzxqCd3PnN5TprlxRmP6ugIq5QUOuxUNpchcEuqXMEB15gYMxuIHCU2RC
gUGuka/VEgMLPRhGYlT2ZBxMUwKKlbmoBNb7ALU4CLAttos+BUKn1/9VuuKypIrJLuddCoAE6t0S
NHGS+uXfsRGdoaThpUNOjLqf2UOaFiuNHLzJTLT5OTYBhLw2/6z7WW2e1IejkvexW5KhigWBDpH6
/6SXkWLLZ+TlOtxswWpM6CVH1JSZVIu51RAyD1i66hBrzUjFMtO3+Vkt0H9XWCyR+cqp+glPeuE/
o1c+YBWYTMxrLq5FfAyiuQGWTV4ayqR8VEnght6O0BnQR3M8+2VfRDTzH6nIsSPi0/l5baXO7O3O
JskVpf0h6BuCCwePLgibSy6nCSgrvvEHEBYKZ/nE+2WfhyYG8f+2M8Ja8pDMy2z9eiK6mNYd7ltf
OO8kV4chdRQ6dUA92YDNDlm6s3xHCDEc/RvQUfHCNDgPVW+TMcLjp8U7zpUADDEYnXXEx76Y0GPW
ZR5IjR+vwtg0kKKMg2rrk1jTWErbeSoaoOtOEkLOeTUo1f/3xCIeMLCje9VJfQm1AuHiZCPTeIQW
TrH9mREfNlz9lw1iU+FdiAdCFdVtcip9COBZztXsVjam2HONpFO5SRKQQaM9QLT5X7Eo+CiPzrYO
MewoWKS78wiPrJB60GwUgcolcFSjmtBUlKMUJc5A36N+ngeLwDInW+XtufoHdrli5xiMxnyjRor2
pXVf69VzniSr2BKN6yUSki1H9CMEF6dvywlILCUBu2ppNhGO81IfyS9OqAA6cSHHtoIU+LvNvfu3
/Z2Mz6x2FyhoztUX0kfo9wazCHXkC/RIim4WtQGavEbqONSdai+4L9RTCn1SR1MnUHS1kgaAtrYF
NUERw9dMrwadqmM/tJInB20cZZ8WAtoHELObOvL/5mXt5lIT/Aii+gN3A2ZxqwB1GZR3WJLABzMF
B5X9TPxDP2h850Kzc02fLW0E1osbuDF8JpU1M+LXO2HsONHLKFFm2yfpY7tLNNRiCxDOMPaeKY3S
W5TQG6mGtkHfVKHCKzUtaY7uX1gtBFY4EiBiZXHIRgKU2Wh8b/T5wPrOLZdKMGMmpJaxr1suuD04
4QDYO0j4+UFRnVVQdwbUOmxj9USlsgqMKmG+CvzGD+kO6SDQup5yX1NvUwFo6m/z0/XOu2zk2Btm
ndCoMGl2i7biBkB+Mry3Q4RriK0RGViIDEUhh9VPMXSFXoX1ddSvSABtcoZeN7+6QTynhaxPXzXl
wcLBB2+Efwh7/fLbOo7HmVQntiBAwQivVUC9ulU32EKg6vsOxcLJxRQi3+ybc6V43gnDgtPcxShc
BYUJZ0lE+SoDDAsXcMSXDMgX+Ox3XSPIbKy9RzllYNFO9wmSWutms8usOf1sitg+vINDZH0UOAmp
CEda264SCm+8ZroPFbLBv/XE+AimvagQPmp0kKIjNEIudP7ttVmlBgqhY9NNGbAdOOaIm5kBha41
DT4002VvfFt+52S2yO0KDcwBeTdm6CQQH03Z6f6IFgrnzfRzTTSVYxC9DU/dWVtvWiBw0JHVLq1G
H/Ie8gYTDZ0GuDLa78bYGbDliDJyJyLWaxSjG2bH8WOYG3AtQgSo0U18BTfHyY+/7gIC4cJdvx9Y
xTQOpe2TdjUX23ktweYbt3rj5/QC76s1rNpvF0l+UCATBBELqZVGKLDRr5jAVbonw051dm4+rOq3
+Yi8xKzf+/BrpfskiZXV4/I76Zjlhxuvfihie50SAK8MHux5x0YYq/Cdfc00CeGrw0GUqbQnMjql
I+4HPpiAyMITm6FHrNqJvot+gq+Sg7zEjzP3H+1GH7I2gmH+992K7yLEnXwnEnhIDIQCE0h98/rO
ITp42CpSydEp5MpKx+pNj1BlDHSvncCtl+wm+bo3JqpISOWwLdk+Pzwr9+QeQ2fZvlroSPo+Xkbf
0ABBmlzy3SvcswcPwQ/qBGT33C6g2DlNPNNTBjHEJUUBQWpL+Cu5SpRWr3eTxjBsXuIYR+WWCvY9
oS/WTDvRQRvaq7p5vabmssJB2GhcD3hS5qGSg0M+Gj9ZmodbtTrk/kAvgD7X5SL2PKaMXKhVI3Ww
dSSETP3qWbPljYo44MeaVyBqz6PIv+zrBitWZTHE7kS3mGuNsjos8dDw5S0czcV3lgmOfiszINGG
/iP3v1WZTNF+FPisPVw11ipB/xf0YdCEA698ETKxonPEIBPZ473n2KdeK9IDjwHDUPKwDykfkf5v
jktiVNyc3pCBsLLrx9dzFLwIBo999A3hyRhIJPsPzMB13jw+vPesePPlzpNcGG5qfdA2H38ECT12
OSHtiGTT8evA1IO6S3pKTid4SfBmaXDbPjvrKkQpRn9u2XpRxlckFGc8Ct+BPudvei2I0nmxsLiF
PSink9+KZ5tUBmB7CPG5YFVHiRdzmyndLDYk9+ISa6z89aDqMkcOLMRyQymgipT4V7Ei+J16jaGS
zw+hQygi2OhOvUFE+TjyLEZPxYJtHQfBg+OZHtVnnSDrDwNs5+4U9OtyAMVrfRPu4lDUYWSO46gO
HPzI8To0ZcieqUlbaw0tUZYaRh+z3Yc4Ep/+ISQbsRaeYPdmfQrs281nUjPIe4rtwzokJvwgkp0N
xO5HJZdQSqzGk/+xRIooTmg1qZHCh/ZLbRCuQsJtR8pR9U/oXGS7i3/bO6K6fbPu8ITUys2GaLZs
hlKvoCOXHuqjTeRwG4xk1Tt9QKZ4GJO7e6KVSK4ZWMb1EUwLVhGYB7PQlhbfg5yU2OKz2ah6GxMg
MhiGB9lEVMyzdJCfh9SnCkJoATa7n2NizapuBAUlRaFeWw1y8t+xQHkGL19+wGGg8if44fsvwcMo
hsJkNLS0MER/Ux6gOzmXTwaaiPr66zYDFfkl2svg7fKdLXRt7VHIJINBEYVGlrxO5w4Klo9H3I97
hf3tsZ9ku70/iYAi6V0HIMuDFyUhDsItfPUYGFek/UXnXgjorATO1NjeCIL1bC/NPQpwwFE/chJM
sQjRa/wwtUcvWNL5PyQ1oTQcEj5ZHBAgKtU5JNRyL3ReSt0azhDQ5BC1WGim+hHBMgP7SbNidjpM
JwjK9C1xO2f3lDP1JKX9IswlUzMExJpe+XC+tjlOuO7QhbUmZdajMAzTw/dOTrJJPoPZsgQiTFWI
EylxMEHTA1zeynlmBBRQacPiwK/5K3bMbe3Ht3fEewRopurCCRECLv5aSGXm26Vk09I3O04hbOrw
NDIFLl3Ni83zG185BdZORLGNW80xeDGiO3SoGWtP4nbI6aG0sAIoJkQrqSTpbA8/82MAWTCEHJ2p
+ckiClQE0/BD/p//7FpiLqFEbgVo/rgykORCnSfDopaBVoaeKQ2V0tRBAtqR7X3squeXbDrMfz5+
Vu1NhspIYYnyN0iG0C+krCiKaFfOK4OJpFVia3pi71V/3AlALP6toyqqrhf2ylY6H0+64ZkIAeQC
06rILLET35Owwsr/b/COH5l4RvhFDk0MXqqMYDhXj+xk99TaW3/OA8q3Pxn0RhqfaC1enJ+cQUqU
mqI68QBNMLcDxx5qmrMnAEmXm6ABN6cE38z+HbTPuZckl7tDvnW/0Slzfq60ojU7XyX0QSCXT4/n
zKUtNoQFE5AIvSfRRsQhJC5RjYcACA55Tkj4xBN9Eq1a0NZTCW/RFK7CuPLnBuScDGdeAPvBTCx2
nLr0kBBYDXICyylCnMVsblli4P1c66CC2h4SdbNCcg03TZi3nHrhfD/rtAxKdUOCx+HNCT6++bFa
vUkU69YKRbVl2LIFFjaePXDs1LKLuvwRqF2wcYuTgns4HlV0kTjbMl/FxOsGZe1B9NbfZzd/ChJR
0SYmw18Qmd601dNFnjja1SvR+2XXNUbI3twCyrz+8GWrCvtp3WB8Mm+uqaj8oAbB1SyeGa9egXdv
S4q2vnKZXWEKHrLjwMb/CabH43/Yf/WcoJLjMIFHcVO/Y8qLX4a8tvXpAmtEpjBfSMRKiirFihS+
24NDlLhnfwYz2rUIwkWcyO8ShMSWFie4kkJXuaj+T1Raj4HOBfbIdf5Qlawrnba+Ea8S8dCNbyZP
Ml/NEKeYtiOjG5sJnEs2cgoz8eDk5snnNRqu/SKNC32k/Xgmeo50rAVZo1T/heAI/aJAXsR2dIg7
bqWPiIQpv7PQhVurj3qwLz4xAE6KrnGfuw7r9xj4uJjnK3B0yamfj6mZNAeUyGWrJ68L5Ksuvy2c
U6C1ZEmaKxdC3pGlnGQMfwXvljdRQdZ9R7uXHgCzSepneBQVQdT7Sp/ZgfG1Pvyyiy/jCxbQu+yc
78TkmSgxFha2VWgw/HMLMKWDv6eMLERSSrKo+mo0FSgZWNfQzC+hO+H/h7nTpS0RZuBTCHSYKptv
RsH0paDrx+h3D9pAzBUjzID3X00DiLCzCeyeUcqU7wmP2rZGcw4vdk/x5K1UNNYbLa8/l2sP114N
mQp2f4JOh61r1Nobse//WQDrdpMf4KD2FUKXbH2aGOl/ae7ACeiz1R0L9izCOwkebuSv+zef3TyN
/QQRVIRlTcRpS5HSqW4kZ7BA2eKzJg+6AbzFSgNQlnO1DXs2UDZ1vujaqWqWm44j2C5w8Q9rcK3A
UCOxMvMyZ8y+d3QuS3LKFa4KsUYA96DEmZ3ztpNgcKGGpakBnW5yGCLwk6a7NI5CKcQl1ZT40PNE
NqMRYQ1HMiCOBHp31elDOA5QChWrXVN+mplNf0ItHw57dlCA+HPtQfY45T6vRlfX6n4AKbW15rcb
WmVrdbN0KkoCnU+x59gjKCU0JeeRlKZFkqGXf3+yITHlZ6kdJSUGg38WrzbTOyH9KR2WWLBC2Ij/
AR4cENnNrnZoyXmEDAflKm06qJe8jKuTK1JC4xN7wcOSUEYsP5j3exwvaAdVBhMi3sYMmGSFrL0U
ojeRXcDC3TtkuA8d75cFk+MOYplRp+IWxx1zaTg9EJmeQbpSfREs9GXJ/PB/M72/cU3CqqZe7G7a
Kn4nlqZdYcVKFJk9ADiZr4aVuSMX60g+PycgdeaGeYmgctAHPBXWPd2N5q1s8J9Wi9MXnCnly8Jh
JeV5T8tmCl3CoiN5lUoesl8LOpqSVKNaDwdofZvYrvNtWVutNesDxMxsDiiIjs3slT72n1wkXoER
pOWU+Ae66dlTotG3GudNOSQEaKdDGKUtHWkQeSayqGeS2/VyqUlxW45Y5j5AmPGlyqY3fLWzxxgN
ZVjVeqzUw0ViqzOXgKS6+9HJZeMXLhzSJjXLdCjOjuNwSK5wXdkv7K3Y966/9JojidzL1eex0+Fo
iQAXdq9Yt6fYaF6QUfxkpxHYQmY0YNreuomuhEIxxXhJBig+tB1JNWwoDmFMzQUylmerMexX5o2J
XCPr8qiC/YNkztc01UrVnsmUl1be9YTpcEZOwYHlRoHHE5X2Y/GL2ms2oFtUVxgAiP4xf7c8PWcT
mIqIJwTZG8oo9cyhDxADaMeobZ4kRfonnOwJnp6De0nRcniV/NWbg9Rsm2LNPrJgvMa83dR29HMs
3vrlmRKoLzijXSysEECdBlZvIJMZ2QrGO0s3yInwjjIsAq+6f4PoZDVGMb7wnSdguh+HIAQXa5y7
EUI5iqxpufqvIMLIBjWJ5MEa18hu/eU4kX7tDJljpvGb+YpO7yAVnPBX5Nq0EVTQkH1nGmwNGG2T
vEpNxKZSe3RiK6nL2ZINx0uXeLJeYLqPHxUf6gOewpIe9P2tpoOS1t8n4XdH1EwuxbLUlHDZx4fj
NOYNe7il5b6Nugfk1703iS+H/d9AV3Wav5LHfZdLX2f2mmPDRiLRnoWgfWI1XgX739WPwmaTSKMu
XYocny97a3nrZdgR2fqIwftYuVk3yJjTpkoX4OUqRiPwVUYA65/rNPG1+BOI+0ZW6fusA1ZhMKA5
dXj9GhAMCWa6DEyH30IZz6KxZClHvE7q6865NYVoACIf2pRg7UtCl7jJWmIdm2EM01pMTlvHDLik
CigGGQVg1wLYkH4wSYB4twmZ60Nb6OING7rVzStlC+LsCobWPh+aukxb+6aK08GOyZXqZiVZeeZh
Kjd/Qqft1viVm7eIZlo0JCSGaRJFrKe8vs60+gxN/iPduevcxzLaEVFaMrQkQW0e3bvA4MYfxcFj
fy+3QiL5nf1mUad8GafiDjRbexDK7iIFa/vOuy2eOTM7FB7S9yZcVp/6NRR26NNEfAsa+k8EMqJX
rq0ViLIDBhT74MJ08e1PwRqDJs4cxh6m3eoVgoGCyYOmHV7ElVyFDMBy1fx3sO7E+DrYFQ9+Zwb0
xnufA9nI/3ZqPa4HPzCB1JAFv4vDEgY30xbjDuVfK7S2GWmE2cLCmo9iJhoP/Zon8llFywjZvkcU
/YHs/m04+305FzPudmmCYWpc4tM6fmBNuZ+3bX9drT44oNVMtSMk+5E55FO823GPlglmAnm7tkdO
QxdrJz6cqBG1i+oTzCP9QnGrCoQNYLblT6F4/DM5HKuBSS3gew1lRrQ8Gl31ELMkrti2FAgdJsXM
y3pyPe2NUPHvwgfMym0QiVLtMtTFwk3CQqLGm6ZtrGnpmL2pW7EU5BkD1ZXkVm26ylPks+gj44e8
I5qJnsjbcoE/Xt6lDhS+CkZP9fexnK3uiHmhS1pIh0gTwUJOMNGY1Xytb7kJduMf2/tEjim08jeU
2j3kQEzTCUZMoSWS5O5aQHSH0oiBA46llaECA9GirfpmKtA0jASSs1prnK4Ws8n/E8Qe7SczFvPH
09oXj1Z4kEov/xO1L5ulnDB36gX+VldUCn7UfMeGKosE0JG9cC/G0JJPBecoX4bI4PoGsK15Mn7S
lGHufAhSRjJRfn6VSlnuglhOmDAAJ68RUHbb0xGeDoZYnfwVsUJ+U564Yede64oub5fWpMgdGshF
SrYmBThbSFhKDAj4RN4sbi+0M+FoocyxJOPmMU/mjz9g+Zb+2TX7Kv4ZyNM+zWx+LY6jjgewfRkY
gFGnvglh2wdJOEI4F7z9qCorEsZ8hb5Jei1PMbdAbEwy40Cs6GQIyurdnLqjuLK6vGvTuhq30bpq
K0ioYyJEigpMDyJsPdmKK1+w4t6vAEo2sdCSUfKYfybsAZBRs9UUjnFzhGgiPkHzk2R4ULtj28ph
RbhMR2wgcZ1gs4kUv/UjORy8muMuhMcDb1YliZcVN2WaLmJeF6v9iwHK9C7lP1p7gh+CJuSBbnEE
/7ak5YlO2i2QoUQ0iQFU1cVRDe1cgdDgMaZ1uFQlxX/C6t1Vwu8/wJd1CU0ztRGTK5MhAWbgnpDg
gmXBWoeiRhunWm2tLFKl9RaGF2ZDkL7U06941E5NcSFUvz/eIvDcSINjfdvJ2Dg07ty74NV123cf
UnTz6KN5F5oYet31//EL73VKQCCMSkiYZTiGRRI/+RkvCzWaohsKCvHsaQt4eQH5k90UF0Zn4ato
ZyBJ/qdmGsKRn0nk1h+W1cXyTAvFBGlrlH8HQKSDvQ7j9iZ2MNJB3tMbhJ3fHYF6RakjOgeY6wxz
0wq9LJa8SYEiDGWcoC/qulDb1tAV+K/g/azwLaQckRFtEFoV+PlMQv7oM+4QjxZGUDqgoRcIJg4K
rnMP2TBfhZEFXfsFqDfeaCqDZeo2tbE4cnYpaHauiL8M0x+5+M4Lx3KaXMyiE58Hz68OqVbEnYnJ
K4QqtC6VPyEOvVrMrzGeuxb5f/4yrEjmkOTtWN20flyPCcN1xQu8w7vPHTQCpdksBs1+6onwnN2Z
4qOEBoFUb3P+uyNDsqKebdryW6eOuIHISxHBMtRtQWEOoAF2ToijC8VsbIiPXyiLeN3jm2TszlcP
HzBqZkh3IjB4/yx6z+E0UQAUWMR2SQ4kQ8F9yP4vYRcvchsRroT5MmG4zn/vPNTu8RNE5Dkz40gs
7Y+1GmC1ZX3hfGTWAkmnFlxCcrUTLVDhwrtI3d0NTOVayyzBkCKi+jj8vCE8kmFibs3Y4Eu1TZz5
6P/DR2Cw8tRqTgd0XkSOeMDJIDa/hFCPMqSmZ29YlFK4c4SiXyBf0+bCNogK+bFn/EKaRRh9PraX
5F1QQYr9D1covNwHdnRZmRjP5rAD/bcS+pvJHiddIqRaP3jvHAt8sLZc4GjYC6KpaQIjLpbXpZ52
MJziXw2X5RFEc2V1gZXSn0t1yPnZrzxSCyvHaOLuqODTM5iImE7LJuSS/w348h/1yFfNTMxFAHU5
wOk1ndE02X5CWkGZdzH1cMRw6tO9wV/SP4wxnzXGRVltt3BuWtffY9/elmblsqyaqF+Z3RyKk6X2
Cegx+U6Iu/2DlBQBVXdETBoEX+rJKQZh1MJtaYh81M0HqqrBIFcxS4wnTZsiZ9hofZOzqT3FCj2v
PrjrpIR0v+ZzDMMCgGPCOv7djMWs2bU9L0fgcZcoKRB4MaWhwEYzIGEipP+zTSTZX1zW6nzL13IU
I17tfA0wQz8qkWXJBbT0aRUNU8Vs9/CDAe9IZFrTXvyI9bE1OsGRhQSNiFRmVqL9A7gTztv0Z2D6
EuqudeJFaz8fEki6OR0O1eBSxlgdLCrpmQDwlQKieM1o53d/CEp+M+sTHj3/aA6J5y+QXkrGOdiS
tRANF6M55tycc1g+YnJqhipA7YynY309ZRWiC+lBGH3mMsAn5xckSr48+PpEaL6Ugga9LhpCEXTE
BW2D6FigXdpPnZZTLqSlBtGzRk4xC08ag97EUDFlIj5u7OJB58CCBNNpa9ixnyrY1DvOqnfnk67E
g1HDpFtiZFP3DCr7F6sqQPsDVJ/DsNi8IFg+kfZAPwXk36Ntz7qnEOb5ymd7L3CuTLe/cWQ2546E
dBhOaEUthXy08N4eeAiiZJSdxPtdFr1QBCayu4k7Bd5wx+0EnmGWKON+1S/V3uRQr/nbDAFUmg0M
bEhALg3xBDP3ixV5ZRR39sJEc9Upcvqpu0efV3RppXMZvOx+7A68mZHa0IZi+0QKWlMlHcjeUJ/n
w8VsYeS2mGZwHWAE1B2D2I+ZcF/qDI7+PdAY90aDwd7KGGf6c1QGxaK1vb79Ybn5IafHuZPErHv+
/sQG4AebvHS8xEm5E6hJMfN8YweNGZzAitDhmuzVmoZ+QNi8tFtI5cRHTSxEeIl765bsqbj74MqC
bSxRCPabktNmHhX8cvF2ijDYsrwraRoYyvNpWZYN8P0AS7aJB3XumJrbJ77SSjq82Fkz2k9LsKFP
wtJmoZjvSnow9kIV6Xu61KJ5AZmUQyig2q2xMakFnCBpaAJZyCWIC0bXkSqgksQW/MrlsJPLAD2o
rtUEXqRgdOgqRf+DIvUY2EkjalbhppADMhyJpycsIRdZYDiPapIo9JgYh2L2GoS88PyvbNtTpGAN
T/uaW84e09CDJUGhwbwGFK3jkcMTMe5VQBIaXn9/dmiQhuZT4P9tdIHtu5wXd1UW6EtxZnHTjHSL
V5PQYFvITj6HFjY+qVcLCxiDcGRMu/ngKgNccAlby+1MBxxnRxC/BN3rkuDmw2EqFg2lNmDw2Z70
+ccvu2nzVNWimxEeSF7RfhaLRST2vt7fgFLjHnxikTAj564BgVTJdy8vzNwxHVXHJEjkU6VC2o5H
HQlkwII0AQ2t52fu0LKLkSC/YcZZ+DLgb56h8hVNPiJ4ZThvAJny0uyFURF3JVZyo+Ltv4W90qyi
0JHnzsp+bIKLC6jPrAFmOd4/3KTX4IcnTOYWx9VCEqCWtm+znrChcxxCiVubEUI5vTZo5ExZWPzD
5uoPmvPa2fkHezB4mjAGScL/1E7RkPI+Y3mbOSbhO8Enu4SL449utilF3/fm4V628Rs+wcCsEiOR
GnM5Guqv3fyumCRXvkDWrrTcjilZhogY4qlkswYu30cWKuM30DMd+auZICgrijagCmzKy2bnChr5
zSIbQ1S/LKasRWH7heK3O4cYXdVnjtkBasydJT4hjHe8RNmyrjb2kRlLm4NHm9vmbd+fjKYURL+K
HukRGNk50tz5jBAIsKhp02dEn5E9FZxQ2DoCTy3jBIF6VrGRxcaeRo9riJs22lZJWQwwKQ9iBWTq
wa1KgxO0QUZDAz5Mwbs4/1HXlRqss6MgmHRd9aLwtiPr8hffm8CpxTkKYnqDPExMfl7ELrvrmzjT
/A/1hXrYvdua9ds9esxBBasPyOxmV/c3DHGdh1dClud7Vmy4WhdY+iOdOEkAoF1Y73dBw4I2pi5r
sANSe+lMOE0D6OKNJ8Aw53SHnWgrtttw4BY4oScUkWybXBWFPzub5y+MMtUqcjbT7tuu3UU57WPg
4hZqZxAWQQkszRxKN5gSaeRA1T9iX+gn568leROdYWMu8EhpBaPx9lI8tiiyA0GYXHUXJf1klOzJ
JaZVXxLCISHNPQOTT+QTkJLs/Vgp1XrEWztrAO8hjde+7zMFx85f85naHtB7qv1zoaTNfCrNBVwu
1JdXwXAuOoDQlf86m9b1TClodPkGFSs4q+dsqu7cv9nQ+M6aUxxF0xgZwdmsEiXHS4yboWR123uS
Nk0GQR9MNOyoc9pERgHfM93kLJDJb0Uih2rS8bh1GwJ6oHzlIygimrDiYu23U0Y1Q1cfB47Cd0Nn
WfyhE07zbslD2gmJAJNdZ/GgOaE0U4N5ZQs1WXbRSv4Aab90YttqYjK4FqICvUUiZuloEWD5B1dZ
Oa8yQOx92iXjWvk8MHKqYOJnnux0RgmiQlcxk4GHxDnRkMHn93OFrlukQ17brk+pcUwgIf+HCqa+
p8xjoPp334MLiJ4RKAFZR3ho74x2lKFwXKlsQbRRlsBcBVJDiN1hlXH+7uvws5brudT+Xni4gxPz
mOSKTXJzsW2FM4ePIr3C1NiKhqCBPwl9BPJeQiAdqRXTxBCIdNf117jueejxxlFc8V+CVCJNQLot
l55aohvgqGTmtJCcJKdiI+G4k6509qmo+yB+5IwMiBMZla9IM4Tuu1yZl8dmFIAV0rCSOmrEqG/T
RwHGHUxH9GfC69BBkM2xpahH7ASI+0yXgDcmwx229slEh6iI1Wz/kWlwk4wUucRZyaA6L0oiR6Qt
PYlwyi+dLb7/vZp2eIutp9we4zIk9ulY8XD/J/SiTYme6KUcpuKiQVnfhgrh5sh7kAxH16I/9qMG
/IQGhETRRHhVHe/JTImGzt8dvMgY2+KX+ENSmk83UlJUQN6xAe4pp0o/T+H+6aDId8VqKepe75BP
qHJtU4+xcXSucdlRI1Zhq7pBHPuferd5yGEt22o7CZplUeHig1xPWRVfzU7SsKG1DsvVOIy1BAQ/
3QJrONSdSgGva9xrMgmKmczP6WkUnUauGKFVN1WKcCBry3xEx1qpn9T0u4CUIiywc4BkTQC3tZ34
Snh0tFH8iWid2ophH/iUtajIq/qa1SpBWWDYZZZPc07SK9V6lV25PyCUkAU3KmFSHW591l/gp3ex
l0ccjnEc3m7wNzII9YdI1bGuV4oI8q/Br8HCPt3Kb0UjSrkZM6h6grirg4J9xptRuwo9+n91k6g7
VQpH9iJaeB+tmVMbXHKtAUqqoohDql49S5gT3hC6r/ARVqnuKBACEuturUApWbZGFXMspnlJFJk/
0rvsyAYzZpjoZnNm0M5MYM4DFRL5uFqN6zmA1dc49kZPSvUGpt7MPgc1uY1aSvFYkFWEZAw+T948
JUSyJ8QrUGRJD8lmekhvRv14hcvAQWkFH2jaHy5RlX6K93huEmHpEdG/5rbraFyxdkZuMid8sRvG
o+IVRdRlZ/eUbLGT7M1Y5kSGl9h+40ThtqsCbWLGyZTGO2KKLhnUJGaDZ870g340Bohe8IW0aQK9
GVubOLd3TTUMSGIpCQ2s8MlUm9US2tOg/7Lq2y7ypYQKmTdpE6ab1xJWtAjwcQD8BqIO3aP1pIl0
/wo0uaDbY5rqhZ9YQql2/5CKgPgQr2Lrd+z/I1oi7aGGqronFjbvloXcoU7H/Ke3uhc0U0cpwkZg
KSSClnTeeV/Nh8XtJQbcwMHoewKfM0gga/NInpnQsjGNgFyviN2TXElBoVt0/fAQvnubrjq6dyK6
Rj/1wBd8EaLr9I7AQYFoImLj1dya5kgHtY1KQ+R745zFM0dUO79uwrJYJCcBcz6LEbiqrlxWgyjD
FD0H/adiUDS6B3sxl0/BWHaN1FAEHjfXdA5utZZgSBZVINIpJKwknffJoJr1pwjWA1SSue5dOoCY
3GYKmDtRNYg/ysOIO6NSeIT2snAxlyus/b6SV+zR1aCQsyQjiHlJXNPPfUQ2diJObBfeWPysQva9
SGl4VVQ55UyA6Nd0PIEHqmxI6Y71eX7hmO2vxayQGDYYaxRYu3Of+9BL6Dmwb7VpmCOI7hHOcH40
YlhhhrbhbKjY7xohX+5rlMKm0KiTs2Skco8ufdq7Ph4nBVdt7cLzANiiIzE5ZrDvm4YebEyNUy3G
4CjTTORGFjUTBVvfenkSw9M5SlcJUnFCRRhFgs/gtrSVRpyBRgb9fRMEJcfhoAT0f07SMxwMESTd
slR3W7VGu7+Btx5EVYaSmoYTs8uhedGqePB4GELAYiKzVbtXGVUzh29Fz7PFcuRDJcB+1Vfmg6Cc
8TgsSdY58MUYrNsE+x5bWEalGDLKEOLGsXqteX51QieJZAk2voOeHu3R7VsOHnDt6vC/FyazQpIR
KtFnqUHkXcWdDT54T29eHzRUAM/h/W+ISNPn9zSYiKEFyBCL0+86eVl3KSGvaLfQeKfGbau3t22s
tZKsfo8SL49Ozft9Y+qW9AlAg+9KUDcU1JAjEgHT3/ZrE0EA7wURQangbFuxOK+laF3ARta8GbUk
2BzIH08upZwlBYRHmmGpTmQQkSE8DgMbpvil0r2OlRDonQd5BRRy/bbdBSpoBfyxnleXdMAmI/WD
j52mFlT5cXSWOIWfn220ykk3mcfkiotWDMsPhhWABaKAvQvD0K5YvU7Thrzw8r8NO7To7pfGVOXd
Z1dzRo0wd3NwebUO2Zom5dSzzT4n8ilQraa1qmBX7XV1kreLP9ki49KEXElq7px7VSZvIZ/6HVND
/CcC9dZXm4bXC4m/T3aDVBpwoEUNBS2eFwvfqkuCheeu8nRH1L/RGxkqSx8DHeYRMlMU1O34KvJb
93wgI2G2ELajQkxpUpCPZkxcv2Et3bIz6OFFILuHJOakvmZadm9QvD3m4OKIvJ2mPWjIuwYx2Bf1
tZx6wh02T0R9dm0Bao1rcg0t+YUrPtZ0miYkUCP2wVGqaoYRwesoYMLdvELrDSgwpDNdOH3nE/Eh
PKcV/yobZXvXc8mMolNS8rYnnAeBqh2t6Zz6bIrE3y40lwnbrYjny9HRLMdygUgxlQPSCmzsNFmZ
m7q2tX351NyFbitmrALqZeKOsO7sUf8NZ+K+lRMssCWxt77pdABgqht+Cte32bG+DDoYQ1b8pSHS
Bbln1bFJ820rJ36eleDGJovy7r03IBDns411S+exh6VvfpOvPiojn2IqJKrEsiEijYMbu8HTWUsM
Y97Iw7TP2nP24WNWrunxhgmL7OTdsg3eRL/btEQLIUIAgVDbKzP2Fmd+v+ZnXsLeMABCRiaIcXys
HE0htxzkUvxyp0tp+DWzeB878UqTabQ5i0a/sjU+nf/2G3hyhuvznsYPr8QWBfaAEK61cj/EYj3H
c8xJzddKrM0TgnyrAul+xsKHsEzNOmPh+43V7QVtQ+gA0r/QndxuJ3A/bIyE70ywTPP+OSo4+Hkj
AnF9cNDaNcGcYUiHdhjlcqruNczAG/Z0R9shYVM4iUQuZgcs9bJNcFhgvWnXVV3tNzKoCdfj5lrj
thNX7ROlj2K2PN6QleY6oinwmyM5pAnnitxynlyUBFksf0dI2463cNpllBhuxuwy6p5/+HpZFzdo
y58mw60Mf80MWCOrZ7mD8bbSs5B9dVwR1ouD1GQGjNlwwJ70Uiwvh59U16hlZLSa/4e1TeJoBZg9
UgY1COmkMJP4rHck2dboRLx81sGhCjxgMnfvBoExhRrvC4vhyH/fhLwUyTx0ZU/wYi1UehSpm17t
7Ut7wyrjwqq8wDVrn8PSKqNTbPnc/Of22P1CagYsrx4rhepghzUep9oAssQJVGCUsCQgu84YtgKV
MF5ri9Diap+jDkybOZNJKkdAHV8y9ufdyoHEgymrEuiOV0HR1L9Aoxp5PgI13q28ZlwPZAob7q6C
Rwzdo5pu+qJ4+8CybUJUZwD4uXglEQkgaANCpXuiVnQT/6acqZDrm0pGg1w5utmRE1ESQr6RgUwJ
vozbn2PHVnN+K+jMoCwcFZa38uus5BWj0lfEmbZYWDvJnT8cCdREk+NpFY2EfwAok0G+1arMVUg7
pXRknrLu5S6X4mLUw3BrdnHV436XoHZ4Hciqh4A2HlKfs3n4/r7t8Cazkhj3KGgVLbdCoYNrWB4e
V5PaVizSNv0dCfdo8b565cdJntUAjYOdeGdT3wL/Km4FNimSi3//coK9J8xA+1UxhPUqMFSUaR2i
BlbMj0XROqvlFUHdLUcaZYLNX6W88cfyVwdN2wB7iutsLfMBZ96S7oxyZ9vElyQctzX0MWMw99Qs
Gx2a+BSQmO5/BydOGEkIhk2Je7T0oCxedlGPmgO4FwILr6UtJ+j4+1My4ythFD70U4jxdDk+o0Lr
V71zkcujhhEEiwTPqeB1mbRXAxoqX2efjimsmAUQbcLibajvJsVOA307n296RX+EnpU2ig63CKxC
Ca+HjfBYlyQrdwof1C64yBSaH4yGADjMLzL9MDB/bl6EpiZVp3GCE+Y20WtSD6odDXHDOG3zHkoT
HjHSkoi6llPBf1R/Zx0PUr+GEkgXhxqSbSjmjRunYpiLEWyUV7doRErozlJnf8YJsAsJok4HgEP2
MakHicpD71qd4SBNLpq9khPq4hhBUxVHGXHZK+VeuJ1LQmDO8JhKjKQ+J7b89OG2OblcTF+N2DSU
ffCifNpP/AWu9ev0ZYzxpuHZSBVDQ/ZLkPlrMbPQ1q411KW1pjLsXaS3i3zKuFG/bVRlPFOC08M/
14bSl8wR0NB3wNRGJ7OG9fBNz/uU3hjTyD1sAFqHrfSExdZ29unYgwSf+X5OAGSZTMnzRR5sS91r
5JiJBaXcg/YPt/HjKWWpHMoUjKsEIF8tSpiVa1PqEls+EGaaodDbc6I4YggXSiKMcv7oVdLxBsGV
Fk4ntJD+Wbf30rlbB0RazFtVcpPkxsKvvW8u0uv7fi5+039ZZjkQKO/z8SrHHksgwoSXf8jwr+ET
BWrqXm/HT6F+bR+ZIm6WaDX19NF0HHYZ3jmQjWo8quNwOuYAjFYPvLc0sT7n6L9MxoYb5qIzOJCh
6oXRjLEaAItPzRXnyHy6W7etseY+Ht5PNXKmwPak/YW/OaHfamm73o2A/p9DigxBc2klNpWeLyFU
OyhmHJjITBeU5VmuDu5c5Kwbd4PwY7O3nOjwxKJ5JrD8hBxd6lWkgxfh/e7b9WT+NBQR5N1nQ7Xc
wDy2rRS/SSFNzpqfUerw4hEtbbs0vGvmt1I71pyEr6SsJ/EdnON7VOD4y6W+xCgPNoxFOVJQ/xBc
qDcuLg8ta2bJImTwabz1x4/7xSydf/zhkNAZIBWsFPWLPlaTMlD+oTgyxBhecL/94xMIXc8RK3Jd
Bndf+bUnpJ2KsOKwi0UtpWwE/irjVhJt76wboPT1ut0GAkI+Or843B2Y6e4WKO4WEqWdJJ/3FnJ+
667zlVd/yQJvhqUQG7FU9y2N67OHABEJPEVeyVEaOQc05Mktm/FY6ZPil6XsNT7y3MnWHobJDXIH
p20u2QHxm2fpDM+aay3ueKDl9pvyKpV4A007Ozn8DVMrXust3sam4hS1zkVAuxMICKy67+VJG3zk
J649/mUBm7Wi1ohZjjEQlVFJgFPgeCE7nj7uGvIToCrqdGUq9hTw/289TSsAM/7lSygNj9IJR6wB
JRNrn0Chk0+ZdA1PD5tuof1KuF3p9jMA22VeTE/9+FU5j+SU1Pc6KtkY2kbLPDbKIXxspsBnLQyu
n+gQYgjofEMmQ5zq2RUg6yu1/fhiaM9zA10l+QAR2SnSegrypgpLnckoPiZX5/CLqc2aceqxg73e
tp72fpZVs0lVa15tgX8H2m30AfxYE2aNtNnsnxBYcl2KRVlX/SB3of+pNNkYj9Qsds00jqbkXVbh
SXGlgJZaL6nYHUyYH9Qf6D+Gn2tIBhoFROBwy5NF4s0fVUApp7kgpnJdFJc4ZwRTwV8bsrZRFHeY
HMwR7v6IZFqbTYQMaKnkfKSSqJV5wcDj+U/Vq3LipTaCwf4qFg9oJ/PuX+4UJWdhhA8VtQiQFxrX
09dJf+OxyYYHhbfyxe5+aOI03Uv8Q6CDNvrCtyEr+WAq9j8IQL45mjcIZ84wXYB1d31jj/GNDCyE
Kv9xcu9gW4mgjoiofCaIKfo2ya+pqRBwyW61sCLc7h1ZCABwZitdq58jj9UtPBM+AlWxsAhmwyxI
5qsOZgOFyKq3EH5uLmD74wT+HtI5dnfJVPzYHC0YUs/hdX2dntcpiX2qU5XZBq0jjGoUzz0Ec/fN
5nPAtUwTbiy+U+b+nFm7/mjAMM9iiMC2Hoy70ZyTZgMKrDZE/b5zaTYgXLoVGrZXULjgIZkD4ijc
3CodVkRIDSyeO6bI4PtQr04pRhlZXEVq8tHkpy/mUQwuNrQyMMamkIDX1pFM54X5a1LBbITaXHlC
cE79Isp6bzH3+xUSL2IwSAMLcvId2nTdYu5qTb3kfQWjzsZ/wJYKIXqa6mIqTQxCQiaz+eZdbzkP
6h/h+cAdJET4VJxjAURqeWhCJmCo+7chtLlWzyQw+AUAF5JBcdOjMnD1pcrxEm9H0xLbbB5Mj0mQ
n58VlVwkJHUmQjS6910OtPaBTTH/h5xO0D3zixEa3OQxzvrgrsuNZIaesKFbNxcHM5w/BufvCl3f
uiErfghi37B52yPzipR0U8aCWkq94f9Z7ssXJXOCFpqVE8cc35Ks74ANpeDDh+JPpF3kgc7BBzPE
YlSGtJSFu0BKev/VurzaB5jeKRVD6WroukdPzV2vgzAwnFpj75eKJoUUr9wwdZHXjDXw8mE8j4ah
ApHHVTDHMBJMqnwRO89onyJWB9Z26IOxrhMUfiu9rB76PZqQGQjDz58gbqgi2JBTH3jfKCxpbS1r
CaEsC6Lihb9NMV8sKo0Swf4ldAxmaY8MYhMLrMge+SKC4RJsMoeH6CNOf4uw9v3/eTtNjuJdJt4b
5WQOSXbFbVBQcqc1DbpXlCX3XadeUFxgrG2nLnzG/TO7F66/G7MgbUAC0CXWeACuyWVuHsCKE2ol
exoep2BdL0n3WsNvnzHc+in8Pa52IVCWXxZqhjAVmiUVD0Xm9zEmvtlmgiYklIpYMDffhbWgD2wS
MB3v9cUHl6zErUh5by+FjqvBgYh854gSodcQuH20Bj52fBG3UgB/ujr5q4wOA2cIdP7a3o+fJlsv
k/hRYMEDiKfJyniEOtTeBjtllUCwdSAm2ULDqXdux0H/s1yaCgLNWdj9lof+bC5tOoOn4X59Q1Qn
yvEpiMsuK65XtSpTxiTayunKYALTZombIH+DH4rWcdoq6fOOtlqU5OteA6CKYtl0iAZnsjMqaFuY
D+q3h5J234gnnUBdrsBZNC7yOLMplxi/20/tQ6XA042P82hf+3nRIGeT6LnLTBtuaBX2bPHfOCwM
xaEN/GILGH8Hrzj5/3Vu7HedujwMb+6DtqwONCLpcpR9gbsq2YxiM6OTynWgcqCeBMAw+woSUBKr
nNBr4VC8z9ALsxGjRjGBG/mkxpSGbgBuc8OqddNZ+0ZurHqsvmmCHZ5VN4JIpOt3y14v9se5w+Of
Dbuo+KN7qiVKXZUrwSHszu3k5zHIJHwIjs7DsvWBFr6IFYF9XdxUQ8xC19o7+muxPLEE70+YlxGx
WP9cYRCtVHM34zLe9IslFgQQVG32LgcWCHWaxSrLrm57sc4jml1rOJCiTlDput+DYkbL3aPPaIbC
ilzhBO6i5feHKwx8juckaS9uXiJ2G0MR0mpCdzeTcBar8b/lj32L+Orc5/BFrJdRLejSu8Gk7iY5
13Dfqpn8E4gqSH0bZApX+diU0dfyKg9qszN+4LM5eZOV+biDxo1dvI4WdRRw2/cSYG0C3wrBe3bM
7sf78Na/QsLAfVrm6HSDvuk4JlIMON6L0FzybhCYKqyqGTsdZWgWD0XY6d3fU4hApfCAAIAFTjpM
AnnJY5JSXOIGJSr42RmYdDHb1KGy84lbnGpyUEoqkfTULfYgzxHaThjSntgr7/IgdFmnqGHpl2y8
oo4crGiVTax2+FvF2QoZnNZfwPR07pv8YCmdwbYiRunt1UGdw11EkpNCp5oUCfsuleCzd//TyFri
rpJmaBsTomuU/KSwTzpQ4kNDqUzV3j6fRiLA3qgXsrPQsPATWAgTv3ltMwGzxVNsOxd7n2rX4HRS
XBcs+z825Hv0DdSgSdKuBNM1qXSur89287n6+n8IWCJOT6MCHHS/0uJwviQdZdUwkornaIH3mq9v
GU1j7f4+caWT/on6+ybOgzuyZEuC3LtvuqqLtu7j2rrgHTi2Fcjs04YgiCyqem64nMZCEu/NC1Ud
n1ip+agrwOHr4hzqqCmqgk+RWE4YnkSz8Y9N0t1fCaKoAbB7OqMqP/GBeaJtpdGAtugne01CL5wo
vFTZ+zk5SV7MDhoW1ksghA1Q1XAl/xjKhqiR/t+4qjElcXdHJjzu0k2G7TO2aJXtITygu8NIcCNz
xPBguOO+3ID5SbfpPT5dPdiPqlMTM5oQEceL0WkNOfPkS57oz7lp/17uNlStzDrGo6oUtB/fdiqI
7gqoZpzJ6HzreHqxcVkHWv7Vcfe1GqYZ51vxvkt00hcjwgVcfxhlGMKHY79plHsWB+l78/hynTpR
Mmtb1XGirelTwXlK86pmnkGaGbCMpUQ48qWtOGE8BQ6jgnWUj6Z57gYv9Kvj4pjgYgL3Mu8kMUV+
pKP8y2uoyYXjsiYlR2TZy/vPXbz2SIehXuyzoOU5ffA5eYgxZHkZMqJg0giZBRinIxJ9A0Axb3YF
4QwGzUGt9u3KiBB4w25V6Dhj1Mmx1Q1dgZpgIntW8zk/xJg6tkhINRolC3FSbjeRfinipKggXuN/
ltK62I1Dnzx+NJvvfZtPIxiCQChVhjBz9P04qqnYCK+3v7kow7ll4cJT48bSim8Wt8SW9YtpOksx
KFzlZzatD8dLADkkWCQv8Dt0aNb/IPA+NjXNHQ3Lg+62FmC59ouGMy3BD9G/QDUVadqQq3VOyonW
jtCxg7WBaBDE0a9hvlKC6eFvf3tKcDk/bRepCsZFiL9CeidL0MDjOSXJtl6dkjawDuLymytUC4s+
NoclqImeLdITxUGpyGsRQkQfVLwnVFqYVScUqJzeLvHHKoZajN4bVX02QLfaJDCVfB4G2ZFE1KFh
gMOkgoIgZxRRVmbT1uSYTCgpbrvxRCPSmaVfOosM2uD8QCAjySGtRQ+hzQ0vXNfyiYQQNPzaikq3
HRpOl1iWIR7Dj027Me8AQy5X/ma+8vkMoAACsafvgGcnS73CiudLCpQ6dhtUC5k4Oekf6FmqIiUQ
A8anTTXLO1I/ZwIls0pPcXR+Okq6hFVLtELGSt9LNoAzBecbCItLWm2FzlWv8KxnOtSjP8GeQaWG
cgfnayHCwyi4fs8L1LEJSkV6xmu8GRXBLps5BKMxozjhd5Mayg9srV5FSJNCcWcHrRrXce3YVu/3
MGcw9ms6Xdw6kGR6Ekf+8oK3L3kWCmAbiBs60kVsp4YzDgf1V1AaHC1prpWl8e3pYmM3gmSeRaLy
wM95qTRIc/LHqeFnU3Phu9fSym+YSk+mIbn+gxb+XvrzMn+U72qaNtWRHso9gXVCsXOQv7nkHQ5z
AAzRURZTB5e9UhLXVbWZs78gO+t1CKoIepuyeSleqzj9nx8rEgTPgFVwwG9pklf5Hx1l7NWgE1Y6
eGbaQvDDZOh7gJvgPu3P24f9Aaa54DfW4VNMwX+0+UitESprf6D9XTbtpg60vBfetg+75x7fihaT
QTaBmZQ3PYnqMH8SCV9uhUwbYfx5+MmBA7nPleTAqNhwQszi+qOpG1tvrX1wGgheoEOzzBuAtHC9
Dvfi9Clq+izkDcoIGHvHojhx5G3CVX3v+nl+AqQCGZ5FJFkwV0+001P3YEgG+Y0TRVlmBvJCH1A2
LG0spYrKLPqJKSFuI4+LHmBg9F7Hh6Rh8HNbQ7xUTQrSckBJv+fiD3cmGv0B/9+d0es9wTSv5qrX
+y1uQNcHON4FnFNMrSp4FpSel5pcsCAw7z3htmb3DIIkQpy8f1AzwWz5FRSfDSKI2DFmx4/28FS7
mOV/MoEc+gBaCOwT3cJPzKuWLpz0lMOKua9fajXKH7RUyalWBV9lf27DfIbKQopZ3iQJzKO67iF7
u2zUhe/lWMEs0xjExI7NytUdU6P1SnS+6EAlwlgUCvnE6My5zu5Q10eOQgfqdH/tstQ7J6/x4Z91
h7UZ7fw0yN+L/AJQo92jfx1OnsROVJZfRQpJfr46fiyqsL8Ti1FCJ/SzcyAemuRFXTM2JyWSSmQI
Ii0FX7ESF5W7Wg2hrdPoaoCAYyOiKE6ybhBG425kvRil0+zuBmkmwzgSKysoku639cO3rtS3mnhi
AiP9fkIeCbDWNrlFLgYe3LvF5Vhh5XaCHhe1kVT52LKqpqQVCI8ZJt6SHIscVkfNK6NhhUI9arCO
V6TjcgF1/Tns/mKOmLqVsk64Yh3WE3xKKUsIxE1eRqNQlBeiDvzTTqJHRxFD3jh1pHpnOVBWvkMU
c06r1JijqEJ8nzOz9akrYOtPs7EVGNenudYm3N1OIrKm4aWNGFTP4oRhCfVjNmw6/5Pej2RCvqZH
jv1XUeUDL9dvDEmWth/R5Q+Z2AiplYtfMMECyarOb1wpTzIUBsl90AUihtY2odkPB958UkhR66TI
dpFp0SG2YihJDPgw2mYoN3igfMYMsHeacGYPLDghbNVIARA1O62F5iNMJcEW93AQ03uH04RtvaO/
VOwFBIRNtRTGkEGpBfkFmhTZClOnx/Zb9fEIl5XKf2r+Tv3vyq1SzYvdODTMmv9HSd3Ix/EVywwW
AMpkXc4pQRv41nPnxr2KzarwVZtDIvgKsBQnGwjrisTVRaKX4VSijfuxRPV4GJmRwIRD3ngTrI5A
O+Kxy+y8fG+j8DkTuTXBX0Pa0dnwC6gE7Q3S3P/2NWwxpPmFdAKZkb3KD/k2LpqKqencOzVg3gVn
ROXZ7zsg+v1kLq8mwVFrqxy5fgMfaZMDz7QLhGz80enV0KEYJoHQVCaUsk6Cb8kSvN+IsncS2G93
sVHUyNqo3f0Ll6YX7Wy67qqYGhzERq2lkdyph1/Qp7Hr3jOvqBueCjID68u5vjebYvsI0z42WCPi
F3/8Avc2rUyCNi6iifnBvv4YJ9DAuTFRKjnQn8USeEpfb5nTEjZ+pX+1xV8RcYnRdyLRlbXIigco
kAoOd0sa8FwsNH1eGqRlDPrf9lBx8pztRi3vrXtFoupY004pnOLA25yM4mXASrW14C+pE2NmzaPr
nCdUIvSqSLuiba3EQ0qpRsH89TvlXJBp9uxv+/L6QOUymk9SNf+j286qf1IJYJX3owwquXjVx91O
pDPLetazYCqEGlk+vWJl4sN3DFPUmccrFNcpTx5atSAD8w4JI+7IRfRMByJZ2SpPU4HsEnViCsFJ
FJ4wYZvgCBTXZp/vVa7Qwxt/PvIWM8Qix5JePm2i2A6GC8RBldxzjBHZlKQoLy3ShmqYDZOOpm/O
eDLxAuQTTl8v8sTCx34kCeLc3ZiJxE7lPsVKpygfceFCd63xy1JjIPmDQbFA7U4u5K08UeAapG+n
aF4rKeMmmcIPK8wezREX3/m6lkood7JUMGwVA5kVxsZK3ymmGiQXGmUnTdqmhDPj6COSQE+3DiGE
1WJ2gPp6qJhP9SHVoHUagJJaHUIUQ1DpMJKailGQz16DHMnSxU3Qzf9yjDebst1vzpuEMGUa0WEd
xZZSdttGa3FRBwdwKrg2KJ78LpYVzafDOFCND3sLkcuwu9/UofYPSLcNvz4sm0l1VxzN96ggYRvE
58H1eWRawxExlPBr3v6Js1L9GKH/rU1R4/zdoNWMwmbpexCbxFB8OH7WAmffOwnTx76nZ29VkdlW
CAECP/2gHsQfTLmAAsbEUOwFzM6ajwsm/zSBrzYFd4prQqT/MvSe+ys6fEtNDeYIjm/4qbaOH8hS
/HB8n9DDc72GdOPswQ8GivYVW3yY5Le1FPU02tRcgJRu7F3+YTYSuJ02QMBGiWTSD/1UYJg4CDqf
MPZItDZuJGWsQ0jru7XJQMYhiKICtdFCtb2x0R0yAMjjijeIS68vGsExnZ1zr6SehAh7YikKCE53
WzBgPTX7mNlkJSZnmo8eWjXLLQcKO8O9yuJVdL1Vtsa+p1zbAFNTNROwubpBDe9WyjZVcVturHbH
EZuMH5XeI/BnF2oXq/uD+sdvE7Yh4KalMbG6K4UELYY2DECFRR9X5j4gWUhRwVBJ2moIYXB+B8Bh
DC1QOXvDihPEUj3wu6cqufryzCYNxYVyLkJkyTFFzTNUnaHtwecqqm1BrR8GEuo1k++86LAsUiCw
3N6LAO/1mmQPXY0K/izKiQPQXujN7WU3LEaPkuqqzWBV24FMRJH83gxnnUlA4zgnhsJzfjE2+fhr
FqDtfP5tXT7UiSgyDVN8AX/XNcFATg1UNUXKWfB3v8VqYvs+ab18ZeGfKRRQDUYLa4JxdpwF0XFt
qK+7zTlKqUPD2U6rHcsJxo7RYmVOO3he5rrQ+cYr8nwkw073xcJ4n0hQCarDovliaO5kQAk1IUVc
qPMNLdM3NJXTQ8J9Z4IWKSsi7yCIHXxaK2gsvWBFDAUqN6DwaCXzwIaeWx5JMlzyE+CWhwrKkh+C
ru4BWGXsp6aN+KMfwWOBXIYzswjiHTbWU3q7egTbYFq4sLZGyLo25HjXEHh4jwNywV4/GmCPwTHF
+wXmvvgEm+so/dAdW5wvmIslUZRVZ3ZmO8S4Uc3/rhT0Dd3NetFtc1b7wbmLBZlYtNevU/Z5aXD5
QrJ0dRqo7+yhjz9wWCrmOA8Re7Q0MekOaFeMht5yDfbr+Dnzt2pwvexxJ0KdVqwAnUNA6N4/p8dG
z+xnv+6HYAr5xsMLiA1OLGllMQ3tzJuaEkQ8+nLAU82jype9Mu9Uf27UirRnPm666Og4qCj9MNfb
OJ/y9XRrAf4WV1XKwkZlvEzD5UDPrrHf0ItUHZDKayGcsEXJLxNU6PgH/anCOuHj76YPj4zYO7D0
xeo9r90TIaTsEW7pCeh0IrMKbjbKkv6JO7c5ASlHkG6G7Mt5KY/E2zAY6TE/OwQfk/MrWKIERsp2
+zIjnAuFq8a9QleMztHjsCIPvtDcpfWi7+8CsRM5sG5Ny6RqzYDm7ixMT2gp5S2SF/N4aykgw5aX
OqdprB8jR97hJSIB4uCKQCTrlRL7Rn2LwgWP0ySsG77HmF+HmtIASAhq7C2OvHEK/nRaz2xTRQlY
bMXhOoQCvZot4h1mqX2yzS1ouy9Up6MPK7to1v7D9gBpCZ3p0P5qh7xSxiJUtyOikxwHSAeRMlNZ
E8hLaJz00PZUpQD8dr6I9H8xAyXl+zFurNPYAWaABbguYgw3o7MM78Tw6vrH5jywQEo5J/5Prcbt
D0nCu0+KwLHZwVGxjSJpYKR3EqKu+fkj76M6cE6klXYCoORjjBHu1DQU4IanyGik3IPdYCtvNVns
3WqKYrL1khyIJa9Ht4c0y9bk75aZ+dUuZNn6/tyU1BHH8vSM62JR6qAm1IhLO3n/1sWxjgWWIThJ
tNIrHp9RoshVg/12g4rokxvp0a4JPQ9nPg/q10sAjbv+ZiICfACo9TsTkF3UnzbwevPZOIs17s64
wTWma86I+EK4w4azKy7R0zSAagiaJtmaP9Nw1L2ZAUJ/bQwoHY+Uga7nAIDBp5zQtYAPtwbmXzct
bCL0Uo+4LpgVQ9ETVxWJmexKsOIFeLWMZeHatMcQRrdFNx7UdFdO/rXHRf1N6fWiETzq6kmJv9cD
6Dd7sQghE4Pn0AmkIyMLi5Se0+DjSKg+Z5H4cR43uVs4VJ06c6hGbgkiFg/Q09/5HLQg+dVp0GXh
iAOlesTncbEGreOZo2qMvVcrm7kKT635GWfgL4GctsiywLExwxFChkTOf+qQo/wxaIbst1OEyTyz
uLUmruSIMl7qjFchC9JBaAQTeI7oPjCLb0ibKAmHdYumvHvUfaYaQpWtR2dCDXFrCj+777dwt5Tb
Dlu5ibsU9tZjnKeAlVOdHtXR2E63ZFp0X0lv9KG1L1HJ/NJxHua56Jo2hT4aOMaydZVjGTo2s5ia
ZgSh3nTjQrZe2m8BusO2f6rZXIWc6cOlJzTiDE+GgF1nxRT8GQbDtdbgCQqNGnBDerqGl9kwRhwj
U4rT0IBtK5jdOUBaf0u7qGEbhcDE0akqlJPcY/znpeOq8Lxi5TXTc38KcXU0NhgRY+xrpA4iYs61
vokTG/J9MBG9o9LC4Te07nXR88xKlFTPmIrylgqHun8nFtUKp0GtKyPPLDDJHVkCt4g3N3u9RXAj
xlPhiT3QjzclVYvkPDd606FftvW47Dx1TYp7lN4xiH3Ov8Xvzgv+skFsVjuEP63OL8ixUxYl55ib
uix6sJs9zs5TN60dXHPZF2Agqf758x0l+pfocB+yPoPGpW3WvJnjIxxutpfg0LZ3F5HQP+ICYbQ7
iJMqVeBVH8na6CpRsaaayqdJQXyEA4OGo8o9MJ8aDopjGLL4xFNxTgDZR8/CNID6u1RC4F15jscu
7f3t7TjmxKdBzHGjxX9Z/oGQhvVQm+1+mckNIQUhamb9F8Ojk4c7mlI8AKZXBWI4dCiBfu/g1dQ4
D+Y9dtz9vCbcghQmXpOrM3HLz9AyFGZlmwlXI0ELKrEj40rMMS36bhUwP/KGldF3rXJV+mWq/U/3
i9dUjVK/sSxTH6fpoapR9AJwczX3XuuBKdWosadOsdI7ShO6hR5TeY6YWedg7ifnhC8HoQKddTyp
05jqeM4RG77cbZwq4oDWYDeE6ErfXKP/HcICrO2XW9Kb76IV87XuygrUFrE+NRYv3zIdI2DucryB
n59UdfWXPApmQeRORSX8DMNOBGVmur+9tbi7FHyfFNVi/txgsksu2ML8apK0uZEyGGyP0xCv+AV3
zT73qs3j4A1oV1sZdYOo7csB4m3Q88MFg8n6sfpn8IXdL/KPEDh0hOOC0ICxUNI1xg+Pg000IaRG
xqcar7kDliYsKpCNRDo0pviX/3uV9v2tig9BUan2mwhBGHuPgNRrF+A1dRZdGC3t+OctgAwxZbum
fev9G54bkR6u/4/FbujK/+pu/dqsGPrI2GsyiO54AG8noppK/FKTxj4ct8b00MyE2XkbrNq326w9
rjU4/23qq6tP3R6UW1SXJDf40ZXik7godaW08qaWEJomQ5sK/ekNViw4rvNRSRrTeJ2KIIAB8xoQ
htD8M+mZBytuQ9WPWC3F60lSui97SlpH12x8iOwQ3NRyxwEqlyHTEqEfiteGRi+IurCzo0KtB+Z1
McsBPSiT/w6zC1Xq7uIN1sOk3Q+DOzvkbiMOiGamQ30/xpFqNCjJog7fRkqHs82ylg4JQkSCJU0f
BIhK6ltRzBVbQ3B31lEtjpUHGwpTImnaPTS39tO/NoMnjdQdb3mcR2nmKQQgTLsngVjQmo+o5Ez8
ZSGbmxLUsAU8dSzE2yEUwuRXLyAEwUzBQSf5Zqt4dQTJXlknqD9569/YkEm15/Shz1X15wrCIiVU
GJOS69ynaVw9DnQjv7ELqTaxMIiHDqBNpxKEAIFA/ASacaIscKfVv1+KhvTmVbSRr4T+y7wmYJyp
9gJP6ZB35yNXhlu+rtpMj3JZJsti8Xya+OlZPFtXQvUmebdQHyK3B5Htv+Sq513e8+fXYW2cwlO6
BbtXWPlT7nmlikgVOyhtXbmR+NJZb43XB4NUdc2Kg5HbrlAliBSIwzqaTQ48EhF1dUDMjrsUbvgq
woScSqZHV2W/V3f+inHPDK7YtDig5MxwXVa81lxZnnRIKjV6ZmIM4a9MsU2umEOWMR5SiIwIeLnY
XD2GzhxxbRkEQ/lKlAVfukC2Ut8fPaP8TFFOQW+JYtXjwzRcpzDDokQguobeXPguoMXwcxo+TplR
fvSULOrxvCICh/VXWQgkOfBR7FOnDXQkpb5S7U8raWA8pPL7hgcUkEZsbj6aL0JqWIlMYQ9QkPKN
jHRBUGTFRd31+FmWqJlrLLuduLjEPIt9uwTsoJEmRsddzhYbUbKbg9oNZxxqbD2zH7SK5jysqFwl
pEJZpmlgKf5X0vP6YyC3OmgC6T/B3FDQ2cUdGvioncaxEPORPqDRpp5IYNaLt3ar0JHNVBKxCmHD
tLNQqFtxFjoISR5BS02D7NJNXhsw4ZEZWNlcZ+juEMKtgIP5QusQZ8oJf1kJRH5OAAQvynAua6LF
ZHAOrH8vSWvfvkXVGAT6pHf55nqSwlqpgeKFk316U1ZbZYvyrPP7T/furAfyG5766hxXIEty861a
5H/LUiNf/BN1Vqsfg2g20KOtkoQgbYRg9fksn4vIVwwBUpCbBO8cM1HfC2FzM/h+f+TMzy4lD9Ba
uwDN/2MpaDKDQjRRKS47BqW9cpBizx2wdKKDgBKToBHA1pelY5S92QAtqf7qmXAMYYfMTIbl0CUU
94saamuCeJ0VHsMB0RfetG1KIFYdCUEOA93zvnUpX3UTlonbODZPBhuErWx3WsY+sW6H4B4zO5aY
Jqnn4eV6RAM2LiweQbyFeS2C3KqrAFLlLePa4CfQ1gRuawbM2AGsHNHpsLYxg656j4zsP56sUBXw
0J1afPBFHMm0WccFqrImV3O50ewJW6NUYUMW6rx6YtTGR/9sS/BDFi2htLXI95EbnaY7NrrWEGqT
F5nVdrL7ou8IpgXl5/tHmQY79xyv7Y4Rs4HLl5Gyzk5ihynRY8VfHuks+6LP2T5V9F8twUk3VdHi
3y431yH74/vE/n1rQdiTPTOGcPby3jdmWoE4xxyQT18SaY/mibzIMQuDISMpW2NWjKKFT7mTiiag
bPD8xK+nCWbhWPPUDJhDhFYfOBGp3/V9OhC85BYac2sUqCn2oA7axvZ/DfmPUwK/g7EcPdp6S0+Q
wv2DVcN/pSJnie0PU2B0got/B4oVWcvLLuNXRVdXBK4Q0R0bGJxtnrWYMg8yvrQ/EeKmfgDnl3xM
5lkoy0NOmksY2KH0HnSm9PabMDkdWhUADUdhjglJD0/TFJP4FO/EYlODv7JfrNFeJbsPbIaI/ey2
7QOmsb5Rrhtmk611/VIk+oorTD5cZSh7X4MmmFlAzVtqbNzMUIZco0nHyYGX/idCPLwpkn5Nv3MU
JGPWm8JqBJUVd6wYgLUih69zCIH1bRZgPGuWcAzDf8pPx/d5NunfSHpPyWuKHQ8I5RHJib45Hxq3
kOeaoCTESnKxfGZLDnZ4Yiva4S/y2qsQUReoerHpa2xQmew3A+66QGLu/ghZahIry4YGoQf/4dA0
+T9HmfaNLrpJUIEv2o6/7R+4JKWaYUzhicr2Rm0932SY5A5fvnWLX75fLtNqQYDEJqXmv0ADWSP8
Y3r/3xtA1CHh7xA6LsqAum2AfQJ9LD3+ux4KL/tfyjZvAEqSsS3WCcAVoOBSX4qc9NQYC61ThI4/
h0YQHAJQKNV0Ob2gaoZ9KRX8QPDz08ePfL0KpJU3Huczu8/0cwhlDAYV1qkiXlGirbuYCaW+R5Ea
LD85E4KYs4zgFYgnOxULa1mFr/6kq/rFJBKJw9rslzDXWX2Vf25EJz9fbZPgHxK4M42mpnoVCBHT
NvUHMkwCuMVMRXUmW2S26RikMbxLjXNW7OOITUahpcrUuaIP5i21O+6bk8FJ+WF2+urDtkdXd5JL
THrltDsWUdXc/GnFL+JeH2zzszZYlyWVVu17mr6rngG1DXe5wjJQYJ6SeYvySOpcaXXc02km2pvb
LPmKY+5G3IaPri5Ksu/nTuT5YAAO6tKHPRVhbONYJ89V+giqR8a5+lsiuhs/DJUtYxnxxpccWKgZ
effsoNs+DxxlEUp6CO1iBKZHWjLlr5crqA2OAv5eyPyrAtv2SwWpoA7W/4TX8OjUJxPJKnKgexv+
fBHaxBykVCxoDiYVoMbeO68I5cplhyaUm0HhO5aL06d6GH7m17o73Z6DRXhkp/w6ZlrblY3+PwjE
pRVWLBMfILHxsrZqtv20HhjTiNxHF55QGwYuDNJNKFSgqUbvks8MJe2bvkgy2/7BjqisVyeAfeCr
p1/8JlFiU4nJPHvNMSAmufZ/bydtaZqwVAkzug96HzTqKvVy4m3HJY4QeN1XM0YG3iiMHLhNho8y
EmC8IB2csWs3t2PT5wXW/DF+nVWv/wZCSD4grrpPhb3pVu3pi3cUuvr5h/A+st+BfuP83yGgANL6
kKLXY2S/yRJdzeVg5MoImx9V6MLKBflQh+ywrurvFDjwdn4xTkueI9Ta0Y36/8GgE3y5NlSh6Fka
XBH8aOtB0paLP73ryivITy69SGMoDRoX24LvZtsizr9syOevAI5qiERP2/ftRi6snAPbXI1X1KTa
rfP41LASb4MSIZQ/tNNiicCNsWo2VBejFlXpUGxN0iBetDj/hqyg9zSZqnrud33MQrVuZNHB0jk8
h7ZYGXLgsHzVHy13K4vzyKlX4OsHxXx9WXaORcRO1f/td743/lV1QLjRw77eHb51YNXDdCakv9cB
00Cm+Jw58T+wTfDdhOsM8e0dYLBIjjI9dBUk1e9g7JnOUujWIal9jxTFqOwLuwlr8vOyy0nU74iY
Uaz8pTRFqILWPwnUV/A0SlsY6rxQh2zbf6zzVRUEIEAnnhHWCQUhNKA4941q4TYPWmLqkUO43Ha3
MV87VPDK5VADJCXKR26gJtkatLD6lYmsXj3F2SgSycngYm+SxI/+9GVKAZwu8pJYObYUifjAWn0V
mItLT7Pn6+M/SEAKUSBrD29r5QQrZjo2r7ByVxiWzoVI7UpZAvIiM38/cyJ+Q23BV3HI7pjLnyPC
NNqf9HJi6jgWIBBG5Nyb4M2DXoWOpOYDgFCso0EnpskmPKUmOwxhkyBs8nZfnTvAnNitGcIh9qqx
yuLnthH5X5Vj7v6nt9Y2bB8R9xkWjO4UutnmiLd7RAtXbHEu6DriGYm32d3/ZJZbdKpElI5s/Hmj
rX4Ecgw4FTK5xH5ovf6FT/pzEvpRbJ7oG5VcOHX/gRhoh2UOCxAPeDGJLyoGpAMhlonD8S3cw3SC
G8ERqsLvNzGx5HL7GuDPQbVJrxRF6IdaLmp8a38K8EleAbz+s9Ds7nPnL1Mvpy36iAuiQ2YqRGZC
4iLIyxO5f5Pg2TiR/4mfUhHTrpaAanPoGyNUUY8nvqwPzxLHCvTTvFEpMzYLh8ev0WkJhusyrj1z
Aho6F3CAHJ68/iVT/jsmfWXSFbTIcAk9WJJ1KLFChMnXvThOi5EJFW178/E3+xufhin0wnrpSTVh
w9iYEnONMRrfvJD8YSVFuMPBNpiuEOVSSFzWuusikShDqnG7//ZGvOzOG3pkXauj/ePkIngyKLGa
KJSFqi3WDftJUvZLs3/w2qFU8RAZGP9zHeHTCdvyjF0DtBXi2H5gwuEcfvQankEaJahSOCd62FEF
hfzzIgrgapmOlItyIpURg/Ws6Vs18aZayeQR4tzOhBi07mXvg76996K3+eUY4MlO0Yq1sUAQdHMn
iOrO8UQTb7EDszCHdz2u1sUVN09s5wpBuOlrBX4msuPs2RKAb9U3GdtS/WDHH9JplfZ8iE5QTj3f
QeLBoctwCjRvz1ZzxiFk0gfeeH3p5+nKhbWATR+4d9k0sx7AfhpKs7tXMXTMYdZLeijS8Ixm5KhP
K+/OZV4H9457CcE2M3mEyZBMDjt/PQrkeRIUZTvvBOtzvGnt90LODqLCViMhR6VjgvaqWS+Z0P17
i5LQXb79Q6+XamegvdzxQv/bBFhJmYzVV+01IXcxqxuB4VedIwYREDxzLQ2p8CsnT+dS7fKhHWEK
eN2Gezh3YFkmHDkqTh+eXQqeglm8kf2uD2WjtgA5Jt8NdxEuYJ7718Ka8KVlmOCNfCrGfW8J+Ahq
LRXUVkRsDcL5nX0nh9VWwUDWrWkJVNPJcxT8RZ9EZQKuFLoVT4Atzmyaujz80hT4+O+CZ4ldm2DB
sAl8xU0kVVeXfzSF68yPAA9eHnc9G5zvvxhyNZ/CPLV3N7dh8mlRvtUgy34WQK2GaFqZhMTKlyoO
fT+13yeedsst69x2O84piZfUqyZCEGTV5vVE2SiuKE7rHO52HPSCaqfDsazv7lt6aAMvi3cWoK2u
I28PyeEm6LrIBUY1VUR4fvPj/hIm38EakgTWyOzBOVcXq6Sa31Vgb3HrH5rjD80U7BEntgo1ljTV
wts4XmUZprHOgKp6NCN3bCD1/CeqEuGF29vR73H8T9gtTJ0Q/8/793+Eq007nc/JHBo8o5BCTaCm
NItEJscHQs5ZdJNdMiOxE5GvvSm9emxfHc9DhTuH+WGUPDtK9haZugS9KS+6WmDJ03mO6w/zOVFP
3M97FqxfNou6c+vRtRrPcThTeWwNix5ZVxspyvvvvgZ1twohntvafz9POZWfIb/Do0xbcG94Oceg
tcb2JCdM01JSkVaTqIJFAhNu6AxdqlyOx3KEOyw4efT7R3aTKLEEoJmQj7Q35Bkn1x3jSu/pKa/T
a64aAsk2OnIyXJw0BScGMjy71CGjTCyIFB0B7YKmpSRTMwdC0AARA7qEYxQ0woluu+kUQ0KbQBNR
7Vor4DEBiDjJU/w8+NZQkW9lirDSz7316JpsV48cfzeiHTJBhs8anjpRM9QPvtdOTRivAKsHOnGW
14Y4MyBvHBnVdlj26kcYjhacNVFTjV6f/A6UGL+V9S9SY8nzFguppDK/+g9tnUOcAytXJPlzw1aW
qzDpXAdC8Zwo2qnKUxXV9LYShuc1kZs6Jbq04hZe8E/d+sqjS6VltZlGz2gGkcyWYvZqysxbUr2x
f0b62VcWx4xukPk0u/gjzn8KECrzKC1r3iacLEMiae8oubBNrflGgcXJbc6njVvtWuqpE7pAxE1l
9g9VsRthC+Qlf40wNO5+KOHlZUqL5zThdVvMQZXHidJQFQ2AA0o9aNuWuqr7v6Me8mS7k2WX7l5z
0zA4an9SuhgwrY1VCzBPmFKBEae+TrDwG+NHR161Ff1zA/L98rUbS9ncjz1X4kEH/23CWMt9BhA0
FfiSIVSM+rVXt+Ekv4IHZCELXnZqyPc2QX04OmLcVWDZIclf50AvM9EJO8EGdYaiL/azF7kQ617i
OksTjGpElqAPJYsriaewxGeZjXjQX8A1FMWl0MCbKX5ImzQaIQLkqgaAOTkoSE8bcRQmGd6fxkWE
j/1vJupQtIBJpDmNLEWjz5Cbq05qDVbdrzJYknEXLzCVZuJr5c7WynOS/VoJUpfISkZ/HyhZXfyS
IBUgVDXPE2JTP6B4piI3aqme2FAG6fzjv5BcH3Q8nxDljexTb5vETqssU6JeimJdtWEr4TzSUARd
ubJkpAmL7iWsfAm+i5qHOc3WDYRr6pyEyLNRTM/8daZVEykeJLCFj707ROj22KaXluWsWRPOY2JC
pHVLfhR8KXjRwylLwMg+6RVuWMeHq5y4md+kbSIFWC9zCNVlf9C8mN25jYjF4UMepXnb605TR2nl
ccMjhdTxrKVwZUtQsPmI53J2AHnrxNfjSNmJaSWQTxr1oca186ld/MSZusGSn9eEeHpT+K9MWpvE
KjvD20kHeoM7O8G/JrWjmCJXcZbO/c4XenIFNnEo50K3sBL1h7zBfdj9g1Jc2sIJLACRf+vGoOr1
TdKh8XHU2jOMSFCmDHlvVl9aD2qZS+PhJCCasbEA4foelxNgmAMfNXwZiWJJQL24qY/wxDyaughb
8WRTFtZzZ3kmU6DPKrPupj4osc5aX46hSduvHY8MTQIlJGXmddstKjHkt1DqNb3etWbMq3YzZrZv
MlnuX4LBxY+/0eZR8Jfym3+4gcnl2t3/6oLPOoHqIlPOQTbUs05XHElovBJNdygY5IskmUZhNPB5
TOOTkT3T0fLM7tBXT9dhs7jW3VMbk/XxaLQDZKrIJQB075whGwInolxJXob0jzc/P9wuO2nuPKws
hz8zdS5VhkTarFwqWGClYc96Dn62GlasDvwDYP/RulxlpyYyPo9m7vlM419bmvBjhsS58rsZmhSC
mGP9fFmUb09YHXPD0RikKHBVjaAZH7NB2lJFG9AL3i3nAKYahIYdaeVQ1ZL6MmhCMgBfAAejTuGe
8UHVTwvL956tZr888dFxEliKr28V9JLM46e1fzoGhh9CmwcozqV1fVIDBBcefCR5WCHNrANKASrX
TSmmtUFRzHeOCMeDvrtTjpwad3q5p4xBYyrP+uIn9gi4Gcn8L2Sxt9377DG80dEuyk6DZzd1Kmh5
Zo2tkf184fYZ1jmebfGWkC7vRbzRU6S2b2z6cQqZQF8cmzzZDSfMEuKgOoem66eRSESQCrFlgFt3
aiE3r8lzzkdpGzoXI5XiFpYT0MjD61tmSZso5WbkFyxzrndwzv9dupEYlNoy3PCgTQCDTntuo8u5
WUEwWUxeuiPYFgR7RdYg/lHuw1Ru/tU4uI4kpUWpuECuhQPQ/7Wh6Qa9LBydsq9oc8/Pigg4VaLz
EDKqabZakEiydkOFU9QEM26Mn4EKsio99d7taC3bIEdeXUf0fYnqEvVFkAUtpDme908hF412XHqt
3angNTQX7UjFkdTkRkwpw7X9wq9Nzxofb7+KUSctIAKPRUwTUrsz2rq44Yn+pmtJGt2yZr2m1xcp
NZhCCz4s7wrUuFDkBZvaMURLPbyJNk80Q92YCeJjBYynOk0q7TotwIRa+Ma1agw2hVrZsgPuz0Dt
MV2tGWa7Q8ulsyp94NE2GXaF+qk8KDGlOtAnHSmc2trR25rGDL8nnHCuAJtzbfeBB/RZ1eWWSY4e
y0L12e9bq3pzZ3S2sr0hZGWD/2lNjbrfb+kBK8HNpn4LRHuWDws2baY6x8AZxbksPXdjD1qzUOph
Zp/FCXHY+jr8FRUA114HLdPpt/shSgh+w3dNwdHJ6haYQ6Ng0MugxwA9yfTxfvsAkAM+3no7Y6No
iTPwg+FwKFSu5NDkotbZRUCd3WsPvMj53wWzf9vQE5KtwXTjxinKPyF6+OHIEe7RS0nbrvicAbRC
We5OqvPpQkx8eFcP+KfzK990m2RBh5Of6hK8d8IResBKqBeGc9nY1oDUAdia2ZwmVmi2KRI33CIy
A/KwZzxWgZEb4bSl2eDUxUFMbRbWNSZdzJGesu0gIS5+q8rO5gZfJNEIkHr0x09DP01hy0deb7n6
g1xAJcJc40KsP6NaIlZoZ+2LgJsgMXHXtEcE86swd/tF62/t4uW06B2njtTUdhX8IUC5rnHWYPQt
ekD3yikrKeLrlTJEpww2U3dmW6wgKaRsW8DY5J0706ejpc4DHQupc+MzfbGT5qGSs/rneEEYtm6i
oOW1SLKCMd1SlLPBGBq6LO0Mbi7jZlA0pBdEV1d16ajnDLVsFaHJo3PFljCRcB4+HscWWsSxu8RO
CwF+fGpx8yT1LaFZb82MR+XOAHJPzskihXsJ7kVGqyQ9kyEtctKm2Rx2Ea+KAyp9Aw2OT1aj5qot
V//4rq4q8PRQmZ/y0fzTNXROA6VBAmmDBUSijKEuiCktRycTwFpiSBafefikvKM8fL1wXC72gbJY
PUSKcwdNcmuw6qpcFk3O4QNsFdewsGTe6xFIoJAWk5pwSEgBCtG2jQXtBYH1Bth98Gq1K7G952ae
2bTCOoNdXNELAm/vIfhVpJ5Q5eMrn9Qjl3s4Rgm3d68QLIPhQ5+ZEC1dPusfjVq5U703VYjO7s7p
MKVfG9kTvsgnRNkGsFyOjVVtuWRJBJTLPd6WAC0m0D1f6eyIM9C4hUkPog0dUyHqRL/ifkzUfVB5
IMsbgHp+5OYaP/w8o4darG6obxZF8Aq30UwxnPpAu4FfNEDk3BCO/Yh7zob5wNbwAzpl1I7Pz7zw
oLfPFcJTj+VPAwXkj7GizEHgPGKmrK6d+sOj2mfrOYe/Swrt/yCBzQNngCWniVIRcHIjXg65mqtU
kTpz3BYXEJSjQb16XU0qppCiq09D3zt8Bwd6fzl9qBkVgfYAY3uGwFNM4ekFcuuKxSiSEVAbPHHY
cVVzoE7uVYbBL6JQMcUTaCS5uVzu1V+fcAmzfhzq6/1CR/GtLEAw2BBoE+jWpHi6vIkQWb3RvecX
Oelrkc4XhaI3Opb74yYvLLusvf2xvtDm3KWFpdkPqKs704F/2KCbAv3c9rPF2W34Qu2JawZymc6P
tQOd83s+2dxBdeWShsSX48S08l4ppjbwEY02aBDeJfmPfUwVJvWA4dE3G0GmsNxrAA5od+GeK1tY
GROBCgNsGtyfGiN5qTJfJ+jKZD8t4mXPNoh+op6fteYUJmuI/CMGFoLX+8pP7veV4oy/oOb8PNSJ
UzQrLVi+GIIxEFmQHl0nzqBPHpYJBJ6CJViMT8Fs0q0KhpJJA+MMFbiWK7iqF311viKITo/kfGH2
E5rLadO/jQERjpe6CMnyAlncMUcexfZU3whciW31OunbEQXe9PmvFhPA59XjPyxcy1omDavQmM0v
RM2m0P+GQcXclt+mcDMA/UnvN3W8M5/7KwTJ2ejtgVmUrUNJDviGzjTqjfRkHHNhx7k3qbj9lknE
/f//sf6M6nfFizMyzPaCnXEI8ZAUEJTefVVDUiETM91plR7ygvqNoQS18g5lDLRPzEldEUhco2Zq
xWZqsiRJl/RHM5CMnX0hr/7pb7a09NJn3agqdpqot07X6u9tE/htoMXlgoKsaYxlZVfsOwKQTw6W
/zC4YGilUFtO1KtywIbvVx01zcABccFBVBCoVVSGtxr6T5U9QQs84MCwQleA+a93Owr4hdLGU7OF
f2gkXubNW7X8NuDxLQCYyDNPBGFUrdufe3kbNrNzRWDKgudWGJtJXHgcg0uMeWYc+p3fMVxUH9Lj
gHCwMHMmJBNB9JPvZuwFHt8IKX2Yg8ju0d+JNLSsF+vc4/clvjHv41NGdhKzJOyhhe/WdUWxQVCR
3WZTdoE3Du9p7oibrL/1CUwYiyiYcW15/rE40bFhBkPBtMtb5ewvhI13sjhIZt9g/lloCGPPk4Yw
YC3fiVuYmBx0nM0jXtwU3o0iJ5/evVTZSrVwMPwZ3LLoUDnvMdhxICXW/LoRqqbud8C8hj3+mjXv
/v99VYIa/uO7KzW/YHcuQei3xlNYjxMtihD0vrr7BgxlwdevErBRCq84vHWaQWXWhtbA/r6G4kQT
TbOMXa/9SOz3XHd+bJNuSIpbAe1zirhJBWFzVhU9rEG+uuMGxSucRoEVW4vMWEAMYrtr6/BYh/Wi
8AHL2vwI/9DOFxpI2SOqe1ptdbCXAkoEDb7qciBiADvMAAdv5D4BW1CgHHHPb2MCumof0v4PFWsm
Qfue0Tz5vui0fV37+GRCtmFXZXvHFuPJCfk0l0/nyQLQoKuA7EfggDB/2G72Kpmjh9rTEbyyms+O
gFz8pgf7nUQv16TKROVa3D1txBxCLVGp5KS7i2rQA6mTrXIufovyvuLP3McnDjWgQ6bhVciRmQG8
/DuPzMNnnZ++VgMHTlZX0/SyeVJQDvKd0Pd8FEwNmic0tz6TYX8uqgHS/hTs/v5EUZovKudTHOl7
tIeWLzZDd1aQMcON58ldLTq1PX1rWnYwPOKo7rYhPkS/sM1J5KD8QVUwdhNvMs8z/OormlKfUN6w
UZCPinE7qd6oqYivZwInEn040WFlFb3nYgDgOmYyBRwvK8ymU/wVu+7todpHfEgHo6XJv/UuHYCB
49fi8O46rC40oXEzEGAtJuGMsk8ZE9HCYGSIIt0liZWNiSgIlQJQOoj8nsNJhMFDHRIS95CWIZZR
soYByr1M2+8ZhyvdJpgwvtgvqOIF/F5TbMuQaO5RVShA9aECpoBUxKvs+vJki9DtH5sGGZURRQyR
HZv6N66ynrY0DXJzKUjqySt1/ve6HA6yES+20w61ky+mZ7uYxOSFatAFV8uTQ1HjqhqFlhGjD+cD
3n52ncd7ZAIHqM4PJlJp36in51b2P1wQA9jmcg808t27pbYK+SeuNHC+e2/SQ+C0Hg1HhvA5kj+Z
18I02U2PE+AsYa6UQjlHT7YujoOl+NPO++McIs5lxDJyt4+bRxRlCoBG2+vTTlQZPeUUFYpA2ySR
gnXrM/SGVqnasiQZYGZVX5sa3egpqlXt+WwFd2ZdglR5s4ppila/ovEI/dkKgnT0caK9SAdvmaZd
XUYCjUcqP2iCRfF572qXWnu9ULbGEl7/ll8ku0DKs/1KkpipSGdLJs2txbA5h2YK9ubq554TobTp
DGmaC9E5CEzHVzfqiO41usgMFynUydYtcltw3g+/KhUJgrk5vhmOVJHCgsK7U7zIThK7Iyd+1LCG
n8kniJ6y0i6ys7chm9eYPVhA8C6aT4YJhVg1il85S0RvaEPhXyxI9E6BmGxRATuGnIRq82pkVo8F
MdOwBnksepk9acpFlGQ7Qx/GcaAqxyxJggKEZwUHAWJmVl+I81CAbs1u4Wqw2y2kTKiNAZ0Pxec3
hVdQqvmds6zNFqMjPUEe7FThF7y2Xwy09Z0icIDnIncd4XekoXE0WyqQz9YssW2NGE2lisI3+pcT
rsNgd+CQ+CwVAL/zgPfK/2myjpKc2oidxf4+MmKcVz92fj4TuGH6EFNG7cu6SKdTJ1dyZv2ZSD32
4uKcajcOJbFDdYw8Pv6s7Jl/G2jGE62BR9ACB8xt6WAY75HnrWzhT9ygJSKRCzvJW0boad433aju
j4MwMsZ7OSmOmu16xprhoRt58mxTfOWtb344sjRzPd1wbVqm6R8Umn+9Ztgme0SGVkVEa5HHhYEE
DvzkbsrkqSz8F9rSVrefyQfKm+A9Y3ua5wxFVC00wH3TpyZuu2FJmYaA/HWaVk5/ik3C71z5brs+
n+UZlWB+rS9I49LmgXIYHq/arnaLH7Nv0hHyavv3Tae7VIPsmUt3FjJe9ojTViJdxi2YI2I75ciq
NbkGJUZoYbW1LadWxXhDZG/Mf3HDhu1m+8papgRNc3AzGK8cNrE4WE3xM1c0iGTJL5zY+IHYTO9q
HcvenVBosT4hqgfb+oPTt2NLmo2BC2T0hl+1CQpmCjUBWFhJUOipXPUELW1Q8XCYLc8VZvSQIGgd
3F5ZgAjeZw+r6U1C6Rttu0gKi0cNyQ4Uoo9dQEgnlw7CXtr4vq8QqWyLEFdXlMkoDbqq/rjjT+R8
tNOugrdPWiife9FqkcfmUG+cvNsTjfC11noZt3qPJjofsMBftFzZBzq+LkL9tdsPsTeLJkx3tofE
4CEv8LXFVHMPZEqgk4CpjuT8JRsWw8+GBOyuzWi2dO1VzBXVmwVUrWer6jSO7nJQvVhM9LWuCXie
42nqS4Y5gsSiJpeaINfxPLLMWSZ/j3qWUG1rwUYCeVMlfFtuXPnWshbX7MpWWLgRVCznzfm+WsOd
ExYv7ITaAbxlyTiAh33gmYlf7zYrcMYi3vBga6KwC3wfolUGBGSvjsjQDWJT0BpjLwmgjlXsqUkj
mVjXvHZorBi1cami+OFFXCq1YWkT/uqW2wecMnj77EznNQlPfozWKdN9G9fE5/sPai6auLx4OIk+
kqNzC2c8G6qdo+L9RRxHxXqsEC+XejTZRkisLtRRQ1wCmhng81Eq8wEHejDMOzPmMm/l3GStQopg
qqaJm9jBUVkMYRE5JWVWEli+iFhpGMB/1FC7h5WLn3EI5HA/6ABNQ4T2rnRxqBsqdljZWcB/Qpga
Tv9Zp2ii1vmtO0qMxXCUa4E9YYfmtoOYktWuhJ/ACRpjZ6JJctjX9MuKWC5O7OffNqTVHi/LPf01
1Yxhn+IHwiLZ/KQ4IOB9/izmIkCPkJvpupysaCF/pZnF1srOcXObjlyQ0EiI9UQ0qeHxjq532Rs6
RKIc59XeNyJYkxp177gQIyUJ1jOiK0r5oZoIzY9zxnrBTD2vVIvfGxfM/DcsM4viUEguM8iDUWrY
jT7mOfu1f4oN+uYaOdh50s7ETcTKGsFZKoZTfkOgqcJ3VsAyskyEaZ90fTApDQW8LM91diA3ZnzJ
B+gc0lc8eYueyrpC8c2ic+aiofnlLVK2tYAu1fy8tXGY6C2otTVTOqLsHyIrCk9ueDtJP5KR/1qi
gHaSS8RPV6BagNQqi7XU7di+L2dYbAPAwekHt6E8gM63SYa2MSZLEHy6nDmS3l/GJEGSmgf1H31v
+8hRg2iq6hZ3Qpg2vq23KX767dIdukBEF9NeDIuVWj9jC2ve18SJactY0rCWHv17faBcKWTv/4wf
exXo5XMnHOhDnVhm1motO8yGUm4YcueeNXBDaQXfE6PIWSJvJjgtrssqFROYj4C2kL15PlKB9LmQ
5HRvdzTYpxtro77oTLCsI33KwQjtkMmHL+dKNsItPygF+3iGY4JuOdsLommiGD6Efl4w9m7GUG7c
eMyRjx6BLRzrUt4lhIi4WTsyQNXUm7B+Z2H9Lh11CU52jy79ezj6JvAglNPk+qB2EHChn5oAJ64M
sJ38GZjZ2CJVU225xtG+Y+SFx7o522+VvwNJMQGX5iUjFJOFTFsT82RdaIejmb4/QUQVSaA9TFtW
D9JY5bUet17+DEj015K6OlEsFrFpYjRUri6pICB+dLa/d83uAtVE/RfdeUHsYvhoouIOuG/xc0TH
bTkFpZLfsK2q/EUNKXFZh6KSNvftEGxeV8OqEaBjNxRi6NLsZFOsp8x2ewwSE1tPd79UUaoKYi43
hORA1hwWTCS0WakA0RYttYHj88JZeoEIbo2oGVnaJPsJU4KLdOJ+8PTXZfu59ROVTqUgzjopgKMc
aMuPnozQIux4pwH2j9TaC7Z+gxKZpcboeqDmvDG3u4kRcDS8w0NflwMDIfvQpSwcLSZ1ngw/vB7W
tIMeFWzK9EtJs6R1yV0dwIN297ksicea1hRx2Eb2Q83VeOuiC5P6BgC8viMmpSOsM9lgbyytt+mJ
fCT8Kz1p+Oev/+1GjYzdti0B6orQDB/jcWw47eiMeuiNagifrDLtCxPrTMeGfiUJwFxZl1F/UNQd
ZrFub9d+4PvlzlOnTSK5nVNaQS/GKV1TN1sxbz7OjPe/WvF4PfIPdY9w5h1AEtmjvUj2mF/Ms9AS
rpnSGuctA5uH2qlIJj0oz+N1qz6rc4WX8wUnijBFoicTPSYhl/f17IgnyDcXDWtqDui/j8429TL9
zuWO3xPHiDjRalNBORsLoqDUNOWDSWVOMNtPeZ4d9eLIXfQyISGvW+NiR8BSvnPyqbAowfUTo1A2
MqiZZCJmM0hKsPKt7wdEKSbKJWJPEVHFZSQJO//t7iuxvDmz8KAaFSquWGFCvmjRhAdmQbttYUqm
+vW1KAcaDTkl7fR6OU7O+xXDJ/1WkDeVc5SEJcAK/94hYoM3Q1CpoMz8R3aVwOFDogghViAXs+Qx
BTyc6y4GJ6VTs8kFRDmeqVYu+JGoRaKWohNLwOqFsFjgV9sgqUEtqEr7iCbMdCiGqlJCmjtFXW53
u+xfxtx1ahpbeSpA7duMyH6egyTYUIM2x/FEe41aoEvaAJOXAsRK9M7+g/XGQKeHdDAKCSE4RISF
CqExWeOdvmEMU+JQJmFdCSzO32SI6ZbXW5tQ5z+GrG6kF1QBeLWxAjAV5IWJzYEGgB1etbILLcnF
na6AkC67XAV+U0b5b58aBtBCBCN5i89WOwIEhDEiY9bAXTnb3pkwyvPA0210TTGd5Y3K002dZo7m
XYPRcs6+KouPiC93N38amJ0PFTlFBjKGun7/pa5FbqA7RWycTJLw4jbtrKOHUzDspKKfUtQ1ew+C
76OqTyKUdcsBm+5XViLxfIGKR0nO52GCptrBJvPsv48oU1uKPgDOAyOxMdiv0Zq8WTIh8q/s8d42
cI8uTILKzDeAUzLxvrpUrk+RNiIbOR9N411pFtN3c3fcWSt57wqdY26CFuqnlg5Xtz0KDsi5bfFr
BFExH5poNb/OxWPkC3ZYQ1H36NLzOBcFVdbZ698H6Ft6WdKRZjWAbrL1sT3AdSsfR/hIp8gZKJIi
Be/oYSbpLrn+IrDSw/SbC1f+0p4R0vKM8KYGqzPUBL9tZwpsnMrkpPGaZr/a1/sGRFCiggqhOXBV
v0f3opPstG8pU1UIQAYJV+XkkjOPmRxVUBhqtf69gCiWi+n7kr2x8+2VWFUgA42sAn0vY6lQFVzL
FtyoGKyQMpJYha0+bOkDPRCruXhSdYW8RTBamV3b2bjZf4+AgiX2kmLcMU49QgTsPkozvj4Ow4jG
DdD6Uh7Zw9o1agppOM/QMKeikM7BA9+YV5MhQuozAFyuxNMzgfZ7bb9U9EJSNwtvqQ80zd/fMjn0
EJanRCBkeXcVUzZqP8udtRPW9y857x7VWvnmVG3ew5p96mvGQObWsa+Z2GNk1VoOTLiKEW2JS9cU
AKRQPDqPtjbhqnoGwGgYrq9x3eOt1bbOvIrG+ziB/ltsHHGw4vUx15xFADGOE0h3C/sxnXhjx0nd
4zwngm8rUjqTv0WLK+oedI4G2gvsVrPNCk4N2lLWWTnPiiXGxqs3hvYhRLfpJ1hu4fSP+zgHRbOW
8H610im40EWNJmRxZzQTYjKjHNZfBVRkEoeVJjaIPwcryq39nTng4itTfwLRxtDXHaJ0Bubmfrq/
zZgyEUdppIBMLv952ZV/gIjyFisj21s/Cv8Ih5+dZjwTkxy5GgFWo7djmy6Tt3ebNfS4SYpUDh91
KdJ8LoNPBFAomsviONNXrbiV3DdNkuMjbBQ7yTIZgjPKRpnVjb4U/sr/vjM8bnC1EGPdK85n2HnG
u/0tKbVc4oc1gQmL2x4Kv8RFMbzdQXFwv50riPM31RCAcXN0gBYl0hMo5JzHxOvJkVU/8SmB30fE
2/ct6WfqRJx/R1LGWtMRvh5n2ck1IacOC6kK/IUXl89Sd3yd0wVr5DI5c4iox609rFsvmr0FeERC
eQ8atbiiyFAgrQErCpNGk7JZqN+aVNtKK25ksNcLfhdD4jgIqugfT9cSVOsyS8K4zotwDVtZUa6K
K7DAAQME1YS5baMkFHIibAtEyooAb8BvXLYyOQzUmw3uxYQGIuvynpp2n7OeMVq6wUOFTLCQQnyR
eXm1aAx1a3G1Psh7IjDjtW53uKop9/BgWkMjF8IY5hWpvtzz99DVfQfaSJSb9xRJUNCy38q/u2ew
nN/f+26vNb6s7TyUhWskGQAu8Mp0H0SSJ5gbVMeNUCkSHiaUaXcryYm2vMif/+L+ntULhUhY1NKN
IrQVjN5ONIALc0+2zfJ0S9dR9x03x8dkt9b3K/fjhaeyCla26Rw5BNeiQSpHdBg7D9oc3iGn8bUG
i43xlLQ9lgRAp4HvT1DuKbAgWDHccqVL5fkzKFwETvIXjE4EU2/R5i4lTNRf8z5tSQVBYONIpYcz
LTciNLXG2itrAX0Gw4Bc/OuGNgkWEvSmljkFz4lfQ3QQ6Cs/nj95DP7AWsNKH4KU4vbHu93Bn6tL
IDVwZ92uEMYfxoJQ0/Ku2zBsKYUcSTf7CF5EpmmM4Rwgk759tjnYgUBFaf1CRSCYLBDnnLoH/P68
pMmapXRBBvlpvRH+WpR0lzZzatp7iFl9Q9iWFJf526GQXvTW2ZFdqsvpSyLn8yH93HOPDAh5Wqz+
M79TpEik/P+gtlnS9czUvIH+GZ+pblZSd+T7p4Ump8yA0A7rbQvRoOJdgCdqDUKKqEGxVNfLQT69
aOxq/jBR5DBESk/hD10+E4WheeQQsEPXe4HqjCfY5goPsSNOHDwV/o1DvDUVWCQr8AdLVX3kfrfS
cqKK7jww74spR5JELj93qOh8t9mvsbYOS3i45ORiC9atLrxDq4iEqsXYCLbb8iKJKVpl67+EkCmc
cQzF0ktwfKCiJM9hUNjlR8NHkQAbsGmLv9qa3d50aWsLQImYRfX/7et3IhRg92GikYt2FHflUFFz
55sRpPqE9wftytHuayKA9x+gj+qYjSZehV5UvtxLFkDzxOnbT4G+81JF1SKlHvImlyEeDk8GRobO
Pu3vzn9yiRsrhC+DZ3mFasW3G1L6Dp9cfnqB0uMCZPyBGaK7HhPbd84+6vQAPZMNGm7tlWTHbFUs
Prx95yfuN1MBTXq9wTKquPLzRtHseSrstSbfQsFTZrMiDhuqdTrZIXCSS9IlWABaxHRDHWzRkIMD
yZpsFaz42MMQDQ+t//xRSSlE/lg3VAih2UnhUrdmXKainlDv7ZDSWwj/tMXv1L8CvhnzXmDzPAK2
dmNpVqbTXc4XU6NU7WFvxANfkIZUj/rFdB72Ih1yfESfF4W5Q5ZFLluJllCjo6Qv6ZWnloXXH0yE
qBxIKLYdm1BxxF812wlwqVNDMvWsysr2aAftegALMt4d/mPYTlaph+X1m0WuYwKfhpDrsZXQFgLR
x5JK8sm1ohqahHbyyzspnnTnLNrCmld0AypCbD3zax6AGJAxrLmeQ8QJwyQh4JIDuFnWZPcYcBvA
e3OPyHmUo3jWgeiZFxLndJtfmofhaBXRzTMlH3Mmr7hvHtgg4cMvvYLlBR5LBiJVHvNeznbD9Q7D
o09FOkS1sQNaQcuy1ADKAK+kxGJ9fDJez/KJ9oejzUhaZEIDzsoMInaPL3A7OyhZYP1jN5SLVHkR
TDqH3FXzXeXSiUE7mbhEf6RYIrEpcGy82VexgrP4mEWKWytQrjuMIVLX2JyjKjp1S02+32WLfiSQ
SvOlIE+2UpznvaVJBPfhwKuVXmJB7A4fczQmYgSx40wG4+f6QTnBL5/Ld4A1u0D5o/zf141Tn6FE
Nzd7dbgZ7sX28pBQYNEIn3S3YA8UCKMeZQKbDCYAsu831C7YabiVfrSHf8HYVSkMglXWXxtMuyPO
FvIikzn75Ue0t7cb/CxEzhtXJhrTF19PWCXBqaSCDV2auUK1Os5rys1BRW4rlzAk2B8d39x0A94P
Flljea5T8v0GbtjMCK+cJldDfAn4kcpDwxvLoragRAN5f53ofm+/EgAnuGuz56h6Ox9I6LONbFsU
Iuxm3lpHUH+KRao4D+ORS1kWJe4bfTduiVazjgdeiSfkKM8PyTPkxzeGGKZp+cCQp0Tnsjw7XmaL
/vy3cxnIZrKa9eM6Vohriex10vkzK47NgUuH/6pVojquSzSHRfo28LKFIzTrChxDHN8q4vCSpBc6
NN/LrIyVUAKzvo+F1uYEpa0pBBPPa/HAJ6TA7+6n1NbE/W/0bFy+KywUuuPFLJZAnI8MpBZ+LeL/
4qV+nc9oKBPxhOWwUBnolGQqdhm19LUH4xjjNgXERHXnVGXMVPh+04Sq+Zd6ddtNBf8gghU4sOwf
Yx5nyCIMXby9U74EPpQVgxsKjKp1UeagfqgIU3+MXHQSWSG93qdQIP7LrTW9bjDCBmDfhCzD0yJk
BQd+kz1VCmaw+mOPqdwlIZ3QDHkLjSwYRLrQrKOpkYcEOhgMX8tQAS3BIxPTfW8T25mFdni329K2
3hDn/o5jB5kT+WyDPn5/Knf/a9KDtzkxWmVq1IPwUDioMRy8OflCkeHJMaPRrg0jioUUMWozJWqy
tbpx3kaQu7Oifodv1NzRYKJpgH7wOQ3P2C/GHnDdSzoqA0XuBBclR5+22f7v1EY8SRBUgzqwNW8n
4cAQy+Q/XBJtO3YiM+FARYQRHy1/0bDkMDHNTRhYRrEV5l90VjsVl8AZib20/7vBqcI6FkY8YVWm
v0mMYZSYa3wvDTXmelX/j1sal5zzSCn6naUMZ/p3XRN5QHRbFuIe/mXVP9tpL9K+XviudO+gWDDV
Gqbw9y09xABTOrQCL1DXiRWc/VvcOdTn3rWtOYKoG25BjVOt58uy2AKJnkd5hFgFIahceO5OrjEi
9eMrAzXBVt6I4uQHXZtDcTacDtnwEcZXAHClQdBBkVk9M3CW9o3qxzaOM0um9fuvvlqHgV234e4L
xu92yji0d5R8bXZcyR7oCSTBvP+ocnkgi0wgyOaswtQWTnH3gXI5eH0Rvlz0lkBlqTij19gx4bJA
lrrOBckOP2fuEn1PD/MUPh+S36x7LCYxUegK9qJd3auKgddGz5ero4tEIAxV7PL3xcXMgkDpCpzC
lCjqjLAzEFvvJ9Ntzv+2P5XADvjz7INddojafGwsMjlNSkDaGackbtDy9KMGniBD9jQJtcOU0KpM
ZLjpwUEAOD5hyHTF4dqUf13imVC2WU1e3X1P4fmSB0dW9rxyUoEwSAtnj7cyvEQKlePy+qM0gwQd
Dsmm5/DOtrtlQeR7siXXJRZdA8OAfjGT/4AAL6PDP0lXHx0r2GqT+bl1RFlFZgQVXrzneeOiK3BP
8tacEv9kk5dsMPg3ohLVrRB6bT8ulHxwtDaSsmAal+H6ZybxJqajHip+scPhOE9YHdA5bhbjfDRr
z6nmVh1/+iwEMELTj1obspVVpmhmhvcWnK9QK2spn7LAJrJoryc+zOBbH6MQ8/4vHstB1O7Pfp0v
nFiX46ddSxd28kfEx8iTHslM+y7y9CGxYM11TxbKKJUIvarPvtvcLn24hSCDCYEbtK+3d28bcYpo
h8TNc3v6ewXVDvpP/n5IpAaLx26EFNsFKwxbP3w9aEwTbER96/j+90OXzO1vhKS6ixzVFtq+8DC4
/guRp+gyWzqIPPVtdBY4wWyh5VPUfIOGZ5GAkz4WqwMwDvzdII6tgkm20h5DsueetuYOvQSPXMvf
92FB2X44TNGGPkP9mom5l8zXIc7bbccRqOL04jGa7J9jld7obYdmn4RtfDU/arVujLOl6O4yp41G
g583C0MV0/aZPDhzGqTRXEmQvq5NMEahMSiqO+K4TrSqlqE8L0M18O2lQpeeG8yYIuIUG1zvjRNs
S0k6QR9zN6yHqManzi5V/wS40HjYQ6lY0HzVUFovO8UZypj3UsyZeiKJy9gexHFvlH4ssWTr7Z2x
GFsxmJqwl4pD6GZwU4TSrwFbysX8E8hcD0pyfJYGxkQIA7tmYFrxAaoXIxXLl5nqw9e136Y6YuNs
aJj89rj1KFpMg7gspBaCN7fPAZCTosDB8K8pxYLTZsiRBmVFm0AyrEEUwQGDlhoSjK4BmtQ7bRqt
IZsLJlC8ZaGnMufKyvc//MTYdvIJvqyBih7kfQXM28zB6ag/o6AnX3F1VGXD9TG2/IkY069bPci8
/rfdmHkMJ7dZOu9gDzBvc6gv+NqF35rTAfnDF6Se8QBUP7fG7AZCDULyx8TXCWw1XpglTrD36w7T
X9kpAkRKpIDLQWPivOXqehQ+VQRb/sO2M7ysFcq0m5o1ai9se8jKlQ2e6SY36YmlnInCCLN9HdNe
59RNxHJksoeWD2in8oUd9zS42uO1h6an5wW5n1ls1k66V7A46vM05zaZkVdt3ryI4KqLJQdSb4ir
uoSlKixo8jDn5FknxbfPIFAlwlYTCRmXXXkgq9N0SHkrzZQeRqd/7hDKKm3aKAo2CxkVo+ajve1A
/0iQBKhNeKOQONpU66l8S/dgzatpYizbulrikhG64wBmn2A2mdnxhiBRdOJSgoqcIqxzVUKfGs5T
HmxYnlO3BTSgUCLwJSba7eua4z7fdpW3IfuwdhmuKNf+Oijd1xNzA+TC/MiWyXu6kGZ+QSwNz1hP
hUVLeaYfUtJN4+7OFBeeCxuX5VYt//WsqGhYKzodbEaJXw2lRa6ZTrUDhHCd11+CFnzbSXdTJaat
J+eIN3t/RpEpRQPMqibmY2RCiU5Kj9D3HtzxvP2zhbfu9l5A2tK3V4c08J1QzuIkgK0OamZnnX5B
caOZTg7vP/fo1AzpSKScqSPu0qNGSehVI3sjZa3cO/eV/IXEEI2ArPv7ktAQfueObGgExOi+uC93
RY8yQG7T8y6jzX+j2rKYiFJGIY82Dxa7PvL1SjxzlOfVc4BH/6kMlbWsWEM1CxihxkdmfcdrbMJP
n11CuyT/+NwEw5MaHFfxFr4s9naj785UQPJv6Mw5+GQYHneE163T5jJBtRxwb/zVdSn80pSXDv0F
Jsp5omo+vsQW22Ucd+DCZHAWPLAG2tPHM9VEc6DdmZ5Bu8eTV1CZG7ncUSsY21HZhv02LqnWSQUS
qrCpFhdEpeC9JZb4qhv2YeLOgLxjPrqTgcaE4h5qNMGkrmhcRKulUzcXQWWnkWzNjtqiorFofPto
YSlkJ1SjvYShuwOwOoEwtYzDNMZHEzy+ORxugK9bLlHKM1Vv6xImpjIsg7Vkiu+xps/43KaIDPWg
NehwCj3xSqf6rzUNkPeykB0ewaHD68uEZeOlFI/MZka85WRfj7VkNUF7CJHQjnW8qCf5Qr3nfwJA
AWPxnI+ozu4GvNj4cPPysqcZCqVmUDBPxnh1w9Gj7UvZboAclcvPrSyMRY1CRj3swX8NDmruDfcv
x6nNeqiMYXwD4PfX6EGVPeqY/WkCKMcETWRiIXcOGLwidpUxibhoGr5OPkEaiTJP3Bp+cyrAvAYg
DT/jW0s6mXZ/7YsrGBDyvHqGTaWrN8f12qJztMJ5ySeGmHmpoe6FRayUQ8OSiyvJ5vysXh/9BQ7f
Z6+hsLtUekCd6Ajrq4D0Z5ydcpqYA6rg6KASPkiXIVBZJNqz3UVw6pj43lIb+qt4g4tREc4cRPB4
V/8/VvYrbykbgzwae3WPDOd2Eoh0YbizErkiAXiXmabEO44GG0IZgViGgKGJD53gcYvv4sCDTHbl
BolDNeQ0bnRkHlM3UNkh3HP92R3hRLC0MF1i2dRQgsii1B5huOLDFMsLPM7BLvZJuKtE/ely5m5Q
OjVNtUUva8oNqHlPqu8uhk8BYqgbrxTRUG4gBMOIQ3G95nesonFPgxUuDxwCX3kzuf+3V2klsG9X
qWyymxkaSQTEQXJPlvl/5cXuyQXh2ekHNx4g1IPKsiBSSxbkIBdgcVte41x3uV4+dvs+rLLYzBJd
BFTI8X7CVTE2+fS9cZOibGTVWXqCEmuaLJIbyM4+HDO83U0EPQOQBgYRDvdtQeSSb7nDa7fw/7Nw
q/LjZzQ+KzKoInJyaERt/+LlvpOvhz5yyHn+Ce1T/d959ZEfQ4SEdRM0SfKuLVzyhAubBnjlni8L
nw4cDI/IKZ8URwCKOtRmO0oU6dRfNM8cEvgk/fqfHKRH+KZbhEKzt5Avrc4c/bToRF0Ki8RJPTYR
7iXN/lT3SCKZ1h1MxJjnMV3SDps/ayJKSPwHQwOSzYukLupwEgHaTSA1/yJGastvFD4gEEckVlMD
Ii37lbAinHuXbfz0J+PQN/tXGmLRAoAkuwu6P1DDU+LTsRJ0sslK/1fXdY2HZIZWusQArRjmgWff
22B2rqkVx/KtVVjfRsmG5kUvCa2XQRQs1KadU+J7HrFRYL+6oaogkF5IrJxK6q+wzbQ2FUbXgcju
oW9Gz4wtc3N6u0oQi3ZiMbm8ADVcPtPcFaTfT9PuDCN9lRDOuAdgGLf/GZOmkv5b3Bs9bK9RRkwG
03D/9P84UGUiN/ADjRdVwKEQ5f+OaNr8N6eUPXiU4e7j52YrUr3NmsQUhnbDn3u6FT7DTZR2fXAe
LIaTUw4rCrVCFeWDf0UePhCVFjdeMinWVaQWws00Fg3zc/aLr3hjKJrECyQDzixAe10KNCv41adi
ErUQedklMqIsAUg/3yOZosgyOh9effOG0hslgw9LNbzqBvYdQiKvgKY2WpKYKkuWAvq3xTBn3j3I
EWRlmKKiLg7mE3a/H6Psr9Usu/i5rSgbciRJnUvXZeYqlBqBa5fUAdf/xWNIay2lAHGi2dAaXI8O
5TQJrvdQ1/bfUqmb14tlXDsjqzt0FmiRD6zfoAb1ra+CjX2QwG3WZpwvhK4++36YhaJqrOlrj+YA
+ExqxMK/6lDVekqm6NDDdrdc42dxKCYeCmmS9LmuQLC3UlmF1zv46OjqoQZew3LwNuYSEksal34J
Cu2GHAF791R+SCnd8wCU3rUqIdDmuy6CNOx0pK9mrw+IZX+cACsfjjfSA9mZ4A3OZuIZZ+aSO5ty
9YVIrN2+t7NKyJ2pB/6msVTTke6ZxZgjVlxnIQEfRXN317gOsYvs3CiGOKTi+Awu7ywYBS4ryxMs
BrPCdf2mwznUejUXKTo/jMIk0izHdlyP3VUEBoIKZTDZHfNTRYxqXvB8cv8fpSNsQpqTxrdM+/Ul
B8q57rQGfAaIxiYgHZmUnfLHN3h1bRxr6k6uD9taPot/JlsnCOJjiHHfozB4Hk/ffjKT5atL89z2
cpH4DKcmsnlcFbs9y1N3H0oSfe7jMKMoON5Xjmm+vgPM1FTm1ZC50UDwMZoekZRW9aIv50brqmRp
fSh510Sk3r19u/yhIUADjFhVFzoBmRFJLUrlgcMSWajPirqGNM4n4Wm2miYneR6V/jr2dZJa08xT
Rsg5AFnnfoyoL4P+KYQ0G5SsVfisCY1O/iC4ijVnujOjwpsyZ8nbUJbLCW6bZUc5w+6mhTeioY9x
UC5LRJwcrruBO40SCHynNKwNt1wqQoYWlIoH29Uy7wbP9IMGZPzo1oJNccrVrFYoN09dKyKHMTyx
WC1+0/yTpdg0CksVo7Lo8wXzgYnQtfNKW0ZbEPB4TtBXGzyHP1pUMvN4BaRHYqvQQ/YmQYrc2B3D
qrMA1RBldgwy2qqYOFhrD/YlyLEUqtBZVnXq+fTdsSIFoYiZ+L3PwcMAGbhfZzni2xJGNPU8Qe/r
IZx42KI7GOqlHomVrXK9sr13dVTMUD+1fPe5tZJjUdpfbvDcd0jtWNXjeDAOSFRpZyc273Dn0VHy
RucbPIsrrxeaM9ra8S95FZ/9GkZqg5zTJuHdEHdaTdCn7HKktwrSQxLmv1kWtiT6/3iMIwJfS0l0
iYtqMrvF7yeN6nRs6+h91WLVKn4kghOwbJZ9reGaaSZGzepxv++DIlud8FPRGWC89DKlhicjK9Eu
Coz6meYKK+u1Eql/ESocpqLB2Kb74+EIZc1p0myb7m9aoIp7FTu5PYsBThKJHwlD3DmNr2e6saV8
ik2ojpyUd0YPpImrStzueL9GOT3Fk1F2xOCQbmDR2ixQq4k4rjdgzXeljQE63q2DTAUVnXeYEIcB
8kX6ukJBbsBRM+CSVTBmBiv8LhZfYSEWbhrBcUSxfNUnbcGNnWiuN5zdkTVod8bpjJIUCRXm9Kr6
3uygTbdM+ENHhRlPmsAS0NTfKOBGh1/LRgW+CSrg+QWO1COaedi6eJONUFiKjqhlnlwgXloedHs2
FEF+qwNgWmZ0ZIGQCQpKZvcJr8h0SORD2gKTLf7fUhGrIPogv/WC+ha6HOni7/EVQ2Z2AGg8NWgV
zcHe09SY8YywrbMKO4JQLY7euY6fWLs4XMVEXnFe+78s4V1dqDuJLGP3QJMBufPSlTj0F/KwrWor
kZWbLgtwaYXJBFzDAWpzj8GzkSVK9INvWfcA8t061yetk789PJhS45D8xg8k8OSS+pYjz0zPODN4
0+kgHVhLeT3uN/FPs6Rx8AOZs6C9zK8y+bdLYurGz0fGWz2Y/dFX0RcSXlKxynOOucv4+55xH/7Z
NOliIIMcjdPfTKr+jCwBq74FC3zNOm9AZ0oW1n7grUoAnKhOSTjBINBMIRfCFAfq/CJY7OREZONM
/a8wR9TF4x9WubdM2X0j5fkWt6h6JXfqoj9K9MqLClqGyShc/WssDZ/lhF/Mn+1B+NzPX11qEe7u
fnU/JHZ7pu4lxFwUZy5sgqFS7rv9E8BBYoBQErk5vPbH6tGxR4pyoGco/OLqiq0y+PmqvTnY++0+
VkeUvKYnVDpNQ5MY3/foeUQxycJr16Wnb3rTqkPHSuKUZp6WGh03IzzejCkvOd+eWl0e7gjnw3Ar
jcr+TywSl8Rxh9fdQLJSUIWaB0gE3UvOQ+xOMOzUEu5Ft9zxHBeVWOHiqnQR1eevSlOGebhb0r8B
tI7/XkzwjVEppE2YaKkYA0SQ8qcJTNY4HaW/AX0pysGBvsiJJCG/iMuh1tC3htPVgHvXZh1POxVt
KlmmwdStTe0RayiVPbArTO3tYlk0/YIg+lIRRKVP6zXN/xTRjTy5ZZsswhUwskBBTUZnsuNMGlJc
6vm4YUxNqTVClljMFT1C7huPvIyf2BBcxW8Hofe2YImK3tCNsD9sALWjDlqUkkBcYjhlzq45x4EK
N8cClPfMdVv8FIPLL5Wh0yQCkFs/fx+arK0jpzS8nM7XZL+GcT0LrJ4u7pi3FIiGjYSVadzV2UnT
WUjbcKcPTMBhLxJd4Sr5XH8BXliEJQ5SEZFMBPpoS3AAsQuWUK6o5Nx866eQJ6KEIjCfRsjxcemP
mjrmqLfKJKxBCm0kNIpWe+GU1IZP428TvlR8PwE5qLtNoltEjlPVS1DPNVJBPDV41nC4U4O5R6d4
UCv6cU9tlNRpGFwsdhrRqr576LUHwQcEmHC8M8fFyhVrJm6Ba1I6bMGkYaOIkHwU2lCn9IuFUs8y
Xgvm/25mAEwz+xILgycobbHj2mWG3I367ufidKdAUPXI5r8wsrq/5JiskQTlfbhmqkhJPvIcZ9Ch
uQMbMK2tK5O50Q5Q1YvbYCRTj2BPoq8Ldil5r91zZuJCINWG0kwTR99AU300lX14InOMNahqJaNY
BsdtjijC35/ZahuMtDtLuVGyVEsdfJqXxcP51XbmXRUws90ZZ94RRSulzA69ACLMNiG44k5jUODj
QaBFdtYvHCTzgL579uctUIW2BYcQcz/bteivjopE8mmGx4UAIl6ovHKD6ZRztoWSXfQVjHnkrVLB
rpIkyJCYMPT73nI94TQoQRgPw2rwqxIBNBS9gebJqsJuIXR3WKXnbhgIuYRZpE7whJLkx+IzP7Y4
cp9UvTk1zGW4Uk+teneEVlRwNj4NWssDcEaAEK+6Pf9RDC+ewH3aN3Jd8OnQwcP/Nk1fyI07wb1j
IG7gLblvxQKLBlHtDef98McqLUu3fGdOusf08l7usRnVdwkFbXg2BUhhPpyEZi1TOFOSAjUGNafa
QRqLDt/+WMQ6kTAIB57H0ohbTO0pwzkSt+Jj6uO1BT1OxLRwftfN1VzzPir9V1KQkHXEFj9iNnqJ
Ev+1Hj/N25SJ+ZgNNZ9XTVfxQYBGL3BGKWdQmmALKSITUGce4mIN8OzMCv8zawHetSs2okNeju2x
kkyak1rv18ZdhPbURf13gt0Nm2WgPXhQztMetsR/fAirBs2PwM3WMSjAgYQVvYqo/kDgjBqeGFr/
SMVU0x7RF2g2KRUQr8mQ1TND0DyeqB++y0oDuhgeFjCzZ7Lxog5eMYl1XE8e8Jh2VtZObBS4kWO5
QXc9jRKESzt4BTutbh19VMWhp/b1VmEf2C58Kbzcm29FRIot7raMqv087hNWDY/eg3hOhdA6WE1y
GX/l8Yma6H76BoGmuDtOwb7HSZDprySm1Y4Y9D8XkErtD6yzM2jmSjXIfOhCuXx7ndET6Ykvny8V
o40J53x85nmhjWC5AmBaTenIgnd7uXiEvRKZtyJ3pBQ/MJ+VKkaSLBqR+quQoExqeeavClDYb9j9
UOEg6zSl1xL9GbNG0s1mUOJ1XKa6qLxFwJg4OERpU3Ryx/HIucfGsuZhBB8j11AwCYkJNUXZXJp+
LxzA/Ru4u9ly1gOcfJ26JKJZG0+cBhhPKIvK28AqU0sKwlxGY4UsIer0r7zleqe5O3hI7bppysXW
NPxUJD5EZ2EfDxEQGbYdeMNelRdoMjc391gMmvMcsO7YeIx86nKTfVJQ6E/2pDW0dYSjamYQ+c/y
337/yafL5H9cc2Jedy7ucAdbJP894mIsr5lERBfHE4SAewHPu7M52DjgCd1FGZgVramy55yPhj+q
me8aKaFqitNugtrFGmsIj1Ro+3BGoWT/SWXiMC0jdoUkih7Hgr3fSbeEHoNUBQe3myTqj3MXJOrr
KXpczx6by1G/gAWpyh1cRtHxwv5B7ZbCxeuDBv/qNqzFc6q7pKQ02m8JsrKM/sCmwklxIVNGjmPZ
/2wB+kWskvbAgCuyvBD26zXqgoj1dPe42xlrSh01JDQri5rQui+ie3IYY5h/LB7rwMZGNAhrzlxn
v1vFIdTU4liSTeFTZ7IIbmlIkjBRHrzuMcDw5j88HNA1RxLM+2mkqsxMGr9+tEhcbCKUgbTwdOYV
tKUgnt1kF/tZzAcO0fcO/Iq5hjvphJEC0KCPCmopD5HA69YObbxIcyd1m2kOrQipSw5hIM16Pxgl
TcVmtg5UWaQTARudF3SlM8cif+ttberVOi+uv7UB/hSfVRP18b/8VvdF+UKmUHKPx8w4kvslXs+S
jB9ihfuFPoCsF1IJhVN0wxRCt5IT15BChhdd2xNAjqC+5yZTMH+wwgjSwJSGdYmKSXWD9+Gnz273
tjTHcGY7RelkZj4jAYJlKajqzMa+DLjRePR68MGTh7vuVmMYXTfMeSur9J3dHuSQwxB/kpG1ORfM
iperCGePvbydVhSMk4ShBeFpgGjHYZnj1imfT96EZekLF2CCp1IPF1VaRYvgUEF+GP9T9vkzlNKS
cAem+PDmcsHLfF3pISCvMKtBwUoCHJk+Yl4+gBlltfzQbA2a+1k9mRQXlUmektsvE6venYiNKlDR
TaDXVT2lMhRmCcpeN0NdkFHUJoDrU3ZW02hoJIgZZN17UEjv6fflxOD/6MFH1HJQNeu6B5fMVdIY
U6lC7OGdQgYwbAncB8q2i0io92KI6pjlUY/jLeCdt4PdadMk/q9Z+LlqYAGrTI7I7NtU4JMfL942
Qxx6F+59xt8sWGUIRwTVAP85YEZ/GdsEgogiDoq7FWlp0fXoJZGBgCYGkDN3eSMpE3cegSO8Iwj5
AkM66vWEA8EAo26ZyGpet9ZLwWWgVSGkNk6l2Z1fS7FRbg3COYmyj9h0FU3XbdqJMX0F9zlHs9ve
CtASTzdi+uiJ5EW2vI+2lBZL4N2UjOVi1Lgw/XQ6j+co/1lYyVpOp6bbwT76DNyquvc2jzsmfcGv
u+GYhZIPhR9d1lwU+qV3JXMlV9R/0SM5+W2sR6tMe/I+SdcyMJV4dSaRAkg/dqi6hVNrtxOp9gP1
Zx7c+19W449J8Tw3CNF3SQM2GDdVee8IBxpX0G54BmocVKofIAE9c4ajSUzi+v0qBVz95EsyC3d1
i3Jy9WPRxHrwVvD0GJvfujUbBS5NEqDbW8tlAdRByS3liuB0GjNC1VspooaPWIFbG6pQTI9MjUzE
1gruIQOlJV8GXZ8zB/uzj0SM66cGYtBT0108ueAYqgOsmYZlIHc7+EwucliBjoIf4KNSQYIpkAnJ
YgzjoaNAjNdjzkj3QOEv0TkCuRRNIGObbgBS+DAzMAt69+jGGvp6exNHhm4M3xQK2r1qvCXbe9kg
kRg9A1fkzn7gPbJF3s42j35ihqxi5lEMhvyDR8GTpwB2MdIlNhHpjPMts/QpDwF4KyOdD5ato3Gp
tOj2UBwEM6yBbcPkPa/Ouz01z4imnk4wT8ZyCrwopCSgkdcEItWdmehe3eh/30IfjWjUPGMFVzGl
DFF4yQ3aUpvA//B72XMtgcvdQYL4GA33YfFCmpCyIzOjt/wToGNrfQsYRQVdMjde9W+3yI7sgyal
ZAUSIzVPrVhcr9xOVZJ8qDfdtKfkoxaVIOoWRpCjMb2Ha9ZiA9GpUYsayfFsQ9E4EZ++FM5GSLle
ZNZx3dGx++UPIiI+tZoDr+5fP/94InFpXTg2UE1H1c1Bf8JtaypzueB/JvwT561rKTGFFmkZr5UD
rjR6sMREV2qfLH8VaQ3MFyVCpTw/R7ySY/kkYz24SpQbt2k3HzMMoT37VBAOKnZ2oj69Z8GOy46w
hMyfK7LSwTbAm6ESzeq4AG9CYV2ci10J3tzSXPM0M+XSM49Sb11HBugLcRu0hUvbm9NvJlqc/5Y+
2Hy6wnv92wCr7cs9JXA3qi0iJFUz6BCh9t1n9AAiXRKjglVZyDGBv/KhZJ5yb62kv1z2nZkCCTMl
rrPag5pIBLP/RfYCAjqZramXt81wHFpRpJYwsIUdH5eyIM/yXLvkwwymTYe0tORduih/d8S2div3
usvX9Dz6pyQnBpKP/+ilvz7T9eLd0FiOzzddMp3bnkp6rdmvBH2uEwyF+mIFycXOqCVVeCm71+iv
hu+dNuNUsrhpErXciIfAkgQE+6Z3cuW8t9s83+J4Y5pCU1uRdONtlOuO7rMeLo837wPl5E3rbLY9
0pOlQoBsmFO8CR+irxfNZ9Y0vnqv0RU/GrXWHSUj64/MEwziV7VBFSmS81VDxl94f9NgNUUskF9V
2LGNSsburIrOPLcCSkRFsO5hr/lnekjBR0D5G7yiOIHkx/WI6lFVHm/geT5+7JVBuFaaWvW+sW/k
qCKKgYr9QYCDpIf7480nsAHhb/ShX7W68xFgcqQT4RBhLyS873V4+Kh29b0aZTR+VK6aZWdT7+88
QovzXKwq329gbV1y+NFiT4bjOM4ijki/tXaCcFqKWnf7hGvTS1yIUYXIVzKl//3dXhaIUEu6xSLC
FFV8cp7U6mojG48PxyZQdi6OKkJWfmfcRZ0DhVVYGtkmmwC48CgkaJykkgYApCszOgb5GIHxJ95s
eWJyBaz0Cp/O1vMNvRsDwx4DKztKh6oSwGt3iUvlp6ibq5PXOz8rICHKPDNuFk+q2W8ATd4jx38f
PIrhFWU2IqJCoYQZEcy92v5HhU0tnDWklKKDixpW3AvyakeL6BVkbe39JGv3XaW0mjrSlpp+XODw
kL377eleSbU9HNYn9NUYK2455yZQW/10yFxskDHY5QptlP3eBr/Jx302hkTCBruCCuZQ3xEtBcgB
mdxfc/j2KGSj4FNKA/VLbqSZ2xZ3SF5btw9A4aAL5OqSLyGgIsueQ3H8ksy+0PG3PEnHH+rtA6lU
HoiDKAVACcUosjN1FacnUG3gPFpYkBg2btARP3HWkOy8XRTb/hx8absstZy3CYGeMxyCFbj6NRE5
vcvavh5N1j8kDWEapC12xuW0kMBUYPC2DeoQkpWjOueAkU/ZEy3cIYdASVFALcD68yxaUYqSk6j8
LodqW8tZdBUMVEfvMUT9KvIJhiHS60BAgD5oTrDoVcCeP2IbsAIo42roNHnApfTJMlRAexskVs71
QMtH4j2zkPm7ruWIZtJoG8MEpMcLX8YkbgBlqRpDoAXEDzqQ+wT1wKiOStRaPKs+6Ko7NKZm4HM1
XdZpgG1TxqY8phhTzqgTtd+lMkcTS6pC0/mTFqpVEYi6NaBWJLAVN0HmPa6dZEXARpLiu4nZl52T
bGIO4B6aLF+CqXmBvO9aFa1RyXtqfMy0K7fCSzvfAFqLLg+wOfNFVFtG0fuJqPoslFWtyB1urXWw
e7uKhFOubXah+jBvHNt891A0z6q/B3Sfq27r/XAD+vUfJXF5XTk/JHVcbnZnSYrxATLKjgEvUZZP
FvuTFF1NiMHUCI7C7JaiUJWanE0d9Z4xRvfjRRAztAGLFD6TbJfzs8xisa0qrDm1tMnsfsyGWcs3
2sSDv8zQ4pkzdd1JkWXnrWCy1UopwcyLGkt0//HxEV6Crq/5WweW4EAF/06qMOxb6hqBm+t2hHzZ
rIyEGHTRJhYlUec44t3j86IQe0OC7MWDzs/1lqeUROenXqXHU4PE4ZB4qAgFBLwsGvhtT31ywDAJ
9NnGxywwhxGtUb96pOw4lJfYGbbxFdR77a+5j+snOi6QRqGzlaNmqQrkoGxUKtz+aDZxOdwkuRMY
E1HzjmiNKUFGNB73bObaB3yYcwuSpcPYN37fSAaxk+oebMnYVWQBKk3JUoqsDolfumFCdjh6vmC9
XmZ60LFlmAMePO9segB1k28eMQXp5uLhUzIYKezRIlw/0bGHs1e9owpuCHxjtTzvA1vBcZp+sbnf
McaJELBKJlG9WUQTK2PtwY4OLCXSBJAib/e+axORp0mWlvUmvCYdXlamCEN7WqIHPZMZDhiAd0bu
QfMLHJcKEbc3z9jcAW57+x8oxj2j076nM7pUh/lXpC3lkjebh5aIbbKOMa2dvPHDyr42ySGGvwPK
RChC3CXabbidvzguSX0b4skUc0NSxvp5fZZPECzD3TZLLwnRk/owYNH1Oo7paYR67z+/651LSLlf
6o7gezKgxQHwq3BNyoB8OHPXa54FK+COjyBcmNyxks2y/uLWOXwXWTNkfYHQxI/d2Un9gLyEiuuq
OIxfFzfvYSSFP2Imu7mwgBVjPB1ZSRSJNuvyesZpCDzjTlgxb5VsttU2//jZBRRZ+U/uULD5UpMZ
TQonaS/Mg9KWGYDpe1cy/H6gRa52f43ntzShIddr4H/hNS6Q2v5xa011kz2Fdn9pvePHE6bf/umc
XJeyWLWbAovePZjTowBQ4b7YWpWCBcjGFRd+8o59RWorZSu1J3uKPpWdrs+5oDXOkAOrYgwt5Bn2
SZAmExCLv/noi+sgFiTUZORotzKYyh9XcpY9O7t3G7RbXG9z5GBFVVHoPbr2ms05C0RVvddfgeil
iM9lZD8s34kEHDBKVcu//DI0GJv2O31gJ6QjkEbKDh6fiaMcpXwJab7h6CnBhbehi6TkwDVFQoJT
O+WCKeHVUXB8qUchkIDxpQDo8zPSlHIWZFwJX9lR5HWyszjF1S2DmdpcBGm1bUWhMzb1INoyTb8n
JIEUA20VZBGGMduhkg8PaHgYpQJsuT89o5nNWBFxe3IELv5zkxonx2AqBsmIj+cN+/CLIVYEh+eg
XyjwcPa8l0MIrEiuq/KTgX8ykuz0hdyhw3xKIfS25C6O64PBCMkVDoeO4n8COIJygp0fWUOU+//u
VLbQTkRs4Icx6JdZqVfAIBjw+i65PVCaPoRT0zhIDCdj2dcOtshWgB/hgsd3J+pilY72LQ4/1+1x
WffYE7R35miENMGziOl00aKigYPj4bqS4RCASUdq0aepNqlS2bX4L6q3npxdj9fzAARLUyUwwUTK
LxEYiRLW6+VT1XZdrx0b1L6antjzrIsJfoJnibqKqewzWAOZoiTgOotjKYjmICuoImij5kVHcUc7
3hWJmtnpjWk3q0fZZWYXFmH7l2kQQArlGWfYkyjztPL6Oou/Pfmiz/iAg/oLr8+hFi68So0cIOmX
5nfpl3Q/8ZYTI4TrewT4oTRQEQqlW26hnIkpkPlVhdJ4pFSNA13lnZ324msfAmWAXPM3GhVXw+Kd
slx6KUpX6W8uNbCR2aamc+rrqogXMOfC/upj4bxkzbTfsfli5NomZJygMDOVdfafhAvIbos6Ts2H
u1xCqM7417vBP/S78vmjcDLcod6pgFtF9P2KMA78Mcza2ajzZ/bNGMbFXpKKq+/0ptDOj7zRCgtx
9TSAfWCX40MmsmhP0ZQ7Gdc1MX5veDe2Pw02KfZmHs+gOqJ1wFSZm+Yk9ez33noFFO3xWejI3Sag
Kn5hb4/CKPGeP/SkxaDl/gOrG/e91nBje+fn404l8bSKzvtxG1uXDp0Z+97V4v080AnZ3kcpHSXH
T3dbyp9YbEQhEOCF5tvbr3tr5hyje7hHRsSPEiAhymbmueTRkbriy1cxRuaQra5E9pcG2ogsQhpx
b8cw8gMz5N+JPXKiGQiez3dj1sfuCb5mE0zSK9ZWL1rdhp1R3lkmmjwym52qUYv1Y1q9DClErj1v
YhZDVArZ8nTI7ldlrDjItYEoA+/3pJ2Fu37Ta/1uooZWUVZhY5ZdocwAiBb+3fFwkto75PlQNdIZ
XP/RyodY+Yoyc4bIR58wC1WfXPXsvQhnapeepTysOV6ph22zwQR2L1Usb1g8IYlXlHPW/0ckq7+G
WyyZQjur3mE75fr5ikdZ1BQNUf3iL9BIBsIl3GxJvJxVbpmejZ9igpHMd8+4cXch7PcheinWGC4i
ST/ejh8lUW9kvGocyXj2b+1V9TWbaW6skl8UId8XCo3AfEyfHXum+NZTJ19rIy9p+I5/A6DWOSm1
yHt141Fgz6bK/+iwM3LmUGX2w/ujYHOWbSfi4Wkpaxk/vCyG58ey2Q9Gobm70TNwVZ/0VHHo1G/s
eMSCZ00vdcc2izOPRl4V2PUOxrfnyTLnQkf/1ER73pHel5SGL0wQSjslaTdAJ2ha0COCoN7gjGYq
XDhbrKMMdOozVvxHlLIEq3z7xZr92gvk2ATDRSVJEknB16PwitcTfdwgQHRdrzaUoUke9Yy9tLHA
OnPJpfG0bUbWmuD6lV0CBnccZ0fveWWztOV6BGk0Sny7x9RfzvLS+uyRGovzB2bRPIHknp9KejCz
DErsQyS99ie4+bAj5tmnwSXJFmOx4UErLP+dxk3oEWTrjncQlY2jFfvzeMpLhsVXcf6CVSxuf25l
wLxIDR9g/G/edlabDSGfrd92IZkaHbCHV7BkPUlH9c8U1z5DYjZRlhVRyGdNVVO+lbkW1ylySnlI
ZSnkd0rtwM8j4YbwGi7ZfbjAVuYhNgnQXA7IZI3RtR/ynb2HfvLaJh/OPZpBpJJFYWj/qvqjDCMj
l3gz9bxE7Ke8Ob3++mSx29Fw3fx7qPMVzA0GS1MYZ3CeQUv7b+QVttdIkeE+fgYPGoOhxUZEQ6Bn
8l+YUJiU5vCSGHQr3ylxgf1bjPb75uiGqTNfBfOkxAMBU0/iY++YFBSAs1OVzT2D/pEV4dlt6GfV
p9aUm9UJgsaGShGMtvwFh0r11YqDwzE6/Kfafja1rnDgSDPFD0G98KPAcdA5uD4touf6YDBA17bO
WMnSTeCedRWMGMGOVkZRI6Fb8/JprxEv5yqctk+b6yFflzmodRnsLvwmqJIpf/iGDWylVV/iGKxz
3SkarL8BvT8MfEdDQXlUCj67Yf1CQ6exsTdYMpxkCWznfUW7eTjHs/V9XtBFZ4nKJuoLQgKNN3Qv
YAjIYF/Cy0oOLsWFGvDZtGjOP38PtndwSuxblVZv+vE8NrQ3QSEl/tcfFlM4JCBzS0LLzL3fe4ZC
xHJOhvY20riNnjIKDGi58CibNrVReB28pUrhI/Q8joTDjp2Tj52vmPKojG8Rq3b2J8vzCLmEvuOO
cqK/fd9mbecshYxnfa38VCVk+th/Ld0Bh6HLl+vT2TwLemxnAqJIIGSD7F2q0MqORT9vkRGPnx4P
r+01tKh4bFmWsqfEiy7EzPGQQB1iWikxme3Lnxy0jFJOx11d39JOGV84iBfcPnHCNv+VhfeQqgYz
q6SQ1HKeDyyuh71yHVVkCIVml6I3c2V4EyBWiGbhdHXTrulxCxIcFoaKTEUQynQ29kvHL++CxcUm
l45NNhRLqJi3D5GLzQbAQVPQR/2z18cEGZDQZlqhUqhGm8cRq33bgNAUE8zgbMcuUAcYoDK95e/7
q5cp8ugnkwTt9435sGHFiqTbC63OEFScKJD3aYXVK1uE4v1gLqWbkBmgQkaYJGQeDIXM41Ia680k
xInCP/pGJ9Ix4WRQf031UEzY/BvV9kY3EnJJc4Nn1rJ3tGu+Ncf3wKpXOU60l8fbube68K3dUbfm
ohpsgQuci2xLAT0m5T2XYsctFsQrDuEC0ZUX0xY9TZXxwX283nfwP2Q1piqcDdUXzVACvImwONiR
pVXqNGTuE4EC7Qfcl7b9BQvuwA/AndQppEGlrsHrBBgW7Tt1uksqnOcvXy5KvF6DAt6lO4kD5zh7
BPbg46FAAc/atcbLV8KwfbIvxYkehwl4qinxQ0deL5QJxlbQx5i5TNnCzIN0i+tjGhM1x91ijVJZ
IKUufdcwSNX2SIsClJJKM0E8C0wk5UUvaAzyK5RCkimQrVSSbHi3qBNLIl6XDiGMIyoelSTJAqzb
+QBo0X/VESiEhmPXUqBpEQlqQ0Wa8UfKnjoyhTUz2JMRzt2juboHXd01NQsUqsQlg7zIELVEG/xZ
GbyvhHtYkatZMYS+KChfe6TdsLFlF2XTUJkJJSBBn9zwsISdqhvxedSOVOItU33/mV/nGue2SzG5
z5iVYFuvrKdq4lZYvcLKGWsO4R2kw1KMgGyoMvktQSYnlwTUN1H6D6mf6yobZBvWdA1pVSjzLeLx
klXU0tM2y11EwKnQgk688BKyc1ea/LvdNL3JTE9FXk3jVh3t5KfRTQKCpmao3U9z+A5944t8K2FV
20W4c0DBMhFcqFCu1sxdVXB/ey4ls3KESlDdbKyUlt85FC8ZJ62XEJWvXYVFVZoj6L6xD1rxhMuY
SGD2lV7UCaNnJlk4/XNeD1Z1rV1047YQiP61Q/bxLdz723xTRsgHczEtjKbaqJZW7EEZ/+J1oqco
LCcdOpUoA7llTgNZpQ2HroP81m75swgxuX9+RoV5ZklGDsaFkAx3Q5bxtAsUzrQn3+duLSLr50th
cCS24prrB3pe0JUg4T5nzRTpko8sPdxPAymzoL045gyk9ets/Kyk0V69ydLE8Oqsk3bI5Hig+/6R
Ys9ThjRwNLuuUngD13K2Ahj3i+lSEmVHH31PTyHYoStY2nsnxPMvZQazSznIUSXj3LiZjNw3vn8d
fvBXl++dDurgUTOICiHyIeWTwGSZg9cNXcQNuewT/yIzQQdYEGLPvl0VyXSc+ChTjQziNMwleg+F
1BqvTEETYMYexUZpxMHHxe3A7zO2R7Kx18pbKjVSWMlXHkYE9/GVkgyVusnRpFygzBOpMTWrICgX
2S5j6yZPjTLzMbuDli4CwJGnV2NaPV6jYfbYG3A4QMfaGzHE7Wy+KqOyNzxLcqFJvGvrc/Jdq7vg
z7i6PkhlhCbJpltMnCVEZTLq1zrGL2MJva+JNbbnHJAelKy1QkfShDQxVMwE3LQ0s87F9Xc+AxWM
eeuQM+hLmhGqUFbpzq1Z7PdJ8r3T0s10YmPwkXdNdxOIS1xyUxDpOuRkc3HF1csOuAiMElIVS8vq
X4lwmWx3NYet/aCcZ6pkx/eA2npFne1B5nrTwkPUVuWPbUROCfRXdzZZAzcqP9vd5OAUfo/Uomgt
zpqQhVBnCSusiDRZt/dpVKkoujtZ04Net7w+J4jfTO0af6EJpS2gPdAzXhLFNiLltZhy6xezBCJ5
xN4QmdaOyIYod88ZntZNJPXTy1VKbOzepkdnr0PxVC/QLVNhHlv6ocwuUWJ2bXZ4wx6Y+1/C6XbG
6XciJfiVryeHsp6wvRI0FpfRi//PJ2F1TLRp7gGhkvSWgrry3P5wb/3pM0azJwUO3GbvpOgivnt2
20dhN2ekG248GDkm/i2uyxdSfcI8phl+aTWjXDIuz0yelpAVu2xktb3XTOidzN3NWaG5EYBNitlk
7Oy6x5ylaJtjhz0aVNkTAfREgNp96E3Ly1NZLkvRgtpE5NqtVMtCy981Tj86VlEaa3AqexQqzy2k
0ELRzYYxs9WmBdudshQUIEFyA0OvVRKBzm53FvYaFm1Kk+WT8pgRiBnO0le9FBbDRMM4LmFCHW0l
C0vpSNGW+3XFAHUx00tlZehjdIETPIjCqB0eL8Z2da82+p5tgC8bUM+HmX62kJfekJohvi+kwYPH
iUf7W0SjTRYqPLo3xqjLAhxRUVE2gbnCVUCV6DOkaKPhJVibXneB4rBj/m6sTaCLTTtySjd9FzXN
zx3VTmkgbzEqteFF+bNLFz6QY+LXvgq81T/bl6eaCTcAdjL0dzZ52RSKQMHq1QDaABDrZ6y/r9PD
vAnIaomFWmIev9OUNR7nz8Ycs4o3sCDJGW73nG+uF86KCiUuMRbXvbOgLvaYa8bVSlg+HxJPUJAh
GlXluLy1uthr2yBp+9qGdbPbC4vP+ehxvXfA/iDZioS3wiLzEgh31RCNNxPnTXVeSmzv1ju6pcKa
N1LaLUoLA8sBRGweOPxP09RBSgO+9JiSFex00vjbRi8gkRB1a2s/4BMhko+dEN0WhddSNvUhri7O
Z5JUgcdG9q72C9f8RGiKTCkABgQqieDM2/o0sqlQYiItVPtqNbS/tufNdL+1mxDpIPBSH5z4enPo
BjF8UpiEsfcxHZXEj7p1Qj31Ty/lBqsV/E5crwybG6AVRe/ifUtNpY6ieNP7qLRm5Z9PNEqOQp/O
w0YmMqdTbLXYOBrksBG+R8BLIGTMl9QR6MWfec6PSS2JPjurJu9O2pfB6rKpx3++eDeAgrGafS4A
1pcQt7BtZnld3w8qKTswAIkgQ8/RsQtMuw8K5JNCqeOTvlXR9a2tgASjAhSdLEeN0bmV9qLgsQxC
iYSWElo/8dsvmt/jzP2yvNeh1PW59IRAjP92fAuxvGZNrQpN27DJhUDGG4XGoDlFIBShO8R3iqn2
Pz1/hUWA2M6IZdvKnhQBPHx8obh/j6sQhCqoKl72BFvS0TfV6jB8QzrBfD1QsnLQEGm810mkXXT8
/VD7stTMKnMGrj0vXKfN/TBOAL4l/saQo0KpXVuKtmdOf7PQlpnQ+WtGJVz8/cWDH63BTas5R5sh
CzJx8pdea4gwACpOT5m6hJGAIsRZR0hK3eYu3qpvxEyAUX4NmvOGdfqxsEdRduwfRw/4YX83p4Zn
zR+CE5A6B70SuSyR5hjzWbIAiQUmUniLcAha2hi2kkxKW0qraLzza6sUUJLlHltHboCkf4CeGeHX
YR2WkBwHhWFdMETWyJzyMV1T++2i6itOcnMw3pxnpZL0iUToLDoyuujuutIQQHHjDSKJXp1l/j3R
RdHAYqDrVMn3oxy5tM7KHJsJ20f3kiY+uIRuEeQ7Qp7blc6aYsWqrUIbRuHgCZ6RDv7yXBtF5Ibk
35cSR9NpCudx0lPB9aS/ZuiXg9Njmyzv0EvuQ5xbUIRtPjBFs9oRuf8FepB8MKlar6dIQBIwOw2x
0sXRMqNtjLRDRMG2rhsg3V788NA2n7N5JdFmF/nd6mTqHNfzM4sDtTfYxCcVfUnTx6ulMhLfDLJL
jPrEMqE02lRxVlyHNGOiAs6rJ1g/80kfeBctgZ9v+AdiPUWfVwazQG8s34bLnOWdzdE8Nh2kytiI
IxE9q3QoIPdiI9Q/fMsAefmw3dM1VAEZoinoyvwKq1lVLAQY1HmDdZ3MKgIR/cMH3Q99gtBYEyPK
BgS2e807sGDn2Hk2RBufdYyDUvj5xPFFr7ipa95q4Id+lZRJalCu0mow8eCwXfmoqazuO2zA7kfj
x7U8r6R64M5kazfMCF2V8cZiZfsQ+F8PSpr7KqsZA024ipd2xniL2PjckKM9iweGDC0atNpRP5tm
BkghUjsBNfEcqJm+5sR4lDtKiMuuoOsXILxF1tHD663sypBhP4mFrg+Van4gfsp5AvfDCIzjYc7m
mzx43mFQ2dmx+wnTKRvReWyta79bjdlroIGzAArVP5r4JKAkRnynH8pYAbnrfNdFumIFKWq9nqXc
iiGZ8EPl9ax6bDoq62zou9Tyh06iarY2I5aUD5CAUUncZjoq2voOdl4/7tvTITlzmJxMlIgKd9RK
qBv4mrklAG502fwHzBL8KePt+gpEXIc5gRrMTS/u66VEKXXDBLfg72xOCwk9/5zWyFkU5sV6eL3r
QTZ6ZwRYFI7/te/Kd7xSWTLjXbplW1ayQ4DS5G+/ebILBj+NjeZn8ASUsF+XFzmPx8v2UW3ePwBT
mGAN9A7JmyQ+3FQGwc7PdqJmGcfejMPTabtVQRIHX0ian4uCQJXkRs2Um5zPzyeCx2rils6PJQWU
h+ReJFV+cazS6O0f1q5ZFgPQwlxybdHjwRFEi60eAl7Vst773Ji4Js6jUrlY3pPIg5FdCSQstRII
t8kRPgutSyQXskm0OicnRzoPsmeeFJUaiqKZA+u5mCY7DlZRp0WFFy5kG+6O7osDHnBVAWUeKwrq
lMSayldALYQs7lTSO5gNfY2OJ6EOHNEMUs1ODXKABQZ9mtnygBRXpPK68lY6zG7v+X7ys984ad87
irXzmGWTDSMFlag2fBmeqlrWdJXD3FaNTd+RSFn1KRFh6uGE2bkHWvpSgfPdsfIE+Id3ga8gREeA
i6CaZz3EyP0o/0JYUDw01qOAPes9NmkN20J/LivbHfRAj1G0ZUCXfCuEOWdR5Swm8uIDn1+xFp3t
PPj+7V/D07rca2815Te5SpnOusz07dF7z6JCKLF0CuoGpp8a1KfHTKvdBebGscsWy7xx5wkKOStb
QAvoc2bfOqLyzn2kLyYaYUS2Kkf3x7PtbYBDoFlbMuvQzKF7l5+8vYizsW5eeii2GFga441HRPhy
FUwC0RohnEgj/qCSPxC6mkjV/G2gXLmiqh84F5aWtWEEs7ZrrRBdu5cutozBe8hssQoLy5d817GR
PN75T+Uiy/EVxoZVUyMh77rao8ES7C9mT6fvNVZ/7JhfkAsc4Vkp1kB1ykLyfS8fovvjw/HPLCui
MgAGlJkB+Pw/Y9mYqqMAAeOVcJTlmwQnlhYALwh9ZWYHShf/MJdaANmIYXXeAG1uYaMML0K3P6Jt
l0p7Qv2vsvRuNNC11WyB7wZjQMk+zkJcrAFLkxSOIxxAwDlLrKIa74vZAQEDMupUz4z2iKmFYPDZ
7FI5xcQm1fQ2DoxrkzC6YyfZYgT3rNk6j4rpMlSEkDMC8l5Z1EBkMryrASBbp/jVA8tEC0Yh2ywo
sRoCTc8THLE1Urs3jb8c9kmhFvMSNfEXZWa49WjoilPwpfVMkvVNGz84YpPeyTZwyldeA7BvX/LQ
/y8v880okwJwvlJRn1Ga24LeSznHnVcgbWvI2XYepb1HMZIFVpbL+Qq3E+qDhbAL1A5v3m9lEjOy
ToZY4/DLYs292r4e2SVZl+x48bXdyN1ADBK9W69Ge0Q1m2F2vtBIGHa8S037B6rMzIRJpAUq2I8S
U6Y117gJIp4l3n9N3gQrwhSLlUQk12SVpOieeRNaTQelEnF20QOdcP1lYHlRIh/VIs0Q0miPUgHX
a/w4/wthzq3k2pUDAgs0utesaf2gqVGgAHxcPT4LdLHIJ8VmMF1iMMPpOBpKlTf5k4P5PlDNONFx
JfHQigwS8ixNnLR+55PrcY4JUKfcgm51m2PEKREa0EmuZ2tNoaNP0dteMo6tAsDGbhOtqCwY82EN
DFZrlwc/Bb13BX8KPo1/3GSh6YSataUMzHbEwG1iZoZO99O1cvIKrWVeD5CMJ4cO4hyGyRQ5a1bL
149G0d/vmLPQ8hSM/Bvm4KG+IIH2VAM9qo1sKgG/fOQR5adttM5L+Nm+A3H3zf9OKeZbJteAtLh6
grssOsFCEaZUG8L/hjJgFdx968lmlm5UlQ8YqD+LyvvRrJ/IXc/xKNfbDFzkLxBOryh1r/M0usFN
V+Tfuc8Hlb7gXM+JFW66r3uoHnRNZa8oec8DAGjJmzGrsE0W3OqvTFEbdD0wMLdcnlj5adMm2b+p
a9y6EJzlqlsayWuop7hvqkUnbYNmpAUjh0i1Y/u3zGFBdiMdsOs5YenKWBnwwtTrsd40SPDDVVO+
S4LZFjoDsKkCH18yJovYurVLboNwWNYCEKgBJyQE74jKVK/FzJ8y8HWC6PRKL0mJynWUiOVVoZcp
iwZM+JiZAQRp3iddqq+5iRMf9H3YO/2eUAuvwBclV4INEW4WZFjUxSHlo2/bWRBru37GicAyAVUg
+3GOWdvCUfxeBanSrq7vKl/RcfXJgDagSQw25jL4CbcCQ9oRpv/REpq5dP8jn+x2PKwgRo5C1i68
2+Va/FvaIwwjaYYIgnDTmxM61HAf+BbOibikBiMx3LLY9PT0g1d/tC2ZVuhIOL/Eo7caue+D9wcX
gY3Fz/Q7vKyAxuu9cgppdKjQ0H2UdCSAeZ5VkJQikZZz/YwOVrFS6fLG39Sk/YVkg/8e4Cg28i7k
iwKaHWFUQML0XfziJONAP4ERsJ7YIfihaCo/ASP3qKIu+bpru4/30VbCitIHTxABM8chiY+w2c8d
KcM7noFTqgR8jL/PapkdA8OTD6080KLjbZpF+5Cb7DEl7zsO+4DEFc3017OzjwUqI2iHzA+SDJsA
ZNkVCyfFMTgOrx7wx2IeDl2RpNl5U6Ed1K5DAdwKpE9/m2MdQcf49RIuBkLiJBLNc9w2yaIOIQfZ
oCuYGOSuyGOB6QB7HfeSA/5S8Sua1P5ym1EMm6xV2WL6XzqCD3pAUp3xMrhG53m+HrY0GpK3ScLB
kfbCCMdy/ZxDj3KHQa3xwqZsrGJwaqdDHu+OrMgy+rujMhOxJjMoVf0BhvYRaZbg93c6A8ixQzX5
VC/d5SAPxrkTLEFTLae1nEKbq3IOQwRWaIrDdwWGtF0/2eLOw+NUN+yyxtUcdg2BTp3bSrGFUyHA
gQgCWOH++AAQZJ6qSTFa4F5ZuTOUc3xuRcLehegCqfFfrlm2rXNWUETRFy1HEKWpifL0XnjhsUr0
5yqq6fQ+fNEbeC7HY7hGc2QfM8hQjqM3O1YZBnBCCKDEaz/ftLJwjolRhHmFj9t6q5LjvDnQROVg
Ezup65H0GvqOkVKcXmfOjHQa9URdxplFBHkP9DBKfm0SsUDaGkPtHg/bqE34Ceia6BvJH0jLkEmG
bpGyxJ+Ui3QKc17visbZGgWUD7DN0H/ytJh6ae8DkD5YCNIGyBmcTPXtiC+d21jIiI/L50tn3qAU
A96eHzbmpZeKDRRHKaM68BihrDDjsNQ1WshIM9nk4o8zG4H8YmZ8a/soX/h/y5DeuQDMO7RRGWzl
cmM1Ty2T1a76LYQ/JLsKUMwK6lY04BtnXIUxFQQk5LUp4AxzADD4hXwgPPB687uVHipQngfPZI9X
oSORY8Bes1qCfdLcd8HuY+gVUpO9VtRXqXf4PlLyLk6l4bXT7uct6HmT1xGiW9g3OkYP5YUWJJqe
GjTe9TtiGPAQLpTOd/bnaRc3BsqCIizxC9PKyUk6wLSAtvDf2AVmMbkR6ncqz2KI469JriHw1viR
cYch1MXSgaqqWv78JCYa4dTUovsiP8+IRtIcfDezeaYEeQmmCoyrV7IEParv5MkNW8G8JzK1ZxHV
2qr2QNVteCqtmMTu/Vwj2wJW+TMybqTRxOr57wSS9RlY31JsA0QN2/mastE1PEv0YkJ0GtYM0FUZ
rnrpkPMfpWLHAekjbjy72+wsxiW8N2L2ln5HB9VyP7zUhNkB1qL3cYHdLe+NCoGp6LOM2s7DHA93
Wle8dLOGi4PuxL77h6BGtp5dT7V0WWiMRFrp8aTcJ3EI0CSEu6PRQrrowEKK27X3q7O5QRm9mH4V
Xe2+WooXDPTeqo4s+do75wO1w0bmGWQ4gjoM0vGs5ssfgaH+E/MkCy3zSuZoB/7vMeE5crtqz3NY
qSfkkL2LXMfup8pHPYoSYmXT8sAXS6VmuFQUq06pcKEr+yRBSE5qF5v92Aynt7MBZaWPnHhfxRGa
NOmBTXKMcmrHZSoxi5WM+ojnGooq1Gj5LkFcV2HbFcwvlRATA74fKbSbTLK88mBrDY0DAwjSr2Gb
oSFjeKsnGSc1G9GlllW1ALqmkliw2mR6+DoNj+fKrkUganQ6sbore3uQ5bU/0b5We9h9pruyp9SE
KGMDDbDT/06MUgdF+1Fj8j0Pipa84LwR/USwmUEB1nEUQ0pv2knCCAddRSepYKNEdoHUo19WmMpO
hR2W6p5i9wv9Wm/daDznqzga4wQawwg5KZm72UkidVHotYDd2Oy3cfhtu7/DTAWVd7/VC1lCYQ2O
iiscExZtxgjEqsS0oznJz0cRgrUe1CsKc1uyqsIes7Upol6DStJvGnwzDTt9zoqNB5erU2pZatPp
eQhIEEMDlcwSzp7J6senHzmxGVmThWUlIDrpap+DPK6w3L8crw+p8eB5KOVq3MfLmR/6qvXjdi/A
uFahze8/7aZcLQVO8Dmg9/7ddTIevKvN90Oo+QtPVIRFW5nKs4+A4528cI41HTrGphtNriw3Np6g
j6rostEQy5vlLsCuYU6M/F0KI/RBfse54YD7iXvhYA/81HOK980WBbw9Z4gc9a/GvEvm/6RNc2qJ
w9C7vlQqN8tWbmXwXGsSKZ84pnCx5TwcbkHt+Npe6qS/2niNVUFUp7xRt8ppwahlEt0+HwwiLTGt
BPAxEMRN4S7s4yuF9hSXV0RR86/mgAOsXSI41O2Jejk9BncuGoUuas03S04BvFvuLzE+yZVNFikL
INjluUc98r/DxKMcualBnMuCk64zWVCxra2nNkkbvWn2v8OVqFaFK/whak1xbBWQLdHrK1y+2NdY
UrW2V3iL2oarlTFgC9vkvOtsfOXeC/R8XqBfHMLR0lp9cJ/GsYu6EQVTrBXeI/QpgBHI1VHqhE3F
M8nq0kwenCsGnTNZ0Y4e6/POwxT0JTYSXL9bZQqM2W9GsEn7rxHbhkhF/KwX4VG7jSfPob4FkA5z
SKuUfgb9m/peitN57Ij/0HWWr2eMqzxM0lsEVe/ZolUtdnb+bex53pxdchrHCcPlhVGe9IgzJSUu
uaQ3sd0dDVWvDAs/ynVqqKyRfN0VSHPNUDhxIT4Cwiylpgq/Vv9/nrNyTj3YFuZMhxxmxaICEtW+
6gY8S2kB852H7mFmegZuQqedcGRdjcg4Q21rxqfT6C67N9oLvfEZjbuU/SDnuIbBqN30X+AojEQn
psOc7pZ+lw66LKxgLIk3xbNwJLbq2JAdYP4/yzPJ2XqJeCM8MSugjEZkrVtJb8U2JJp6Sw3JCcz7
Up/ahrEh6cD0OHLB4gOqOz+QBqyyMO8Xxg+MNpuEhdNZCIj+1O4GhPvXIlZgFB2H8blmqGleIr1l
GnquHwb/eYHVPXNCJbgqvQ0Xokqe4/Mn/1/p2cxZQNVlwzaOqi4vbEJYJ2bUb68+cCwVJYLN+xIk
lhqDDfur4Gas7lgm2WFGfbMDySwOa+kn8y4a/FM+oMQCIlPstrB4loWAUqopsT2f3X3+iy3MyU4k
xGPJarhKgKN4Yier7f1yhA/R2oCeLjZjGFY1jgtO4SjygXvC1PIYRq2rJ52KE6RP2TCEI+IhV4p9
8rSQwOQIPHzdh4IYv/5Iao3/umxecDU92PCDTaEqbjPt1S5WM7XFwyZ5HOd05VbbzmlpfjLszqIT
X4Ay0yXOvdoo+msbc0spptuJybcWWLa1UJXZEc8WWjhXH1xmtySOOHBssPsLm76zB2lbtXBNq+hD
d9mLDWugaocTeJSbR0O8f4FGKurRkpt4HudGfXUSUckgNn6IlAnHrPGn2BphBxML2bbZoR1d26C8
imgaigy+YJAwPEpojYOJa96cJVH++AMZEwoKYoG9WVLjq35G6YsYEj7HBa4eG0+ZYaV4GbKzuh+r
5pQ9OFP9PGsxf4yw4K1QReH3Js53xubbXvyBtyoMK+Mddjs4cHEVvZ+QJxVCLpQShtCn/nFP+Sqx
NyldrZ62cFhPPU/aHVhQytCWkFsJ47Jn0MYbMeTjO0bsJPYVRbXCiq0Z9hJuMcDlLPqkAElY+svr
JdEL2UCrbem/m/iQUCs0q8R3t05CCdf8tE/Vsqjwdvr1AMda7N6/XJXJF8DTSEILifGoZVynVAEF
dCicyv2VOdY3EksW5/SDz1PxbZDMiAqFzHLFUJ9Cf+fJ9A/CiWKx9s+el0mywoyGUbaKA/YppoRr
diE32LH/UUxmDfUMNAqpU8XzZNBdu17KmTaoFsK3QCrx7aV5bg2KdaGnLM0ijaoVchK9wqVarTG1
AeSq4Hp4jVhWzqoHhmtqVCwOdP99K9X/5UU86S3CYi/7nxwMUMrc0xR8xlozMyh9i3AtyJ9guEUD
wm7RG0TTYd7akoH+3Hw7lDpF+v15KeaWUZ0eEn1KixlrX2sdj0g3ls8GgqYOHSDm4nkEriqEFo6s
0qzgXcE9xa2sXGxUxF+u4buIEIdsbsXM019oOX4+D7v8SHxePSKkoIRzbvC7qm6cOECv68zjNsGb
AJml8wvE1CnQ+0L+bUhKCuNk/sLzgQ2C/W5eoWc+noVeBUYPh79JxDrTJUeGnlGeRaFw3p9q9yfr
jbrPK4gJA0q3lKDZAOrhazutVpavdr/U1dDb+KKBI2Ku1hSeua4Fs3v9YwbqkSej7qY4wpL0fZhQ
C7ky72NyVlFlo0XG3UAoML/jzsAvVgd+evHVLs+ocj/AdSs7drzRGgRDOgK+Fjbalvig1u9UDKhm
GHXG+SruxkOao9JOwKjXMM6P9r1u2p8YtKCOOlcgmNSFZmdYRnJ8ysKZ1YnLhtjb8HSH0SDdIrUT
hBnVXmXZXNKqhw05KoMOHYaLpc5G3qetpv/yEGEr46XxV7fZ/URiDfHm6PzNgAcmSRUtzT+XQfP0
wnkIZvSrC1Se05EjgvF8r3x7KTlbj6/JNakj4HuR3BOHX+Jrjotv1UpoxIC7/+xL+/N9cJZ1ie6E
vLV9cN2WLGAQsNO9vKX6Rxcn2rCeyHi/CoWsayxRQCoHwTPR+UqYUTdP8HZ1TRC9B+IthjXPHpoG
RfXSgUuhbXubSfv7a6ZY2FmkhCijhGjU37roA8Q1ulO7iMVIrnXNzAS2FiA9dpShBr1hQ1sY7Dju
KHnTWncLRLgwtbe94T4p+T6dyf3Jhy5vejOX46zIqtpiceyDfYkAnecvsOZkv8W5d3EQTqLl8VDc
L4fiWaBqyDJq+dUaFBm/uaLt//beS1F/5+29dUZ7DSNEV9O0awFBqhXl/5ski280sYjNlqZHh6gs
MPueeWkoIgH+XDBGqa8yaeSHE3quiWGUH5J70qdOn5dQTeRXQs+k69VgjTkZ3tds9KKba3HI0Lnm
wQcmenxvqpmeQfwef6Jr76KfKiZd9ZRTelEFHX1ggS84nLmdNeG1qw7VdXUwQ75BIOZBVdubg7yQ
uoyXf82dI1NrDi7OAp37wBQQ20ZApffcKOnQaak4wZ07VwpeJXzZGxgpngxudbdNT7dAWlRVgQxE
D0jp1n/pS2AIf5hf8ztHVMLZW4BYySF+yJc2pyN/IsLi4GC1PHc00MsjwRB7QSdlfnw0GqP8yzKE
iwFy+UaV+4zFGyj6XhEB1EkyNjEAIkcz5734ffRtiIBxwjFxi7+tlduoGRJStT2qI9uvqTKIDBd3
pGHPL57BrasMg8nvsJZYYiPh4FnA7Jn2DpHKz6Vu9j01fmZUqrHFEJsDpR8r6Il52qOobKBCLHl1
IRcrEHbRCSsiA/8MB6E4sMYAuDfBfmWuFY7ReqbdeImBY/iBLstieVyWBErr44Grn9zo7fqOzTy+
ejqFwxN+fLMBEnAoi+Ityjj7QkvXF7HNOo2SDFnmVS6CbaRoxpzlz3wrQEIfB2CL8Nr9Juwwdrup
e1hzXX2MNCv7WnGGqbK841dHvrsg1aLM3KNQY/guW6vLmm3w2dAWH7BwjzyO9qWQD1s/0Pvm1AKE
vvCX4Q9q5B5cXOBQOkdUKL9sdCGfXM4RhyJPJhM5+iMFzHLVfGsD9LNsyQy5+guT9DW+sdJzgOyt
HpAUO1TM/i7IJO0Az7rDx606WH5FAzW4mr/Vczq8VElkDPIYc+clLvotT+/IMoT7ri/J8o+fjkAR
IqhSI32464rpn8bK7KbXlTTTOQ1qPKZBVy0WRqekzdmPUI/QIQNNo69MoLW+A5NguBjq4QeT7Knx
o6FRkHnmU6iGhSS1/ZG/fR99czAXu9zpofO0406C5BYdwOQtng4EyVy1RQ7UzhDkm4i38g8zHSlS
FNBL21IVjOraQ6sxnewGK99b+qOK6goRM1xR1F2OdFwW3aQ04oR0o4ooBRWkQ1wNbvybcVA8aSA6
g3Cp+BCG8sFNyyj3MfGCQlJaZt4wUbxFRwn3vZGpL3ytpcA+y28nkQsBoUY3/kt71XxWKnpLXEXe
h6UY5gH49VUHyiQp7xWusAFa1qrf6aebCFn4ZPULRSFRUyrCOHbivr6Z0lfBDpxdjYV3ht4mJVgw
7WjUT9iY5IOioVTHPEMRAwWajVzNYfKGIskkgekf2ypaMi8SlKFXn6uyAJuws7LRrlkYH55gqcEQ
ULE9eRiUjlkBaL+rvCZUNUA5qvMKJyA6+FSd3L4GtBphAQsGxYoDT9HK2I4hQRxMiC2Zm6f1qCz6
b5eFYv5Us1sQBVKsgLUU2tOZtPk03NMt+yMxsK3mqBQwkytFm5DNmtJAo8VV4KCV/9anmzFeJoDL
xoiMLoP2gpacUnwv9dGXP4d3xZv7vD+q+1Y2UQyU6uILK/NIyfPL6QHf/Nxo6ePERLMllYt/VhZT
rq6bJ+ZsGnLVQRMOcd4LPtocOUBlS1fudMBYGu7vhncgM7/rBsgqcwxN3rCFlLhVlPgcbe46g+lQ
N18AinDQOjlyY2w1pIlQ4amg0KFILxhREZdjDmKw1VVBMvlJ2qg+PIkMbzTfp2Hw5yvOr3KHOc+Q
befX8QzGDGTqsoOjGgZB9U2KbFeKeuuaXtAtWxkO5EOjbFbIQ63JqLNgbssVyPNZJezJLdhr4+5P
/ih+Ie/DNse7tYuxxPSY3ycYiDkd7y3ZNf8JptAhUnvJUCKPXO0YadhEYk6N9IRdvNKuBcVWKe3Q
91zo9tANo0WLpcQlwUGWrV4ki10aOe3YW5md1sZgqonRzD0AcHpVwZCImGb/3FofGWbTnhhe9zto
agsSkTjGqwFNYF+2WVAXMM9dCiKr2kEIMogL2rIBRr7WVIq6Zbtl82iPJ2PTYWNKZdb9nxWBhg2A
3WYFwSrhWnF74LB/yYZKbrCXwj+m704unZGh1b3LF+8jlanl3BKJAftbtKy+9jAgIHQtSKEhv90x
d+D/WY1WiD6qcsLinyXsQcTtCjT5GSBbT3DWXok9vvA+HlCzsAda0xy28WeS/X49IFR5HaSlUoNs
PT3jtEvfUgV9SF2cVOC5YBrav6f13nU/JSZiQgHXBpSpFUFQ76qCIoJHxb8cs5vCACdFFO3hU70W
a1SAUkuxD45XoxQY0+yk+AyoDmLQoZpPnRrf2QczDK2hoeAMCrSl3oEnM8Xf4inDf+WBntJzaYNN
JoF9dAgzPVS7TmW8u9UItzLekRntV7T7MBDtHS316x5yqXNVO4Lkp5+SNinYsXvcQZfywj3vou7w
0WfK02iH5gms/dRVy3UMNBUJrm7wlCm9IUd+EBwnxG/3GEWPpdKc56ufbRYXqP4z0+9DjJ9N9VnB
oenCcj+k7kUEtAWXcx7FaMUdi0LnCDk4CyKzk/CCjcpsrj4RGiLBP0F+aS8Mu/iSoxLCsYcPDSja
LYk+wWUSXFnZeXPPvKN7NVqCuyBJ3Fz9nS+JgmUrWNxATBaq9SOwh0wKX8tHnezphYo8xqdUZSv0
VjmJAtAriRV5OZnd5qA9iJaZWRL8GqTGLPLWhySGx6BzSQAW4xpAgXL71fn4ENkdfjNgeZmU2gJ+
BxAiEbvTEm+hpwIgCMPlX/nGTKbF7LSKXJqH2ZtjJBfhqh+BsJeSIPWptUL5jI3jWF06Yx6MJsTP
4KGrgIMN5iyTrwJ1mX6BEo3pV4Oyh+In5dwbdJLB43wRUMXNMHpHZ2tuTJbJdiQEtEKC7a9GPPXr
8pTvnyBK7m2Nn99RQLojtg7AwaOJTXVqDzCO7YWtrvVeyyAyzlb2yTuynDhEFFNU6ol2v90a0O1m
iNIEBLDf31hLdJWXiuYNUfjONhqbPI1+pL3P0LOWtAw3TJHtg7AtCWG1FHTgacAk25dUcVacU6yO
MkPkGPdB8Px/83OTcAny37K+su+VTExUk2I2BiDNMQwkFn2FyYj3ROXrASF1Sd0xUm0dzQBIxva9
OpRWrkwUCaTt4QdgAQ+5kfF0x9T1tp99YFmLPsLFu3vKkUNuOiGJu43ffMLWdhtfRnIsrqWWbO7n
D+AvbIaELGl7eD1xE6e7VAw2uNtg70gdTUiCyLFaP6GezHp41MtivNMxf102MO4aEETI9lpO0DV9
HiduL20WkLyeCHZz+vOZv21Pwn1E6IDdXhHB//ij2lAaqbVnvEAcA0UBRHAiNmB/UkVuoRSUn3/v
T29sJP7kmLWe8osD9RzIVPR25ZiD6SjPVvGcJPKLVtom77wsWtjVIVYxSMJbmMl9AnX0iY4Hsjfd
cnC8QzcOtmT/alWEh2vDdrWBY4JApI3F8625bZ7SUVPvbVqzkdFJbEsByruEPcmH24oTa+TSQcYi
pnD270QyK6jAGmQvNNGnzllFx0mCuk70m6D4jSafyfSO9atQDXKXgCDz1V3n7DqFkqxNRiPRDaf9
xGidrDpuibJOUQXNk91B7IWLBAF0ELb3FahDFDn2ajLkediAPSRSLq9Msh+WxTJAc5VwBWadQz5z
ih7F/698QK0h2CK8yDeW4Gw7NBJ1pIb6RArOTwcA31OwI2zc5DRswa9AL0sADHNqN/RO7S91dLaw
xiSADnjEMNbnF6zHr0XM4P0qJWovPmqDXjNxkJYTjqWSUvzHjSCh/wayUdpSwXKeV3d++cZLjoQ/
pUH5z95I+YnbVqxspuDAFEpNcpyTSdOnCmjmtt2WhzghD4reNdKpa8FtFjf9E498UKH91gAEutka
Zp7DbskdYUeDCUz0Y4HrfZhsXlBr7ehrqTLpATpVgSIjy4UChYuREC/HvYii7KtSlUm9hNIg1iJN
ZSww2xuSH83B+nAlWMuZ9zPBz/Z+OC7F1hBKT5IJaJQRwO0U4d2gsnO9j6gqer0xFAS0t7FCEvrD
JQ17Y5f6ZVzNwyBilg7x5OWC932S6/veIDwYkxFcFnG3vRiRBBJ63LGB6svvGd2ZKvv+NUnVAsXq
uh85P9DLHlm+7Nb1wcGxeiLRPRf3xa5ly0n/ctU9UyARdnH4Pm9tmIp+HU4qVeleJe5CG6AJt6Wy
TQjY4omZ7TTNe/LK9IGyifBu/BMHLAqP9kO1WJYcWaKVj7zE9wLP4iPkiTSehKzig/ZUTeALckUq
y74pjrSjPhr01X+VsZ0C2UHRlO9AqNDrOv15LxyErbv6dQKDYjxy9UbmA9otLViK4sA8iar95H+q
nJDdASLMb26RAWxYDyuk4CLYE3lkwwRv0J1nvsTAPL0N46OhVtLE+lYC2scAVrx/xAUEEBOLdb13
StUKKWwrerPRdny9nHPckpmhm1Tx6k+SdYzyk41zf/P85fuNc8SZo4O+hLln3xI3YWaHdkvRJSqT
jpz3Yn1MOF3CVpFjn4mRLE1t1bx/xlbLAe2oH18onniurw8DoU7FzU6ru5mEclJbL6YoVuFsPE6q
2k0jFY2wjPe6YXmN3Ok8R3pgulN9Oz1ypW771fJWIbfUJFcaoeLccvASh7r16bANchQF73RLZNid
devhUR5puYSoDYuaQzE5UeWu6oHjzoCT8rQ38VV07ppMHn4SPIKq19arh0bd5V7iozDWfQMxg/ZM
mg85E8OYQExsUZjSsA7llcDgHJnmgD0P7R4gjgl9FR9s7xg/jlrgzacjYqhEYt6hFowV+R8a1nqv
HZcnJTsZJtVF1HImyIQwqUjMi3ddl1zNYLYzeck1A9XI3mOcl4e72dSp2Ok/levkAQJGRWW/lISB
HGMZtIidv+Z4Qrh+2m/J2ISy4/ASv3V5ekUEUf2UtVT8GQu1XjAI60xfoo1hQUAAsI/NQFCi0AXV
KnWXwvo5j+buqh7bMnGj4I0v5mYzfg+qHDoTgNVvtUI5dMjyS/yec2gvIMzxJ+BR3AUHtbZ+0JSP
O8yOpXMbB4LOGDMxHPyc05N2dIfBOU9RlvOXslGdGt3RLnc7k0VLApDuM3eFasL+ccUki2SC6E1N
Eq68dpJ454jBxVuFmyJ9uI5VZtpmMHwyk0lBzqkXfPinGQ2XT9G4TOURWkdfmPlqd6g0VIBaztBV
a7cWrnCtY9nSJbnhYHafRnmQX4tqefAbw3QthZIQzFjHsYfw/iLg3YrpkhWI5UvcyTgc5wZINhVn
1xc9ysEIxcONSlosL7MnmConLBGsBdnA8tYgirLLkYlOxYrsRvEMvDsCqH7Fyng5Vx4kaGaXnNGN
easblMeBsxveHxDB51GqxbWZvKr0KyFKhcDw4QMUIoDf+NYBGKZBo85wjWxBILm/nmWSfAh/yTs/
qd6jEshcnQmgK5fEnGTrFJ82kYwHNPLFtge3v/KmM6nZ6/Md8M9IgVMiQCabSXlfxoHd5TXhrrjw
NtzmWHjq8u0X979VVc8Q879rQ+6mmeLuySi4FxWPFQjC4F0iKu4EoX1HdTQhlsNSjIiIgxZ3rAWs
NYZkwvgXfenBurzl2qYzV3gJkZwZwMefLDWdQ3g/0EL/UawpRIUg83gl6pxD4wB7pb+XwQXPJO8U
Q9ZVv37oftmJQPnDGKM9sjvmTBEIjJF4adpTFDY0oQm8ELsrAnOftCbdtL35XfyrzLbAupRptWxT
4JAcJ19jlR42k7FiqBEufp0iRycIzMbWvBT8QCT2EXAnPFIye92spv1c3g83LQ8SBJUjNZ8H2WNr
bwfduMjCDl/zd1XoK/wtK77RML8OUlK3CkmiMUjjJQeCB3RSkXGQfouq9kOp1jrYjjrzA5wm6oV0
iJd0NlDt0qXDYLHX0J4gVcig0ZFVzboBV+7ITHop+CsZ1xBH3JAPCu89k4RqwLi4W1Z5sjg4VsvI
HKAmyqnrbSI4NnPKmLx8jAKgppbsj8v69Su5qOjK7OUIPoYSjLRUi6JMIu8lDY8Hl8G2JEf37GkU
NG4iFgsMX91G23dlu3j8zQHUK6Z9c2Na0/ZOSPvy6OukCjW9e63Adqx53mbBYB0erCwSRZZMnX2K
Kp7igIMxODx/PRzsMSEHa4NPLLqcaTnfRzgfML4ugsQHyoOjOA5LtzNIW9HhNC7GwH4SC7gHeK9T
dE+DzLVralA7mGzi9TznmVaKjFHElI2kdA4jThgu0n002nuI1rHvQtkM359503pMjaReksCCApXg
RVnj4rsQtHHr1VzBQUJ8vR0hdTGu6ocS1aWduG7d6hzNOTl9dAizGnYlB5CGAVfO6DGaX7ogikPn
bKrm4aCuicaEtH/B4lSMVgzF7khU28GEq7FlyahBOiKZuAZ5EqsOEbWNdUkMVhm3/ZlcMXX6QmsC
Kmu7hCj55UOF9HrKMOYVUgx+CBfMbkbDCujZJmmAVqeNlTizqwxeElSexvksRx22cO2w1JQpaAx9
GdTIMPMWuRahA3hlBIpSPw7IyA91DtJxWINa4mDkzyHhqV9Y0shSKAXQJ8M2R9T3idNIyDKr1zKj
6jA6NCLwk84hX60Obtug2Tx56Di+6HUqV5vJg283ycRR+NM73gsJ9/7Lhl2xe3ZlmM+cbgvLx/M8
nngWMuSyjr/MuS4ZFlbN0kHmbbwp0QodAA2z/nDtELF1lLfFQMI8MtbMvOwf+RiPz0xGc23v4y4k
p07HOKQ6COjdrhQZuWk70vEBuF2VbY+ElEGujldultmgac8W1OHMfKTqRTYiRZ8HDFuiizUUNR4R
5fp9jIgDn8Fp0JhxlXVRVeGwemay3BPKFo1n5ORhakvpq0rpYFWbvp3oP74ph+ih3qLpxUdDbfHF
SFfn+w+OBQh506eqNLgAxn6nlnRjfl2dwoFSpymH9RJa7U7qg64+Kt4Uv0BeVenoMYaV6jY+JJoh
xqhosNeQxNLmL+qq/2wn5j12dB0Cx0TFAWUPkUBjoloV01VpvY66fYA2pg3WFk7dpW4i4Z2F84Rp
mtRYP5FIsN3QZfWfLOCCAHmvHDuZ41OakjDkzV/0+NkZ4MsEI0qDC2/ggYAeALbQfVUSv4nLIJvX
lJNFcpMhCFKY13qdxTQ0KsYWSg9aWPAoefjqOqjCGOywdL4IZrBD5et3riOEAt0Dcv0tmQ8q2Zdn
3wFPoghPR+9YNxXWELEY5gNDKn2z+gh36hPjHiaLPmzBTLCeGI5kYuIE9LqhGjovjMvBvVau6g9S
5hHtRVDH1B5sL0VH4q2CODZbnMKfeTx0PJvhnihObjy+tP3vZeBsw6aXnfumEurMuSf1VHlZADR8
fLc568qv4HKTluSftD/3cr+MufmSI1dwtodxFTFDiufIsj7TMOfb4CnuwIaezzRCccNRJJq6U+Gk
vEuiooBUAkucbSdzKSypgBBr7fveUNmDgG8vywA3eaFZRkzl+KohsjKxFLLplo0/J4RhEFFJY4Q1
NxBeC+ywANttB/0TvdQKw2qsFCrlYDgmjd0jJ4nY18mlZ78Z26h26/bsZ5Zc6ERhNIVYS0s3tmn4
6ygCd4h0aAFnHa1vxYTebmiWuD4cz/7B8kGBM1DE2OdXAn3nLvbFG6STEymFDW/dMGtkib7zzbXV
YE489V2W6KW5qknGQSjKqJRw0NS4h6/ULMK7baB71NS0rL4xacjM5Q1jMkma7VOkVTGIKPwBEKil
LsbKA6g3462OiknfUcC2anfJC+Xrl0cIxPqZp9R478pJ4gSRzX3OIv7eMOrcmefUv7r08p5AdIEw
FlthBhCOsoOcbt9TXc7kZwMzCqJH62uOfvDjZw9O0Raaw46PkSu3eCxzKMId4LghayehrTomTNNj
NT+9h9InWnVuc82NWSS9QljDKUbSTdrutIEFLvocEvB5aMG6SKJdLmm3cdRPaVc20eNwtFPNoSDy
pcpLv60ioZlQn88BruZdZoQVSo5OQiNQj+BnEim8eDxAlw+52jNfJdapLE9FqcqdmcKNHuYXbaqf
je8q6Hl4TF++qR9bVbOnEqZEmEa90Ctfz9ZZ951GrmcflhhtHNQJgII9Pd7ayw+HU3B1cy5Ev7wK
tDquzffj5l2m4DRCQ9p40o1WAaP9NH7pQw3z8yQCR+xj6IE7BXYk6GsG6KYRgE3B2a3C3pBdi3cF
zTduhyXP9uiJcH0aAH99vzXhxDW3JcWliWOXneyYWBmrGzVm6TSz+sb51uaphheXcdK5iLAZWcGh
Ce4vuXpSVqVbBFdmrWhfrOF2F0dqZ3qdUVx8wdPhxBjDzbLjVXW0wuEQHnzdntk7uSd2oXtitaDC
Vm/VHE+pftngEsyKla1jbhfgpxWGZSTgj7Q47ob6mNSieTBRVbsnzl85dncKXjLi+QsjS/lG8mop
7bCWg8/LfwD8KnszYF23PilLT5nOsuZxjBPVX2rwSeJTE3hxPypYllF9/Na5Xt528YRtGSdTXCkz
h4egB6S/sbgCsWyuTzuKe3aSQeMNMP4hancez3HiS4dCZgRSdD9KO6yx4oakiZ4WWGKM8dIMB6CL
FxxEdOhj6WdGeIjNvKlCZkAGS+C4Mhb5D5SuEGsws5zjXDU7Pf6TqH0PqHYuASowQbJ/uh5LWI0M
zXiXnap36SxO8Vhzo7PwHAMgptIEVfoo3yyr9wo1sNCPRqiN8Y8fnupxZ2jOwvu9C25kPZg8BKbd
wkG91OUCdqwqatqQhgTWfMriyM2hXSu0FmKS1CLDALfxCJd5wHhziyVmyK9NPjHqqJ0uddDznJ/2
i0HHo3Wfkg3WtHqEkwRXyn1976JonVCH4F4GvwSf+LgjaeUtD0+22XGaa6U/BIvgraSIOGtcs+Pz
NsP7E38rTzoOVbygBUekRNhNEV8NnV5OOCZuT6FSOFF8wbAdoxCAAOeeVu1k9Nuqi4tH25XO63Vh
N6aM7liLl4S1MByrfJvGZu9lajrW+z0Ae9djS/FxxaSeGIPfLBcpX5DaaoTp8AHXWDmSvLdRTySE
Sp/1iGKQpHsHxOae24wsPPb1C23leYKmoUSx1DNZOOHhwAMaKhZqHwRAyiflZXTwHlwrHbVuQ0gK
Mymr2F5pbxE1hESFPXvS7eayogea1H8xQerIaN/F2EY7SU1IGhsrjfbfkNOIr8ybZZStDFSbfsah
cocKAfhVeXzp3MtcNt1Mqb0qOnfekrQ3RN2w87mOMrU0DS+XgF7i7gPohiiR44aR6y1cHr1b1NPo
5+4jNK+6k1DX7VL/cWpxke2oD4vTnfq6fa82h6lfD2HcPwr51I+fN6TNi6344X7BOL6459wtHOxJ
dn/UZB00L/EqcBXSxySNGmBi8elfzxD6GDgAM/RsrAPHIwa4W+C5RVUw20hi66ljg04a1nlUbc+Y
LJjcLdSgUho3bcoeOFkBaeNrcW3v5QragynctFYuZTKi6GWyzR3VJkBFSJ4v8OoH238zaukZwYOZ
HUUaAZMBCFPTY8fmg/cz1rExpri4JvWqppRNCzkr9c16y5OdgR2kNTBQA7QylWniSYP0dht+SwLu
8dTjMX9QHBEOllBBc8uPeG4GtrozirD85PdBamL3F4aSgaCaHbAJjioZxEXFMzOQo72rTgYpamcT
ukYPsCfb9XUVeD9A9f8J6xr2GTcrrHobwfL0XtherKsl/UsSow6b4XWPE8uXr2SWnBHg1VnAIt6b
omG5+J5cCvZRZ4xxjYpKGYx9X5kYXiy0UHNlGuK9qCqzseu1H8rlMFPSj60e8OYNJmT33zuPDD7P
XsBlF5xcVnYuEROcxy5dHRkUbL2No5oT7ulpwK9FRwJ1fI1ssRtBwuvFqT5Jraz6JVbyNPtBByOr
GTG0/tYD3sFYYQ4luopsW40k2wX/ZW9JAqQbslCdZnn6kUGji0P1a5O9RlBDSNbZos029trTDycC
NUn99JnEVepHY8Zrxr03vCc3T8xQtd982/OHHpaxOWWAynGf76o9z70G1atPgm28f3eFQuY6fyuu
lkQTV2RPqi7r6r7ZURBxRUVUAEnvIxGHSqwQkWH7s5zkCQu/1WsHK3WMf7sbd3LO9HVaClcHGcRU
htqpwCNbci97Y2gRnKLPmaHlS5SxApElV0EDEHZpckfh1wWQR6bJhC8zD+mJal8e1SaKn1h3Olkh
925csq+zSLh+qmGEoni5b3cFtp0d1vwPJrS7TWUCVmIJMxIk9wcNr9DcRutalPejzGIs2EUNaMOw
4yINpbTQOvMwNu6/u5eed7bWxRdiYBjH1sK4hTI8YOQGcbc0OIpO95ttUNz87Gkh+8F7E1C8D6VI
YL0bCcm2B7/soWLEDbeWtcKQGPUOZFg98fDQOXmwn+qSR8YHUSnsDrc1dZicsUtLhsWaiPtrLqxh
frYMIzMRjw4yeN3iw7G/rg8M7lGNXPc7OwjSiL7qWK7A/CdJHXQ3ZzHpsWeb/w3E5csGSunKkvhM
LygqtWkkTMs1/91AEMzCBRWcd2rxJqjUFCSBIGDsrzgJF30UZ04k0Zm3K6+8pOJdCcNlovqSj2gJ
71gr4Ia6kpfy8RG8//TNGexQ0z3tkVSYRkkql+fI/G4l3IbZIKNX5367kLFZRWBaOFOkgZIPFqLS
UjKxcuz6SXUOr9oIDP4SxMVy0jE1UX1yDHTY09iB3YrC53vLCyIP4gJE4gCfI2AlFziXODZMHIZF
B3/OIruAovjZokDJrkGbqEZ/o8RZ9ahKlssXlNsWLgFEb5py6Ho/mF/v50O8zNLdphmepChOiR7P
ntAoB69pwWCiNt8oNp90SXfs+O5xBE9MqHHhzn/VCn0Fc3omcu12XwIgS3olEfyzAr1rtSXli/Nl
bgYvZc+q+PE4o2BZ2obcnKSgJVNMM4y95ckyrv+UlqgGMMioHX+qGbvmmKW6wMm98Y4q+aXf986S
ZYl32AHMFFhC7JGe/iMiNt0/070X9xM6GqKVllsAHNJn07XyeD3SF12tkAsCBcn9TUQQMXAcadzZ
qbH+ywOuGlbEe7dTjl2zeSFrUZmi2tJwbtfYi3K4wOaT1t9QKhP4YigivVV5Ba2fy760DRti22tL
P5HNv/pa25Az3+YOR2q/uAbgi5SpbLz/jiFInRUsAoL/XbkJ6nZAprkSQfuA4ktFvqNlS5qWpdCH
jEbWLmeI6CSDHMCIYPfIjMekRoaEhNcsQIltvM3Yp0w7x2EkFzyKZAAvMhUUMW3yhhKpYArrsXTL
tbMI4COmBrurglp8oAyNwsjvtMDilETB6vkeFwvOPDJaWmrMxLJIZVQsK55puBpiWaek6CRcjHzC
A2+tcqVQBK3JSIY+PR6voDxhank2W6e2IxXemmv4dtmMZpaSosO5ZmFKpfu00dfrU1OnFyL1qKEy
KLt8im3f0NYZsLweip2qYQLokWNT8k3vLQV70saTM0AygM0sW8J/CrY1h8kMmWZpE0NfVi96W/1H
RA2Kx60mHwlY10jDAslSkq3A8bNIRajvXPPW8W5rvXcFmj5vJ/C66/atjyuhIZsP6fBWAdtuzxoZ
Jt7cg8rx6bkA6otgi2gQzligRx6sgyqraxqrcD6J/fbA0wnci8d9x3pd59qrGgf3XJANOv/YhOrL
3y7/R3KAKhIMkVroMJBdauOhOdbodaHhGY3h1L5ztI1gFT5jVzB50kLMp+Hvpjw0IvTmAWVu7NLr
sQ5eNN9hLCzlCDDLMcj0PVHgQudukRb6mMzeS2m+DpEAmd3T0pIM7/3dN7APaaXgb637BYW9h+7W
k63qwrbsI9lcykEE1fpnFA7lVwX64b6QQlK2zGBOM25H9e8C7CC9h4J8IdYDohkZou9CANt2ohcq
dxCtBU+59t62sxvSyTJvYT7ABFCUCWfcU/FMPYXkPRMTtcVPbk5NLmomwbu4L2YiLHrbJwVFTGqL
0Da0TUsq/6zOGc/XfqlLA04zl+aOIaGKn0uOzaPgtajwK304QJdkE2s8FjwYhDR81qhDlMSAEMXI
a7o80IHdtZ5G6cXIPvd9bKZlUlegqPIHljwAm8gmt5hJ5qsB/KRvpIuKy4lWOutc+WpLHWx5hKji
+cx19ls9g9y9Ijdlfr9BCU3j5h05hMjZH9EntpxMeHPBqDGSYgKaLFbMSVAQYjMZrOsVTfLq5QRX
PIMy5bFTtrSAfpBh8S1DGtEXj9z8KBtp0cDc/FRQgVVPKcx/ycM+U/uGHoVBNLmJWFa8rgjaj+ro
Ji+zVmq0X5RFQm9dvp3wryLTj1Ur4dnJA1jBgodiwCExRGu+d33ZF91l4CNobevsn+ZwZqxtT1Lm
Y/JmEBLiVRgcwmn+Gkj/CjxwpPs1QwLwKw74/L8oAxAHqajzSMHDrMU+99lZQCg6eYsTj8HWJpCo
CW+Se1bZdQ9Hc8mpZ7YXx4xJ+m4XhvB2cn+2wlbsa8PHFpXRv96+LbYEQ8Rwa7rUkPOgV8fV7TdB
xrU7Oh4R3/CODN3uCD37bDr37BCY572rHBrt+x0COxWAbCcetEHNS1xv1GXVnPsoyiZ6Ghb6U7BF
7eay1Dbfoq7JSDsng3GpP0oUeCZgMCXTBEHEm5E+5C4uWV/6hLsr+rp77j47/mmyYn2xcF4FRiC7
IeYgJNriMQFsufveawPL6K4n3fRLEvfkgLxI5tziswLFMQP5sgFrL8Y2GyYxN+LzyHjtLD8r7Wfo
Zfx1Bt46+FvpKqOsnlnjT8629Mo9/NGGZ7za7Cri1xwqmPpTOeegfRzcbeBiMbx/5tT6OCelONnu
ViX2o+NxVFir6Ks35pkpaNqjSozJCBCIcYp/vq/CxvbPqvDO1YBxzCmjOFqa9FyxEsPuMNu8d4sm
qBlj34JWH7qAXO4snUqD4Li5wZo2nhDgZpxSCKjMqPUcdcmqpk+6CzpdABJV6515O6gx1bu7MiPJ
RYYfEFJzu9pfArGs3FB+uwR6uqNWDV1/m0oAJA12lkGZPAG4/9Xcn0qLizT15d1u+ORtQBaUUfhy
Zq3zTF9XzO1+ghDy3MfxdbRt0whNBrMoO85i8KHysupyZiW17p4Iuwa4j7/ioa8IJmNSBqwEa2CS
ATZ57KkYz0Q49CSIj9Sx4Ih+VorIdP5LfK/8oOmlxBvF79Smrk3NnOOjPhTTsy+tL+pyYUyHprlQ
5MkQ0MnPXvt0X+h/LcGIeFf8WjlNH5fJN9B0xNUpp56Aqg/hznCLe6u7jjXrhW78528B5We98KON
ZC2nxcCiUxlLjzVtAuPZbYTuH8at4kM7t/p2m4/uFe2SlRicjK1EVUAjHE+mBvJPNnF5u9Vqnqql
Nbc847q/sRxPWAirSmdLLZdnXgofjiR5V5dy6pkEgdDO0uFzxLauKrurbNbYT7aNYYaDsEfNrx5j
9wjUfK3MuORVKNA/NHXjKljWFL012QquzwqDmVCxwPQBmT1X1yqKy5gck7Bj/U+HtqowR2Uvehe+
xyiNgNrngkd/ejsFxeXwn7GL5hKizkv5TLSHmr/btYbD29mRN8cN8EovYcarFt07rgvMhl+6Go3h
+bjzQvoW3FVwFU4fJ0NfdfihNosSHu3qxHgcgz1S1M6JgFX9kXJgvorQlI1y5g9shEpOvOeCOMO/
CEBSEraS4h4AXDWBuAWN1boxjEKbpmAGadd9UplV+E7yMMqweaOYVFki5zvza3+9z22YSjQab1//
KZyl5BcFWjijh2BlOuKxs4BZV809MeRtXe5bJPTK2nuhBcrwk8MmbjdHdZ031Ipe++wg2bKU9YzE
AYLfGR6g5BdmJd/zk6ZKvJj/n3Zr+cezvLohKDMV9k2Yew6DAIB8QDVVRyMd/UIhB0i8u2DwfofY
AlO/stFe4cwIPXUM7rETRe/qwDhWQweCmF5cyqrFqaBs8tHTDweIZQKSA+NAHR3CXD3lPIA3unSV
5V1zzV/+YkOdlZJWzix1nqfLJzzMLGLGeRXMnb0rI1IwtopUZ7GNe5hiZ7Zk0W6wWMOEt6i0fdCa
KVls/qKA9tT/ttB/8FwMPBeXNfBprOQ2cFmgPIT1Sga7yZ+5BJeJMWu+S5rtWXdXYWivbvepRnWr
GdAeW6kzD20Ri7g+44643GSGsgp699dzG3AmE8J/hU6WMqxDjkUoKe1MCdSfQ976i1m71SyIkMoq
xv2wdLMQBKUfb4mGknntGPvlAYHgM82vaqiaAXXKooXvqHJlCQY0k1w9p+1wm/ErbNabiW/57s/y
OfsGGDz5inGRY+wZYotaggsIHJhLwsnAg1b7vFivkIQMxjURtS7rt/JW1+DwFYcejv3kYnDJbnkr
89IpMuzijTxlmeqmEegkXQvu8ma8WUXd61FMYA+u4MjHsDzsEElAHLhyplz/YUCYnfkmx9h7wxSR
RoQJDH+GE0/CqIWyaniYxEWE3VJ9Pk68AJI2igT3QhemvfY7GQu+qA5Jibjo6WHejahLVD6UrwG5
CEdAYCjA+86FTJFFiAlyFmBt3spOjb7cZgCvSgkKPtXhUkUmwvqAvci5AurKz/2kujjhcHOCKYzz
IcoeX8RbDiXeVostKhgpS0PSbCXGACkFhPu5LnrhV/lMKtnI6ZCBJ7ssPzPTtt9Nl24H9YFHtG97
mxo4mwH0Xkeu951YxIIrAs8zojSMAjHIpfrj9zTJmV6L2tanVXmv6X/bNtIejFQ0mxITCUupuTe/
klrgpHbx6Foe6fOSXnWoWp4oXBs9UnI+HvttH76ThKmFcMvJ83ACQkj+GRl3na4LzazH0zX7cQ6A
UEqA7hIfayQ4LRRQvOsEMRLL+rT3B9b6cGtVqLfiFhdXwd+SYeQ35fazsz+61Nqo+6snVTXUkDYn
mN+ZI732JY71cqgoe5kDwGxYlNTP6LqSBrwm7GxXQnxHKM49VgO3e1VuvmgRmoHuLl/Rc69KeA+g
TiH80E4UHoWCf52Uu/nE9BxejAYxvZKQsK/ERyCXc5xec0eZblaWHp3//wEo0+xuikdzue39+3RY
K8UcoO393eTLor2q9mrrVEgTNq6z+ZT+ESjtlWt0nqN2zE86mZW/VYEEfytyEwXio+ErAeKZENYK
q/htDMF3tQk4mRs5cZV5aVnrpDYBr2JyCquOYW6m+kLMWFgt/QUjXv11vtLQk4O1D5vIVPfYsdG2
TnYh+LPTQ0zPRKAbOpbEs4KIddc0kZdDZUqlF+7S+ZnEGQ/FLMURlGVjVbvT4HQOnVGeHtZUJHrJ
rlWFlyTIezBERMLCPXipYwq8BIQyw1qcdTu/QqqGLjyYZ8kE1YoA6jo56sLNpf8IK42srn8nnhKC
fG1GyBeWCdEQ+Mlp5catv/dIVIdsf2Ok5lK6wTLcCL6CnQGuiMntHxT/Qbk+1o038Ky3QW+WVgcp
Ksd6/xDiwMcQQ7lnpdf7hOlJkeSL6pvp9ZqdwX161SMEE1O/Y+ATXcpAc6IuhJ2N8mWxT/gbiSDV
IhWiSQyzYpOh53IpgrOD9ZG3l+E9AGvNH1JFMtb4fMznSymHMRRTEg1HfxHbx2q96XqCF3kC9MVD
Wq8K1i+MN4QJjE2emtuyZWysFZsXVctrZkXh1Y+9ozKtNFwPxyv9ERz/2itOCOxLn0iA+SPtbcEu
5k/VjpIEcpJSOICNY5fGBK4YQQ9X9DbxGF+7GuKeWF8WIrPmnB2SrdXyJq6U//bH+vwXOxcSdWlR
OY0z2yby5gZGhN1eEcR/QPVt/WsyGWG0kwvMkeTj/BB9eA6AzaG53bHaCl+fT77D0yj/+hAPZeiZ
9CPKPZ4v6xYXE35YOzg76+i8BtSliHTce18JSb8fnz8Qr0PfJHOncw0Jh0SVwkZNE8xI/LS6t392
U2apaWDcH0x9oSeuU84hF2vZm49hpmcKoJuOE4LQkWfeGAaKyAaClrn5IBhZX4FJi4RHLtqKJFcZ
z34H29I2VnuxsbX6lwLK0IRtKN7GQ1ay1RM43NiLUyST1M/DPkb8mtHAvfHCpZJaJ1eJUdyfqlKv
j+VoVqWw+pEVqZZMG7R3BSuLGt3/kREfNUotGPXUz4txn+pMbtA2/Fb0rHXbTWbAZgDMikTacEDW
BmDwYb5+MNG9oQcdP4ayws0Ndq0mHPxs/XsLFPkEwSifaAPL0LWLHgQzhggDVZ5nawjvUXUTUIvS
e1fkuteuPBByQaERpInlyLkzRaLrFMXeURbnpkFvKp7Fc8xeHVS87D1Xv/pKSyuVSpuhaL8xPnI9
ERNHGQLIS7m9l5/OH9ypUg8WpVBtjALABcaPAQQU8pQM+Ku5OlJz5MW6jzUycS1flUlA97MEmmu7
MlON1q4wwrFJMOP5PD4RD1rNBx8oMqi1NmdCiaAbTQMz9/2bb0E/FeIk0OiaX5HFmC+WNuGdjGkt
xLZnoSH5Y05qiqPd6Qb7fh3yHJUBnNGouyhqGkS1rN+iQH5oicm7vX0VVJ2mGvBSpem8KYXt5Y6Y
pi2HO4HrTYA0mkDXFEs3nrKPsX4MXh6I5CMcfgCHrpLesw+6v7MnLYqcucrZRxb2JkpkvZMlOPoL
KkohuhMHLvx7YDLOnVgDU7eHqNS1GedhNGz8hyUu3J/nU+ecosI8zhO6gFRgmDO2LvBVXVT52ft2
9tD+xkHAjPMBDzwI2AiFrZwrAAJX1OIOKbrEr75U/GbFxQ1JDRRgH8gP7KtzUXg8hsAW5CHCtU2u
SUzmFhYgM2ZTwuNigGs3SzDM3geDMSmowsNXIrrC036Gc4mv0an6rQd8AQb7vmjfbdL2qefkLyaK
woGeAjtxvDmN6KwWfd2WMoXjVbGkZXORfUpY1E4Q71WmOMXXKlSv51TcZ4KS+NtgVLw8xMDUPhFl
x/D5zfzdoMQHR7s2nz+ZFf1GwNNTSfX2EdUMatKHmXtuHfVDXK9sjU7UKk3rYMkZmS9rpkqZnX3N
6/7ySgXm2b3H0kq7qUjUkco6iQCaXkRbNj5rwLISjXJpbf7/itUdMKc6cBVFzm+K9LdHGSf3pIAv
Gy6TmoV5+RNmq0ga26vBG/+1XK3qLhGUBLTHxRK7Z9RBfcKHPZLe2dBOcgYrcI2LecMvOW7hqjt3
X6d82I6UcgEJLa/rfNygcVoJbVY4xaS0Nifa7JBgeevqqjtRiE+8HW+qVlM36jvxFWzgGgly6xqh
xzTX62QAWvBXRV1l8LzWG+hmsEXI9TfsfmhVYRM1RKnHd0rVBqz9s/fFSGgHCFjAXzezwu+Nuk/G
RYRmpCNBjVmhOg9dDp1+niFm5F/EaS2xyd3tc/Ivw2Xq3k8QOWqrD4V+1lzppyggE+VyZggPfwkO
Ti3Fr9QNqUElQmxeyP+XCBMKkFHxKj1fHd54lRuvTUU27GlT6CSbdWYZUYLKioA3Z0bMLRMHsHi4
jID0xk+modXB9I7ZrVi+vtmr0h94mnidNhY+n/igzuugqSm2NIFZ70aFzBNwPoSfQJhVXonH3b4e
9GMXYdajFFq2MT1e0esAIHRraXrEaCWT669UxXLdrkTSpJT52zxD4J8xnDKg2bpWcrMkbCTzhNX7
xkRpmQQ3C/ETHUxsHOgJ8UJLvsWzYC6pvoU2JP7koaX2UMtrzayo+UWNE/RoHeuIetcv3g6ew924
I7zmO8Nb8J3XtFcflRjyycVWUZsKaWvLXs9o94r9i9VoTf4Icb+w55o5nLkAHSyhEE1Mbnrc7n+K
fJOxp7A4XD1eHRjocPouYXNiqURsceoO9s7FsEB1wutjZd5pChhjVkxodJRFrIMyKl+/XBhSXcE4
SBubGLHXq2XC4IcIr3Vcz5PCexgA1r5si2x8D5Es8LFr63K7lo8HyDZRZ8QS6LoYSxqkGHtzi/YR
mf9QFoL+Gsn4fC6bvClxmbDGXpU3sLx4j4SujiL7Lf/2v1oe1wRoU8mCx7qCJgDpVHUI0zeO2xlJ
hXLfckFJzxdUVzdDK1xIRZD56HOxNIrZ1mZtsXd235SXtIeLggZauj6bSwYVT/mgrwScguXtEcln
OZklUnUvyT9dpV6XjmtlnP7Ep6hW7kWD7ZXuTMWH8B8VEPuP/T6AL1UOva/XnezrkH8mfFAjmpO+
hTRJBA+WcTqNxclWZpu/1Xmqcl39xmF9B9ar+YCLZkhx5EaUTcPqoqYPRLBeVfz+lOLyW+yz9xWj
euvOXR4X6Kw7qIEdoQ4nvyhgPG2gdj5vwb8XTXGgNj9J9+1GgFT90OZdUCVL6xSINTZj/NjfTqWj
4XewVnydXkXug00hImAMYbrjGMvcBZf4mheNHe1z1FGemNZdsCUlku3p1uSnKJ5lnDgki8QtQkAQ
DpH8BGz2vfunzeY0/LQsjkKGoytvEdBursmphfHIy51ppRQIasVy/bwKxf5NlE+rBlne7C24u8lP
Rtukt7ENGH/T0dT4z4qMnwFkxQb2eDPoF9ip+MomYQiXGvllA7tLZjeKnvGx2W404Xx9nl1niqNY
GqUegOJqYfRanZzVo6DBaZWQmpXuudB32ZUE2g7uCiSdL+6rFYGk8R6VqkF7TJPRRZftE6slHoAb
k6qeNy4vZPzihDQIiY6V7ZDA7DwdA75rZuFzHpCOdsRARm8HKqpb+eT9+u/KoAl+MlztWih7Ppah
P+FsZWocvnpFaOh2L4CxKrYts+p2tH3KbXfF7isWW+5feLnqC1MICs0lcGFgg5RFQLjktgBlPHti
JwWk/wN59pXzeRPGSpR7mut7YR7Pe9v4qSZA0nOHOha0YAkTz+jgDnJHbatZQPmUgR7Kg6ucu0bf
zQB9lwRnX/gFw0L1DcrsTr8Ygrx9hx5gMlYio7oQ0BgaaNw8XMGt2k9nCrD8jfztb1oMXP+pOde5
FfN2h4kxGTGwfyQlhKOoZlsUPEs8evpi4q44kD6oHtgg/zfr6zPvpNOwFZgiftmDubXdq6omj4ge
/F9l8dpQW0U88yxzJcfMy+l46OOwCrP6jKedO4ovUXW02mazBoyzgkaS8vj0YXiyVJr0/cuAuyqG
fJ911XJJQOvhLwxGY5qLIB8VkfISoYpLpxxm1yuDjzAlOF8tqlhRnNP5C36d2oXCIJT2c3X3+mCQ
U9BVZTcqUqut6TFDzuIZkl/x99Zjozr6UmD2VKxbsJti8sNHkroTrxjBoas+fgRAPtlvZfENYf7q
oaVw43v04FBP0pg7zGaaFDtsaN2aiNew/JoHs/GzFI31SJoNRPHJr1tAwV/R1ePT3LBJNj/N7yb4
hLB+G7JdNX+pvGmjT5iZDImAQoiyaaa9JCXwCHq3JXqpGM+CZu19gXGCce+HDScpsJ92+eefQ91m
CaD5EIVWPqT3q2eyh66vdbDiZi0YdE24e5TbHczdTth9Ho2G95xl9CTsafAO9mqYhHzVp4o5Rf5G
oXGZPdly90v0yrnba/MOJBUb3E7kBCywUqsamkRo2vSKGeMRo09WbbSvY049oB1SbJQ9Gy6Gv5gW
bTuIwcnKxLQlDzKg4VBniYW0iEtBdvYhRiJy2c8W8dYRlj6qWo2CtMHMU6T8wKHp8T7+nxLtCEyv
PmbFkR+F2pP1TpmpdFJI50WwZkXS+gv+buFNckFXQrm5IAsY48grPCqzgUEG1INdZYFmtM1da7x2
KQiVMkXbwSf1ZQDTmKXyVa6bBvI5kLeVhkgh2E1Ks5mx0bz7EtURHSzU8Yu1GTQb3ifVNqOi8XYu
gPrCQxs8+WBr3wgrv5qyRliQKhYOcYi4LiChO7/0olxcTkJii7b1UQWb0N3QwmSOtPqJ3c1ET7BZ
Vj6BdXdS2QtTUYljhzTZTiZoZ39eOLsQz/t0QMJCZRDJJj6Yuo3IYpM75grF7x332UT2ytFaIGIq
WbFlp0D+zSzVkd0ryVf2/7QgoePgrQsj5oY8LUxzcUT7rW67Bs6Fb7W6hYLQa9Ru5ulX+fI4EIHj
fq+/aUnIJ1pX154r42EWf7pqFL0jyoIqQioZqrLQeSNKo9/0ywQYpMeFTbGeDiSHKQupuuCCIXi6
XBsTbr6foBVgoDDSGLtkNCDzzDspm4yt+O9NMyYeYrO3mLdXWhcjHXNNJJqpAx1u5shSeDVui1Ah
Uhw1458Y4/7jzoc6eBNhUvDPxhUt+vEn9IzC9utN+HRIR1iorkyS/9oIEUsntfDuwpD5mQOZeiqO
xk5d+zD1e302PaaMU/KB+lNiHzDziqT/mzLbyg1ecFUiPA2NEgSTQ77ATWfZTOCMmz/npm7sSJ/+
cj7Ryzyxr+7mxEFp0+QCtRU+tTl3lK+feRu7SfZivMz7NvsalKjEEaFAxIh0Ju4ImTp/oE1ftV2/
v0owxZC1bEt02rqdk3hRFW6gnt7tOWampcd+IcFDoM74L7P48pVFOkyIndPrEh8GeAV07wV9p4ew
D9OOi9UjoZn1KXaG2yLzy70EICp3oHgW/Ki29JPNnxoR5KUFWCPvFm5jRSQvStXpTQcWJtryJJxc
u7I6voRkMmqJPyLcxsNC8H3L3Ril6H6wSUBAsLWC9hPa7lAQyFx/tZ021TyRVu1d5XUxsYGeXKbk
DziU5W5bYpfzwNwWoWtbMkqhPScTfsOU8+3GeLGjfwlWPSUCz0RypfBsJCiRqaSAlSd4T4CBZ7Tb
4z6uUcz+bxHjBEhLncAJz+M8EjbjTN3/pbjutMMVpBrG03YLafj0a448TVmwCJB+G9vGI2DrXDlg
GUWPfDehWVo3Stl5sK2XCATy8LxlhioPdSpZkB0Nf5LCwxzHou4zJrIRC3L1t9dQocFHPk8917d4
gvTfujwjvWBesqI2IVGuJBVy0rpgkwO+kzPHFMmnyvdIFi22x1FeZvyqz2FkfBas4kRwXWWSBEJk
D55p5Gm7VXzDniF1v4Y8nUmPu2i8v5yPZ5yOkXymFly0G/SKNjwmCR7OpM+8m0J7SQWFiKADgjm+
rVZ4i4kGfkE/rvtxqAO2EvjFRIclYa85qWSGWfVoLJBahuvRwoQOyCN/8AZXDz7to1JIXsebT+TN
iT0M2+ysiXXmWWpI+2lK7B3kTFCfhWzSLFB9HivJnKHG1N/AzArEt+XD0SCtRkw1YKueIQkClpWv
djgsd+LGyb7Z6xR3Ka0EPd1XeLX3BpFdss/GHnvbVkN5ve8/RW5lz4MvVs7auLqQlFN6XL8i6ekz
KB8hKlq01y0DbqZGnUYfmZ7sOX3ZcUTXhJgouSMq4na7qVIqD/p9KG89sSbaG8wL0tRwnJTIS7FO
its6xh2ACPo1anknKsy54oY1eaCKfOTR5weL2hPPBzywFwoWE7ly5yMuxUIwJvAJyxFK1QIrsgHu
Yd4CiZOv6T0TpZBcT4fSGvLS/y8O2ixnOFB0Y4+ZCPulk3Zz3JmJW7FvMiVjYFtHDxvBWZuAem/K
EJvWy+7WumXkPodMyVP9nC+oqf36oP2Ld1GAtbhNcFisGSUdZcAmwiAhnWWKnWSPN6QnYlHgvejk
ODo/9yjnh9aPsKQD6jYftfNGkLsMgZ6R2CjenwHZE1lJnTLSuZFw9Pofda7Z3Df2GucP4OMDeJnJ
bjo19k8cCkuaFjTlqJ+zhNUEa95vYpct/61C35r1+r9ofecdzdSRpXl1xb+6Sq3ZoY2tsRzGkoo2
PXoOkum+7UTFmAdczH1WboD7iYi4sPhvBbPkZpmtCb9FANDj76vtIetTaABc6NgL6P7bLP98ApN2
1hPpWdvc40TIPOktRDbJ97sKXJdHWWAwDqaMpimEJPzZTu5skXCEDuVHDHIcbAkE1MOSy2Jnezmv
IdTJmSByFaaw79Dcq0lBpwcoVRFeJmMcKQGAr/9+6RD56B5B6s+/ss5YL/aBj7Wd5SDKGMu6W8m6
JSYcqsp2QCAO9r3j4UmaMmkTxyvqJ8vMzqCVSPUPHbRA2KwlpqGnlt9t/WiVDDdd1q2VWqTS22Vj
NjXu2qnXgKhA0E2FZFY6hJ0F+6rbjEQQvlNcJY0oB8VmAHPwXPaCjnpedRJX30W3MeHF1z0uGkEU
gmsS4IDca5iYR1U3IFB+AaDJSery7N5tXDdXfsht2f4eJhLPYZLASm3jCKxOav2UB5eWB9RliNZ7
SrCW/LLZ0cwFDhQW8KMCAk7Lz9ONsLthj/BGxtLq8lO4Sl3UI9yfMULkXtFXSP672e9skU7HJHwe
5aDTJeFaVAtO+WJbU5xJKQ5e0irUJ3VXXyNA9jXxJy+Kcsq9LjNUqhUCbCofdwwL+YB2LdMiJUXj
nkNwrKg2z6PK/QaLmcTBag1RZsD32OsumWniO0EWSISxRLGXfcUVdryJ+zbZ8ieU353xk3/+S1Xs
zWzKFsnIBo9McPvNEJ3Qzo0GSJlrnwbvnzU5/M4MSc1qbrVPrwlYDsSdXoyUFwFSBKUN4+xFpVV4
QAldWC0N6z9ZGoLB+r+9V8uv0E8pXu/GL7zkr/anZdmaSNmPluzO8ZyNnxXwikyz9j86mKdmJTD/
FQBfNliCksnNWMdv97fZmkSNyesbjUkG/M+yFMPTv0BCcK5V3H3bBws1hRPn0YzdQgXmPbwaptA9
mwY3+7w91nL6FPUtoc18v7mmMWL9eKCRV46Lxvge1Ha5qSMGYLXWYaZ0KKecF2Kq8mhaSquc9nQe
9VLicxm2hjxS2VgGLswCq0Ci2XXpxuhRMr54/6aq5jYv38NOj482oInV6FP2AflTNVPUlcKC/Z+B
lctya+mFOZpMKTVGztLr5CY+HLNWvp4sQvWohZUMz2+jqZf/9BsL/2d+sT2VZpSd1UHtV0ZJ0TSz
LPvHay+hB3pZVR1XknLLE3S9dxceWTLHU7XgbPrXK9vPxKyWz16+NXKVvz6iyaWSD0Oe7V6t27BR
vtOEW8WwMk68Ux3BucDaXQxM0KEokMM05UMXQqthR4AVmw/F2STfDsyT/e07yw/MKPY+5BccrGv5
iGC0j/Tz4YE2SKNs8Bj/8tG05ZaBHM2qiLObvMdB1CAl04f9fvmj6Mza6AzLokbyIjiyyDhyD888
+h5/t2xfgLJznlGU33to5S8zCJ0yUIl3legsMU4F53/W4vN/ZLLtWMp/C+l9nNaRYpK/QLmx5p82
n4/HWVlW83ilCKD20jBWrNf6ETazyqpygfAE0579iyYCUEPvdon1K9E1CYrcW1pBV7Dr8k6lPG5n
AYsJ2K7U++dbPhUm66se4rvEqSrjOvYVSVf/LlvJbLH84x+Vg0pZVILYUQ16DFYEOc2wN+VSPT4E
mZmjla1tJ3TI796A7CEiMnYwhbru7Si0Y/7VF/fO337aIdI0O1ol4VhZmp3Ch4jpyNgfRO1dbwx3
O8wM52eRRxyioBeOF/ME2O1gOvZFUEqg7lExFgHdLWM20HDQdTNS71Dsrs4CeemXBE2OHKsWuXmi
H93LQqbMw3KQ639Fl+GULJBHARrZkqQJeXSQaZTKZj5K0nqgiEGf28j95aRTYf7AvAA4XJ8V2x4H
8jnC7JRpQyCJPBx6s70TjgKk7yddUM9PNqy1cvVJWsGslLpvzCZEnDHUuEpseiGfDelT0iWuQvpW
f7nFj85BXxpANxaRePSCl43mQC7VUh4UQp/FUUgTz7atWtSdaW4FTxsxkGklnG4road8cOlE06Uo
zQg+uFsv5o1DwELjYcDzYltUA0ffPR7RCMHpBwoqT6bCR0hTieITg0ELYnYjNL4jdU5Ab0kNmh9T
XgiG/ZpduKOwW97cZnE1/Fp3zTujxVaB8SgK6AyvnlvAy8b3NPXDgT7ZEjlPgRKmKJb2ghBYeLPF
RvptS2r9P2YxVtkdzBwjAFc7NA0vD5e6d6AqRy0hITRQPcnS+QLEiLnVj6T4zmStEbjPrg8xQ5fz
rj1OlKPCom5dvvjIngdtTGDRmak1dF93PlWioYJZ2pTljWJCghlZZLYQTbVo8VLs5GmtCQtgWuy4
LiNz47FmJE6XGkI+UpBf/HafOsoC2U28rf06EkteTPYLAzORO7mcV/UK+1owLxh+Su0Utw2IYSJk
+WAJtV6UpHbprII2fxcrC3J3unEY/9XLLnELcZaVRmfGJQjXlBSTJrD3jjD/DZna67wM5zQNvU6l
+xGe+HvkmgJldsUvEj5Uny0cWmgMXqf3LG5xaKFzKZ7DNfShZl+VwmRXAdtEUSa6dXJFT0INSchS
l0pew12vTfzlYGVjtA9dK44f1fAsz/f/aeMNhpbFRZ8UnRntlpUBQJggo6Ys590jRx5aPz8hSij9
sdAr5/H5y64xMDGK8xHeq65miM6hdXIwNDe7TqZDte5NkeODs47G5lUUN6kTSdoha6W4RzexMF3B
wldQ/Sdrd16vmUBa5cbflZouqycbIBEYUR397G3gc37aoJozHjpVve25M1BtfB+LANuxNyayriA5
cA4z7H65NafPRdIJpEAv3Mt2JM2TFGYpAbbFtmBn62cAAtKgSVSqe5QwjGK9DfdQ+Q+631egrkW/
wKEm7FN3ILiZ2lL5vfCNNzsp5G0d5xbGpHud1iZ/xgonQ7rGFu0rXLNbqSfywNKczQgA/lS2h9jA
2q0Wu3z2fwEl+RvZCXRSesH06aIEwVTamsmpXD1492Bhx/xPYHP0GPa3l2j31yZFdlPc3RajRz47
GIGRhxlbrRibIXQ5eAPxacbaMuVlTygWhiIofOvxhKT1DNWof/cFFmigFbnI7ATTpZ4FNy6jATY0
Jp4X6CUg7qUHOsGl9Io2uEjpPK+TcqC1Rymx+BX97V27w7cNmrjIe+XRwu26ZjAiNoCK6Y5xDzaI
KPB0BX56/tu/H1hEdiPoeJICmoOseF7UWsiKfYsulrSzl4y/JDdQODX1rxF1/wbcvK7DYk7imO47
vJkQkhLG2nHJyNUXXIlrUf0FMhNS4bmO7UiluRmDyWOJHWXYnNjf12SJVHL4RWgaHK3hpuJJ3Iga
myIBsDMxfTApqlajndBxURJM3GhMnc7gt9MXAfe9JwfoJvxSM8BQZDvgi09jF0c1yaGvowtzMPUz
XzOFNBaMzyMXIbqIJiIhy2VCkWNMxapXAZbOBRXcJy7iJ/+zNAvcYY4KdlkvmszaFABiasFIw1hj
Rf9qBcHxJbdNC/eD0XzV4BJLNiP9cvM0tbmhj60bZt4ORqg0td+BwMhmwK5qIFLn3ss9kUiLSP0A
CBkXaLV61390dboxf683U9fBoJzq9m+FBjFid4vEdqS0aNyEM4zShS0950xxomOzukOn8MWpYeez
U8f5w2YpzZlEqouxwRb7LgKduSPrCFH5xrOWOnGvvvR3gBbCMI5uTftxfeli+w425ZoJPvfGfnxl
6Sb3DRX/SQfYYS3SX3VWrQPGuEbtX8lH/Iiwrmd6BP09mCc2QitfosTdAcaFIyf5bHuMIdeg9Lok
wEKg0KPJZOR6ERb+lLdzkiiglVVqm4yMpg84pjcKKzdMlYoioWbZOYCHYPMopf2NVD4lXw9noYJ6
FNQrvHv2Twu6BiFZC0ZcBm59XaKgIQ5OgHuCskA8lbaZMHjtsIaCK8hsUeHyhh6G15bRDkaF8uJm
HtNPCj9yc1FdWuUJlF4ye6sKY+Wr8aTbccOr4ggKe2MD7o9zXUXyQuntXVN7iu4wdK0bHH2sdCKL
QbN1kYGBZknkIUgrY54Ys91Ljh5d8gl2DWQYY+0ru6u29fDFRvo4TL9olsPUAURcVtrLFHFdz1uZ
QR6tyANnJVrr8b+Vqme2o7Oj5BZ0EFeri8+SCX3uMaePTnLel5Om37n/pgH6/w1Hzv3exEIX9xWN
xI+MhhS7VMVe6G53ZiY9MQQbFxqT/MsYVHqQ2uaT5OzZFcVm99Vuq/sux/kZf6uUYn21S45IoEi+
qHgKi19dHzE8Cw5VJaTOdiM09UDtIOWBajZrZXt/F4h82oKOrZ0NrLjBqEMqDU0A3tSPlaJq7Tkb
qO6ZTTbRU+CVXzdoRG6b+8uVlIl8MDxSX8QJ7Y/tn3232mwoo5X5YzKkaCgmRnpu9QCe7eYEy/tt
bPCQbiegsdnMJ9bLyCnbnsmcT6Ax6j4+zwdK9f6t0LWACqcEd/ZCZmrg3wIseTkQOY+eiuhJboVB
4fLBuPCHcIMEbw4zDvniCqbt0wURPUbLyT1Vh5jirykynUmAM/cawsHLkAv7mYUP7N84W5DGSJCm
Qr31tXfe+NWlVTU8ogxTlA9/zIRuu3Me2XKeMTPqMzops8TuXHDDQzh9dj7mJEFpYFSRbJ3tbQho
WCm4xcKqhLNYSI/olhegcqGRl2JZAj1CZDy2+1xzF4isFrSQf0y9uniBNQWmHAWybkXbgXvgQG9V
z9jCF5BI7M7FKF4VcITZdOhk1JRYRWflwUBatK49nv/y73BwkTz63M60Qw/Mplrk1P7InH4WPSmP
QYmpz0/MRwUxLzstatVyMUPRn7Z3xMhYwAhaPyPZ7353enZN8wHBfsYVhtH4otYKkr0o+QBGYAXn
lMrKGaugivZabFIPNUeUi+uCkESaE2jaC21CNQO9l/ivfuUIjjVghuvselE+Fr3Uccu13kJ9fvtG
v9dgaJO5RJqmpEDUDvlMkFAVRJHPVZu/KXtktL/ul3p+l/WdiDfgroBf0YPDJuxTRqfKvi4k0qbU
UU/jxkyZegwPGjav/u36z7iM/nQAVDmISY4U4oFi0bZhtWf3yh/JfeUFGoic9bX3USf0eYUbqswa
p2Drnbvb+Ta1uJH1Wsyg55t1ed0cGgBR+JVriHgNkQsGWbasgRsaf3SGtEtlaWYqppFdARGFln4Q
KUAXeXHRIA1FT2A/q7RZvZzXkl8/IEwsm9Ut4o7OFnOHFArQdgs9+tP0GhSFZAIgtNd9sDaQcGEg
fulDE32U3ktatAZ5XSebMum5tkf7tLue1gY+KtwReMTwTweZi+WuY27mmiToc9lgAuh7+7RUUqWk
jYKjzH24hZ9NDy7xI13Rq1XrpVEldJPLmPAejwOl2bsvG5H6MUUQFkMO0e/orHxQf9Ekwnct1KwB
Uvgb06RO0XhVDSMqzUoetUO8hKKjtScR30krrLeRM/IjmL1XEXgHr57tz7pILCaxEqRJq7pVDD+q
Z7bOHr9WR1TZOHy4KkPdH9x6ce6p8GfP2wFibbJ3VAeyoWOxAWvROgKN901Iu4aX7CMqhyP6Zzoe
/AHjVAjBUZi/z8WFBhoNdEEzIPe5HA71tBT4jTtdyYjxAj4TzbRqNm5pw4x5mZhMqNnvBxVb53Uk
WfdL1RwCSGZqRC7oN7lj5/Tp9ch4KZ8qlNEfQMaevHhTBAlBlx5mVauPNBAj4BjNjYAnt+3HBgVW
w4miMWbXuSU/remVA93C82yanb3x7Ro8v86nyPfQO9ymVWvJGvwXtCuGIRe9DJ2DRpOxwiMk9jJ3
XHBoRb/nAs93C2abM4HdpPslMkA9/gDZ7sfEZ7XqYGM9CNnP+LuUg5gsRRDA69G0/xDv/KU3kR0D
DaqSD2c8FuOJdcz9DNHHib3SPnKp5+L1yhSRSih6/E5GZ3LWygxpydXEAoAnwZKrGpegusGVfNIC
p9Saap8M//62Gcrwnvyco3gSEvsD+szcN0R1ak4PgIjSIw4vQfbQAZUtokem6kUYsTuqkVxaPpMz
GyvApu0c1Tc/4h4aTLyxH/IRFsR4KUWgBib6RCEldGWk7FctP6p/qE0C8ghGaJ6RIvWvZGSuOBQz
rY3+oS6Shxb/eZ7E8aRUkALOv6gH6MQz/U6cvtJ+7vWZEq8BROUr4HU3oJPWfZpT6DmBwUYV+78B
lIKRJ4SFrcDY8su9pd73fP/z9aVYkBLFzTe3e+4FkUGsMdOLVPZqFNCjpfY70+HuJCfUfc0I5a5s
A0afHTVjyS9/8u+KExqfnGATt4oe90bfnXBG/3WOGVlNwjlW0xdxHGO2pRS52jTNCue9bz2QQERW
6KgOAWJr9iID/LcndnJn1QeW0bAIJpjEHolvssdE2RijKRPnZ6wQGMCA9OJuOuIO29akQkaEKHpK
tQTUU3LVx7F7qW3I71fAizf9lSoUq/OSbaWcsGDrEtgsutCeb9zWOywQ67AShBuuvmBjHMNmp22r
MTk7VnLH1OLGek1BRTMHK+QmUsXpJBQpBuup1jgKMe9AhL60aY5B/SUAI8mWTj9q04ynDizPCX0s
Axx/+vfioL4Al6fWsKzZ3pkdCdBUEyGr2rDckCKSM9aTRyneAqAkvhQjpC0UWP8dAlcx5kg6Un6c
DLdB9nn0Qo75SNt08/b0FLnnCqPbeZn3bhH/VpUUOS+GyjX3XjuwReN0UJ2DzqHEzyi+jXZo+sCC
BquCbmyViCdUnKN5qQrID3hwa+YFM36BVbPdxByilJgdLlBn/mLeWtLhlAXHWYBvkpdkDeT/Hq+m
bKmcG8opbQe80ECAziurhOzsIGBcL5NPnBYjwcwUsvVfZtFp+kez/NzutKPCpKq65fX1SMoS+cyU
tIkawMQz9F500SXOyT0JmKXSsYKDwyxVzojJJP4866i1xuglbqmBrJe0SA4tkIIRrjCpkkFtLsOi
qS9lrhHHVpEnM7yrYz8Ifi8VaQwufaquzLmBqDxwEaDx8zUv89vnK2L9svJNSfQ1PV5p5BCVAUlv
ouZ49LoDRzypnzf6e1y03JcqsH6d+1wkXANs/ORBnK+MJvjtktZK2WIVVXPIeJACQWHPFtrhyEVE
sPmoVo3s8XmhX024/9dnZZWHKgPv/bm170VMQl7m4dPjU0IqoW1PYulVeoISgPZdnIUFgMtZnecS
RFyKO6ShQbkJz4WbFRQ6Pf+BP6grWk4NIR/FtYesi1GuV7Km02py11TxGWWpB1blaVDXpAtygknv
T75a670gWPD7BdXBGh5SEvbUfyECCGfFeiwot9qp3+Ej9dYcVLKlAO0RTzevbALa9ym8NMp7/nQR
c5TYuKSvkC3/VkSSv7DKRMWL2pL6gu93DyUZB4vYpvp4UIGVITf6MlMu8p5fqouydV12+XpN2nOX
wOXSk9heDen+Gw5kcGuKfJgT1Ba5dfCJWhAtex9NAToTKJxBe7MHDaB85GfVkB/rsS6F3Lh40wnP
XJr1ovsEOOnyTiyKvr8E8qXlp3UIRJciTvj33Sv9+3HFBj9YIE8lFWDbw+uawwxbeeSZInm4eIZo
J1p8ejkWbeugdeQyG4Hjn6LwSw4oVe0xrxaBx6ash6S/IOVRA0muB9R1HabUFsz30bFRDcAjgQ+E
/xIo4AM7gKB+rZouKuRHqPCXbkwmMqPSfSWltfMM00L6L5XB7WaZyRP3xlv3Mj5VVKjuFJjwq30R
KzuzP8YDrFqAPOaILANUUwXXFN5ZaDJmbFHJqHJyfQj0IHuiil5IJBXDKq+cbMZV/aKqkw7fJAz2
pcRSI46EeyfrZLOpZZxpL3DSs79MKE4JxNUj1KfimHViG+62/pCtI8qiGByZoP0frwVwlljSu2BY
HMlBHyGN1Jde0YlDSVX9pYQu1RlhOoSEpQR7o36PDIi9E6asRkW41CkH/a2o7RuDCpqhKZRAZA35
sgrHnTGzKwYFnfdn1UeQVav3X4h7w7D2D0rdah5O1xqjCDSnk8l8hVXCeXfk5Oxr36bLfUPp22Xe
SpfXjNxcWYjlS08ckvrEfSnxQrv+8n7txdAi38I+JZDoDHmnsVEh0orLvO/370m5+yLUFjRkP52q
ifRD/Q7JjoMlXfwxgdh7+8TWIWA3ML7JtdQ9sYQMh8M4pVsqr6VbORxK7iiPQbSWjnj1/nyt93eL
f5QcAzr+67QPubPADxKPDNM+Akr/WwUrdQd4EiTiydCGg43uxMm5PiM0CKLn7BGpf0Bqf+Jzf52l
YgM+XYvn8GLhiTlqF4ZTla+mVsHjVc4uFCraxUS+OoakQ9WMDvAZ6kseatwvgWBtj60v/E6sb7A2
uiuYHlT3JQiTNsu8u5zjR/jhjs7aZLmsVTU7oAoMxALKJiB7tTZvD43+7bAMwuO8N0d58XrdeNq0
uVaVHGaKg+GxrdkwxY4W+Z+QAtS9PJPNfsTCPjRp0fWPpXcEOH68E74+ioEWWsps2eHvDDeLszsd
AuEYTtK0rt4kSsUm3aOrEWDDNi/QC5pAOJjcNkSYA+k+n41gWl4UrYbXjBDDb687DissnjKuQjUE
/4iFFa2EmPLoHViJjzS664vlhoDe47kii5oHHy+ROz9nqoGmgSIrdfxXlooqy8P0t+E0Zs9KEI8D
y1r/JNKQCQVHxxZbEy/mIYTrLIUnIPU7FyWGabbpqRllSf+KAtCB+4vwXlJ4iUKcLmCk/Y+qnyrZ
z1KSK9uLVeeIOY7gz7tn4whQ8UnZ/8AEI2T78J9mMa0E1tjEuQjQzQiSBrOVpRjOTmOlK1ddOsAU
HcR3aFZgjvUAagWquLy2aVDb+TFe/4Tidnl1pif/JV3Cuz++z6L/+yu8MKf3yrYjul8Bh5RLikJq
rF6d/SZdavmZ2rU4pFP2jDMS6GoFv/BEck8WPIw77rh3grypBEb4AbfmlL1IP2Mu06+CQUJul6Jh
22gtYMAxg1o0709z9qudbIIU1tsaQwWiW2Fr6kiHrzX45ML3LYlcQ/6RuqitR/wTcE0YksAFCaZV
67b+3Za+BVP6X0BAMmxZAqKk6hIfzATEVYAsc6EyAPXO/BPXUfBP1nntzVqBDkLTcUftiaPHln+F
UKrC9sHS9oOgfPZLpnicAv3hGryp3uE3iIMA4E7/1sREQKD+T/tIHiA6ydghN/D86Sq3OjU8Q5l4
TUHR4RnYXJCavWb/2T67sCH3Ynw5KTLV7WgVvWKT/A6gYfBKsRjK0Eqni4URW3utdqEL1YcvbCdX
7Wsuwz1OF8OdftEL4BJU36jmKIvIMvktJ8wwNHRa5nCefqGKGNxzXT19FEjZO5ajLfsmMwKFUtkP
vLZuDOTYFOw10WKVdnRCMgWdpVOYujzai5VnNVIRpFmuah8KOzdgoQMtbWepZSQluUZ+wbx2qMZ6
dsGwRX3YSZUs+BmiCAqfAyYHJ8ib90v+JIbuHAZup/FoXq10FTZ6BbHp5JGw3BvjyYNKFhl8YHIt
rYLdvoqtDF/bHiafnPValSzUZNMatzCGXRDsy7AeaG6Lgz0nVhkyt/mrggNDvp3PiPClgHX+RfeY
xi/CpcX6Lo7L0R/Rvwuo/RHM3yDOKCNsheaIzMVcGgQycJU/AmXoDS0GNgEc0QGuNToka4sZjHLU
MZqPw1mqRClqDe1fmxNbPwzObucOj4peL73k/t+1JfXlzDfXpt/SfrdhrYR1mKMkYunAmOxq6SgJ
rw3WsBMmRYNtRJBHcCsFYqNn70NM9h4dSLIwyw2iFI6TeY37Fu8/X+V70ZxG10wsmCjRa8QzzoWq
qmw2d+SdZ7kQoiIil/UIthyrloh8nbIauvGhIOCeCLTId7eFX6++rkSJ+E+PIvBJRWjbTHynCblU
XYd/gM0kmOiNatpaE/dFStUfnC62dOvTusrCaoKvbiC9NSirC8J/zwTul0cMuttqb/V+1L2XumcV
3LUy8DGlgFhAcLNMmdHzdeUO/fageZ7qyGFSRIMcoAB3tojtw5fsP52oNGPc3kPchNV+ZEWMNbNt
7O3yaRECGcRFGlHVYy1jZBcxXWA0UUibDipeT4W1sFasU7Vy6bzhr0skMA6aBNDuvEMIfoGive3k
gy2mqyMYTOKiX8E9v0QgQFezOgq9ODmdcyFfq2A/0bH46Y6/G1IWS9u50bYroGHsHY4OMZl2XHLi
Uu7YoZGuKnQWRf9cJ/rZU8tdX3AxReRUprbpIOiOROiN2UdjoBsTm3Q4os5/uQY+8wMaPMfKxeW8
0qTcSTh3BDYsIqjobI17TfshX2gbSQmKyMJQh3CD84R1hEPE5MB9JZM9Mdeo9llj52gD2cmFI66B
vUpE2kVJTBG3VZRPmMew0QITbGPaUJI0+ntlrli6Vj09+HNl6yoGpltAK0iPPvY3huIIO+2foPH0
P3t4ZZCDtyE5zWdo5uTmKBf2Q20nkyVfux78tu41ptWzkjMSgKhBY90uVocymXCJIbGHNJN+LPHu
wtWxFBFiJCAQvCYGJGnONgz9sF0S36yoTLEysc1fKsJoDyUB/ER/vBKrYMIcNCz+TN/BQVAuAHgB
nenAR/OZ9RUhekc9G0tehiCvLgzmf97rdN7x8kD7TnwpQpn6cqP9qVe2uXRUL/G8f5WsEQK1YMnt
mtZn9zAtCJ8vXpgH8/itsJVNKW0tZIlkWquvJxsIQVcsjjBCCFSc767y5HIztBaHHST4rHSIpOiJ
pv5+gtf0tNqkHDbl2uYiuLgit8leV8e2jkMFoxHYay/Oar++BpFzEGrvhNqNtvc6Zp7etlD3FVRY
jU4xrYccNnQ0XUHxjDgVkfq+TAnFQGCQNL3euG7kg+dsR39l5vCVqHTEVOn1sFEjNl7TKptE5sxO
XLMtYFtzcER/gnT8dVhFSKl4HHXyC5o6CPZyGmq5UkUVjN7cweXk5WwofENBlfPfR37wOD0L28nk
NHzPEBsQN1QK9ZfJ8hDABGS0e/mSqhuNfG2+i7sVCDedgdzjo4dvpysxlbT7IuCQI+FqzXhmBU70
FYN/RkIGRUGvsW+rP1Ffx9rHXvGalzBihWZXHziwQhASJDbUfoP5rFu9bWveAPBA/qwdtXcA0YNu
qYDfPyYDCXWmG4Z1+lwr6kP5zBxi77QWD3dsdwId7qnCJ1vYiv9Si6/J7hz9Etejff74AYH5A6oW
nWbyDU0CHSr83PI2paedhJQEu3fmpBkX6O7KTtzqMJncPNuNTiWeFcFK+dnMBTByKpC+dZYkxFvO
ET1dog40P2h/TgiQoGfzPiRZni47NwA0ASdn2x1yrODqz4YVQSQ7EDVDBKZXd5MjO+Ie7Mxnqb0Y
FT8Wz32Z1EqF0h8UVN6g73fhChI71bJNwF9C0/n6Xcs7zlmr/aoWyQxSnliXykCAjn2fsec5YWvP
1PHxtvwiFdBrhRm4yVVkk6+4j+k4GeVAY13O7PPyCcev9xYT2g+L0i8cOPJMYP5ixCrJv1Cd7jpy
Di1l/IelySBpraTlY0xCcj3sZE3zOTaqAwj8uFfhgicT/62fQphh+Nf+FMY46T74A8v1DzugnARf
k6Fqkga3glNmbFAMr2WY/fBFGGV4wZcWX7CJzLmO5fB2jUuoUS6ckooGFpP8lMKfYSCmFl57sbZN
mL4XNSH9xdi0W4WfJfIilLbrzRH38cZQEmWDJBEsT5FvejwLzWZguzspj/3WyUZlHO50VzkM94Qm
7doyn/YuE0kqOUvaB3RP9dtmJcsCMtcJtdm/65yruuDZyiop8IHtpdZGiV7Ft0n7M0ASoUteaHW6
lvxZKhbchKuJTx0SkTjOqRULpd/MwmrWCEBVZ2MXiXIdXz4Dq2i8LPFMgRljHbo1T2JLq2y9gjEW
eQ5S0+lGVogy6upbkns3q65JHGNABmm2MhadPA2p7KMhOgDdZ+eqNG6gsO6mRBQp2LqbThT/zmc7
TUUcsaQSb1JPxqxCjtiWIosMOReTxvS5vjIdr6J+aE2t7eyqAUF1mbZirD8GlHNyPPUfbJUvFPAh
SCm352BtALZ9E1BCV7JIUEXxnoXML3oPvRYhiRmRpByjOP5rbc5fY/wBp0kepltORpfn9NSAXl91
+To2xXGnL5ar19Vb1xNJSQ0KVuw8FkJskFiDrsna8JZeKSGDsIvr8wBWVcSK++LeRamaSRk9Ow6Y
ZuplZn4nliCAteVnrvMyv0fyxUofMz1+BKsH3wgHNgVadP5jvLftGgyk7v7pcln1xXttA6GLQTjX
pULTQzMrIvu3zUOEa4Qpglz9K3/1CBV5RZIyGGxJR01UM8O85JGRRVyuwJVT3mKc8waCctBBXBqY
DXEs2BC9Cnoy8fS1xK9G3e+PmhV1+/2a8NCYCom64t5fUxdDyYf8wIpZygBzyWMcLtsX+wPoNXA/
ZvhB1PR9Aol1ldd9kDk6BZwfQpXL+3bA7d7ujRKzKq3fl3MFowuY0mrQVpF//sb/oh3hwQz5xUGH
y/wi7sumSkZ9O8d6a28z1FZz1zd8dLaGBDN/tnd8ySbtz6wBt7sw/UF8vaTb3BA62FUCftlxVU4l
sRjS2E+N2mjHNxznjEkfEmApwwNwgwpcLz6Sa3XC9o5+2zyAfvf8hHxaVnGwXwXVtV+J4tVGPrJa
XRVBRz8XdX1d/tgQcJy7pDTdqMdqqavcllsawPsWEBgxLlYLtd1qrEVk+yrrSKDRbprQgTsFmepI
m6KiJ2RDBpEHwD8GNiKRX9ysN8EW0elhZvgvf0sfKgL2V8LM72F96y//GRTI3Z+UrlTtwT2yr2a+
72Ghjp9Pn4U1UqWmuIgdtNmgDD+eKaYIQCQjnO+qg9zGb4uXlErpaqgE9/qG3R1RxkMNMTpsa0/q
UrCkOv8/3BJoC4OC+rKKcytQaHyGHcHY6YPi0Gn1KV6qDeClwPyICzN9qXlccEsFdsWjILc1VP9c
ERuL8fGLQxTN2Gy69HGAQGddWu8Yn1/yaYcbr5wCj+fzHx+GUq44s6fuNRxhakH6EHKRLClfR25p
L6A3+QGkbtjLxt+mq9rXPGHPVWPhBdUVqkZE3Km7OekQD1oQ/BDDyz3UFms1VhnzCfbkNqmNx5iN
08rOuiX98Ldwy3itGZqTX67gHxdR5iNnJvNorYkWvchNg1R4GFiwZ1WYuaAg4PK+zLQ3FRBmKk2K
JzIw/tczteilR/ZgLPbZijrgNiD9ziH8ZcwfMzf/u8Ccz3GjNBB9AJF938ZfvuSnW+khOdV59MhP
lycy2NZ5cvKrPymSQ7RlU8xY8K7IHzpqTHFWA1Dmu4kznUkBwpgBoqpBNXApjXOAbaycIWhvoiws
30v7RgFPsDstEyNHwAZutThRbTYgucnafwkrmlqr0imiuoZ0bqQ8FmVqL7LmDvj2ksVqBBN87uq/
FNVpTvTROIWk7Nt2GqYA3NZSJYYyu30w4pBIsVd23YvyikLmmdDkQEWTn4OXlhTpcS87vHAkUaWS
ZWjlh/qeuWZ2aZodvB5xhzv6WDw1VVoqqQXotOTjIa++e26xh7ijxiOS8yoFu3gpNg6DWkPFo8Zb
Pb+fFl6Dy+ZF8Bm8MhuL4RIGxDWNyaFFPGumSijukBMRt2sPBd5fpesxjQEcbuGupFLrJTvPKjw6
LFLXDrQE0XS1HyNMMbfGutIfgnguF5v+GNgaKO/TYekcX9hx+2x+egzOGpYsbpcrp3m1PDIVC3d/
sgHl0Lo27XMe/IMwRFjr9xyv+0FpiTaxsuXamEoAjpdEO6isj1Efqgq5xUc3cxtvVdudno+ILAy0
AX/lAwPzVZrTTL7GZxoslBCnK285usPqeHwz24nVc0J92/eV/PSpT0cLkNjnjycmDPjf+elU+lX+
nvBW/mjs04j+xwHQy/2z8K41ZGOlHzu+LMXOTC59s7i4pWoDhX8WsdO+FE3xJu3FbCetiiipejKQ
x6agO0jIssie0HpxBdg13TOMCWqULlki0nLl3AjXHdDmR1yuaVu+wP/FA6J1Zjm+5ZRQkeFgqCii
hi25EbkwdHQyS6wm9ADqmEJSAWp8JKM/V3zKd/edK8PtCUFKgw3MEyI/zwu7vxSNn5juSpXmFvDV
qnUe7mE2ySQiKhmTn6bHniUbHUs4Z650kcy7aec0AOickqX02vhxSEbrH5fFlDwcxO85ob+KM5jq
bwy+7HdEwIQR7IpELno5jh6KE9MMKKy3k6mCrP5jIOBHU59MpqPyu/VBAwTbRgLlYregYc9XLL6D
JznexMPKjROYVw23cRchzxcdipzPSG98OS99qHQqyG/vrWIKFMgxUOCDLgbe8ITgNbbIV54jD6tp
Ua06B8IHzo6rA1APtEmvSKt00SIVNVPIcIMZXce6SfHUA8q4Cai6xum1nTHQfYeE2fmJpTfq12nG
V+cyEfM5GiM3DDxP220c0QqUb6beLyZawIf+wxvr5L4MG4jPNm4+Obtb1egIS3rZEc2E05hoT/zI
7kl1PQkFdg6IfAsvFZC5XMO7RfcVO8e4fEN0kt7BaSiYAc3t2+uMX7ERxwnKeQnmZS7GQJr433Ft
SLV/88hMD2ZBVal+xO5S6eeh95RN11eljwHUc8EiDEFUtc2iEG5LNLE4/4+AopjTC9Y50fjQ+tpm
dFTcmOVpTykB8dN/m/N1as0chxo4dC3fqztshs3OXy2P3qzRMoScpRwKVaXFx2wAPYQ5fv0sMZbJ
+AXHt3K+fXrvKImp9nfBMiBs5j35iPDiuLkVFN3mHFXB5bhCGrr23h16Pa7mA2Rr21XwjpTcDhp8
G9Nv75GzbITxkTyj85NMEBv2tBgVeuDkI9yLTDzx75NggPQu/rXd/Qq009zG5PgPTkdpgFhR8MZE
yvshVIdUKIvSqZzhgsaSzxU83KBJNWG4IMi3t625Oadd3uVaZqaJdaaT/AKY22BdVtBBvYcbVHSv
u2BJw5w3VY//NkekR3U9k70XaNyS7D7wCezlXaPMw0bYZZSssiHeKoROKKX5W1hTwSiEL8hW2E0m
sTRe23tAeCdmiYrd4jBUFdsoUKEW4lY/DhTCLDMmzsEjpOgHG5fJoVBGIqH3Da66abo5kCgZqVxi
0eBxmrTjijWeYmGliYZgd9EhMF9cxVdKq1usm5zrrw2g4bOJENSkwEy6N9uCOI6tGOG6S9AfPRps
DL0LCAGeXDTaZlDZrNMfF/5HtBLfgt/jTJjDba1+5sRc23m0tCS8J0bWJbKGyXb9uRYl7+hdZEhp
joIhNeff0LtQGCC2lhFiwj5xjwaINI1cKEVZUXSz2qCUBYM3tCPAkcl7bS4AXeezgelFWaEWMvvm
KD6TXPC8agovxxQZoDlgNTAOwXZYEHi8ynF0Jr3x3Dx8BInKF1GbUzNPyGMbRvWE5Rl51EsYzX5s
1MaedF3H5YfS+vAh71E0Ipo/K2iFSdbwmQ9f3xr36yj4SnAiVC8hSzWTTnMnc4XvMedGCngyEQXz
NihFOojwQNiGgxkUCrg9vDcofMPmjxsBdS9oOds7m6Rn7FsMk4fQMsP3HayrW77TxD8b+uS84Bw7
jnY2Vdv1oAO80b03EGu66ZT4r7Eo7ZufqYPQpzOGNVUDUZ0o18oHW+P4gBwIQsxVjo1OsWSFflQ1
2uCIJOKxvJzn3sdRUYs+kGS93en63YEnff4p6N/e7WQpCraS2iTdoDLEIuvQ0yTY2Sth1HeCoiii
qgbC9RfU3oiT901wAe4MhZwX0ZKzwWwNSQFhtUfGmbIG2dvoJ7uKnLtCUxbHenQfCvf3Gg8jUQxy
5ujcmIGnmrmnWLj5G4iIOQbJjiHc8JXqL9mmLZxv/jx369kqAx/ypZx/sJHQE3FXWZIunvrEDHs5
4SU6u6V/htJnklSmqDCV4kglgVf8xFOmLqJNl1tNibB/L5Jyt/5X5fTdb3X/h4PCry26FnhzGCE0
eGeI8YcLJF4uQOB3GNOJOyOeeM6LlgdKMBj+s1YH4gU54SFXnTlS0qJi8EjQ9zrKQeQF+oTiKUJC
h/gvmiHt6YDbOwdfJyXWf05VDNasBTNtiFO0OfjGmBp33Jj9474vfkeXtvPxmhb/C0frsTmMkpYR
l7UKyQD1u6qOnfHlO1sxish2ItzQAKbXtD92w0Jn5qm998wImSzqmivQhHyHug95lrN19Llj2Zil
xEmPMGxFjj82PUCZMO8oO4hqEkRYVQp6xNiOD6rZ7vEqhXPg3Q7uuAnBOQuB0LGAYsbN6FDrOkxM
NjvCfbqaPuW7FAvyzkVxVVf8Lss6ZfAXlJSRtQe18w21CNFAlw9f3XYpUXQau+3gn72pGQ9TRkbF
zxLhznmpNfunUBqN+WGi8am5Bpzh2F1MGRX/wOf3BUmrLlOhPP6sGkG2YXxtgbsGHKdX74nNK3tg
g6KzQxfthB690lU1jckbAYq9Pi5GHEU/UjPIaYu9KkDHLO2MkzB6oINy1lP33LAzX/sn5Q/IXymh
sv97Xxv4n7GkS+tb45Rb1GtAzppA6zdWHZNtLJn2rmUfUa+8c9T99C2bHzj9Z8k2ZY2SipedAm1B
PZjJWCtUNT3mJlEi9/9bFTEGgLWi23jg2nsV+n68WJe0EVf9TK2FNsrRNydemKEQrFVJr6q2LiST
A0vRLPdcVyvHuHxJ2I9ZjaXutYuauOZ+xNktMEE4nJvFCZzm5B1bLA5WP0a5dfKubY5GsLjRew03
DVjAqyhX2WD62kJbRcV2Ef/EHMnZOEDiqFo5oE9wTuCwdVIkwwb9+OmAd/IYLeJZtoeOGE+fWCUn
tS38NFqp1G9LBF7ZFPp58cEXtiNzj0btjofb8Xi+l7UeJi06MOuvQGs6E/EqYXv1/LIGsr/1ovQo
bXbq6JU2Jc457aJMffz4Gt1rj0Cm1qk0mDldST1Cs+B0s/J6HlcJAjCclmB+2/oTQBoj16ys/1M3
+/ZufSbo61ilRpwW5K6tLAPJjptJ2cbjxDhP0dd9q3kOp8RS41fKsTQygyE4U96YHo0NF00zw6Sh
5KDOQyNXFE0z3nMP3DZ3viKx/3h0YChK1Gas8gITmDMj6YAiJdicG2sOTWPwHShmvhYL5ml8cAt+
7mEsYSjhxbYZ1mQZbaf293ouxYON59kX9PV1eHZlWA3VAoR4lRORxYkY8okby/2d1X9LyEqRauUl
ox8Odkad6c98mV19BV1uS/y18moUrmzAw6kJ18Z/ou4G1BHlcg+5tp7j5hWgdDu81++jX+GlQviL
gPJqqlu+gZCbIBQ9KVTiaXpGoA1JCDCISmjEEZaRpiTkXEvAIBGJtCaNd/OiDbE1jgAaAfhWTITQ
qzGg8dMHhjoH2bR9y6aVUFVmMg6f30stAifuWRobp3Cjk83J+5+dd2oQwJaAZm3WNVlGwm38J/K+
WnPk6hvwf8D41SSPu2Ov+U72Q/0JPzdhA3JyiPgqxCcLFpa/b8sdkPwCz92uvDsDC4FW+g4OnT6O
iKCO0yxk4zchWKhRicOsRHeYeNZ6tyRDFXrx8ks2aX6PESZ4AL8Xlc/UKpeiPCzDGSCymr/8hHWy
S6qsC2q1/5YwF5Q5JvzmsYZh+59PHLhbBTvYBvnf8gSyXIOch8e9oUnuIFj/fJd5ssHKq4qto6eG
S+2lrwVuHE19pHni421amUu7Y+dF/kX8I4LVMCIZJQd/sIFtWAARYbZaMfc02TRDNmkMCsCEKhNp
i/5Db/fht0WHkKjpas5qPIadDmpnuVFh3dWxMmFtv3vfCkhtlts9grOaoHpokgfZ3NcNpAPEh/Ui
ZEQyjcPUhpgIOiyURjES+hDpq0BYENOVrKM9ECOQL4UlT8UtClHwEKoPaRlkUm+2J5A1GLnQtpfV
lTnLXd3hkgd57Vmr9VS1BRFEwOiO62wVU2We7zm3KKHKZhZeVcOYuN+VB1QCCKqlY0FzrhALvJx9
D9g97TqKhf9m6Nv2pEcHmLXpRIyXNhN8obJec9QygILYRANcM7lzrG4D3v96QRE55TNnXbUf3MWZ
uH42yxy5Jorocmr9ct4z9AIAO63ZZhJTvO1uYaWAKnxw0/YIuPoHg2Nxl5C7Butq5BkJyDr+b1EJ
VLqx2yemh5nL+GUtTGhacB6kne9eRkaZc994JmzzxwlUNbzUURxBz4sgK3wAIbXvjKKrVDZu1Lci
zZVne2RRJ/NPmN+I10nLO5/fZDHCex3CX0Hs8LSq38wyCy+fTz7hRxj/u38dxYR53cMOFcb0o/ZW
QFjKzpxG3olKTi6JeU3AgTHVnIuZr4Q+LuoFPBjLlVXyiuUId0OH6RvdnHAiSBOdjemMpGx66xD4
YynTxG6MtzW9KMt/sdJ2tQtBg9pNyWq/PFoq5hf9EBAXmvZJenO3zIAAMSPbcvsMHrBIjhn+TJdb
fWlSQvioITXMmYwbdgdqsNFjCQMjo0vqUF50FRTTv2WyFC9mRSXJeF8go4L1usPc1JgAU8ds2sqh
paGBKUlQxbDESCVHo+KMfY0/94RfySOLm8UEfG3veoSLMkMRgM5LJjwmmyyIuKTH+MTnATKVXpMH
X4hG3oZdgaLcPCCi8ioYXKrrTAao1WTv52sGv2ylFAEwulROZIUA9yOr/hxiu74tYeM2e8kVCgcu
I19pva+X3CKIv6pkTnuU09xkj4hqmPqWxo/s/wlez9iiAl35hmZ5Ea1NrzgJvsQYNAcYKPvLE0qO
XSaTpSnPKUtaUyCrB/mA8Rmq7D+G7CQvdgeTS38cB/Ln/dU6w//cWcCuK99HgcdIDDKJ8VHZ95Wz
Reumcyypl2loRo4+NIBKvClf5MU6cIsPL5eXX3On59+lJE1rmxC5eVmU6GSZWCWMtSrnE8Az4Lun
m64fyjZ/AJpGwkmitaKc+zvttCQIXxAKkKdULyRSEnrawoipnndmnduh2Z1XENmTxYAfFV8wrriG
7jWeOrfszv3AU3mI4jp5POzbNXx++RQBBU8I/E4JvPtPLrSKa0SJpwBGA7X4E+fUlzy0UsAlZGdB
RRoZNC5qO/JAZTnVraFKbYiCZJx4sYcFp8w2u3Vv3IqtqPIqGe9JJw/NlqcOfVG6BC3q9uZz4UIh
H9yrGj5PhCugJbqnLtKGpVxQ+Ol5IZ5bHmsVxd/bMbTZLLj6lPJTDpNNQ6E6JwjwaGOIHOgcMNwU
5ie5IKLXILY9cfqNzIY9JxK1pKP77D9JlE73m1C8ZW5Gs4mO6lhcJ86F/9KQD+YpL3eC8l7YKn2S
YKw8EpkCcqtPsbFoBP1MpfkENSdvdyGjg36BxO2Tl6IqBNfJpS9q4FIJToo76rski/j6886WAycb
PuhmP7W9ajXpL2QdG3u/wseHMBpBDd3f3FFKcC8SHp34Dbsuc5DKc7TbmLgI47UzILmmknwR3Q56
EuLnao8jzD7PG0L8YRpPGvv7qTtNXIuKZFTyTMdMh9WlV2sKTCWW/FaTe3+zxqiNYzGn0zmjeTYk
znmApiQnNXAwEy4Zf8ZyR4RHMvzls/lB3QV7YKcDjOV6CEwtRMvVfCwQGJ4f/uAVDV0l8pEUYNHG
2iJB8LPyT83alWhzprBmA7DpVlEyedUuihvR3fY7SJ2KJDRYJNuA1d0jE+r5BBYAVnolDt4h4qqe
kWvFvgo0CKUrsFxdz8M5v1x3CM23gc/juao3VmkOqXAgekUms/82NB65nJTHKRFvRHXgLnL5UwPf
DF66GMpqAA0FZmRt+omTtnVmT725Benr/uWyls2+li/5OptMaRssMXPL3MuWB5QHDzc+PlP/S/ZI
PuDMllT+Wq83TOGWlen9eosi/E0uimuW4T9bFaxW9Khro72+/y3uHZUf7fCTeGH+24pZM7SjoZr1
deg8E0ppffcdtbvEo0ZlbCv26qHUjcgX+J4uCR2cQrYgWIH21k+mD+u6YteicdCuis4lQKDAQoOD
BTunz9pXuKoe578lFGPp22zJmRh/abfhnSbhMTVUCm5PNyxKiL4CEbIqDr1DOME+92FRAMiTT8km
o3vyUWfhbCQ0UxQnX5DIwC4r/uK5WF+QR+0Hq9BV9USAwuIX5467kz1B8yCGfKyZcUxXqgzJuZbq
3ZXWHxFY5TitiiY016AjzNt2qMTPGmj+Sz/TBhJhRgpg+k5EAhR8p1Z37VDLfDHXN2e+Zuw6VHEl
TqG/8aMxwJx0v3DBpyctHsjEeZvykvyi1dhiL7cLJHkOBSFoHw8tKxKdLZfkgOHvbLhQ6Y7MAMGJ
E5e9ApHqyfdMpZR/tlzE7nSARcuW/dWNGUAg6CQH2VWIW2aISW3kt9w3w8n+8cOzC1oTN+uILc4L
cgxqO+ZpvQg4b2Ctp3cWZjAoVi7i7T1KMVvukNU5S4g6uuflo8CIg18UgdWgzCF7GFtk4fPC4QPx
OYq/USwXVMpSV00xbPJGGwTO7juC4rPyhRWMtsP9ix2kit/ogWmuD7Nd3yBrcrgmgWTRigzdQRHg
pnt68wb5HMeqw58Xe2nJ+AaReOwcnCvflcOiRd9LxoxzdEewnvE51natvsaAhaWS7ZlwsDbALCVj
zeaE/7wbul35zBrXyxCCHSfsv8dvQ+8Uk+fXiDECEfC3Kqh+KIgkmB1Ztkue3aY/VSY1LYYyKxA9
6j1xH5dyaByONZ9wshs5hMycoDA/7UZN74aecs9u4IrPwxGzohtvYDK36RPEsDi1bvxY6sKnOWKJ
LCGgIBJAYI17n1OWkCfhBHUK6QNssh283t2nbgXCVAdt6ZQNLLNDjWkhZD42txf0isdVZRFxQnXE
iLgENyYwZiBzbQevTcPYUt2nkWuOk26d2ToYOjFLNeGj+sDett6MnU0nmgcQq7/a4GsJTBiYr/HU
f+dFOlGEB0f5JgPpkMQbhNOtXMgYChS7DtWDd/H3DObsS2BV8+yvpDHxUaYb0qNY0c4B/AmPwuvV
EoZlSQrolQbDLJGsE5jDaG9okVFhSkwQpsdPQDViU2tjqlqGhTclEDwEv9voDlPbZmWEKOqFX2D0
ey3ORfj4g88RU8rfyohJyAQJy9TpG8NPMJEAUJp6wWE0T+6VagcAd5h842t+VVNuACR6BZuj9Avp
wCHlQ2iGtRTmozudQZ49IUDnebRm6kKll4zBsKocNFgWcimFRVQNfFdovQEu82I8E7oyuH8UJPzt
tVoMpYKIN37R8apN8uyFtrprKory3uHyFB+qAav8sdVLLIgtTVuRKc6i44jSsPCfW5ItUeWx5y98
nQEv+6dKOpPZnL8PJbMbc2WMZeigLNvrwihYfB0stAAfcY8re6e7Ri8eKm6pxzcwCFzCFxTZvJ+c
EyWBM+CNDE3iEOOHDpLthOVAja6ncomknBAbl66/6pg/EjL9IR97FTjlJcmRghb7Nr/Yc0GnZBXB
lj/a9C5MseNR3r4w1WCWiYhvRQ0RYPN5If0kwfb2nPLKtmNx3iETqhgIBKtwm1uDq93n5lIO+kqy
fezezG/z9L3FO0mjo3/NGar4pGCXDDBYJZ9dcp2/CL/AfsuzXw3dZnIB7ejNmuMpUSHj3hKi0TKt
6KVGCkbnLDBisCTFLtbUhxhIBY5mfVLeiAUdRYKkRjb4zPt+ERdaGXZMycslF+TJ3NCxELlkzhzU
CiQsepSq8IRWcpNyqcPDmXB+GXQMm+078Q1/xvZS9BpLguiWmkxh3x4PwZiOGK6N0DnEYMzp0dlG
KzvQJF5aYeeaDcbCxTOZELJfpIdFuxzRSff0ekYXTfwIt3EoXX/1Z5b2cXdndGVOD4PmmKANp6oW
D6AvhWy+GzgZhFmco2KjNdc+/itYv/VfYyDJqOVFB5Li/BA8wzb7F5y4wug/9oAGWovRN7SiKeba
GzmLPhD6qxdUL8OahtqWqTnL8mTf2xiWQ/MafK4Zg1vt42jVybsSbsw5x4XS7/itIMqgZnJoiimp
XmFJrRoNZdISEY7HqzOV3Grg6AJPi0bsHqzJD2Oxhc2Go3O6nAi0lgfeKeHT8tFkIMGLxLe41/7Q
sLSCp7zzyYUhmgGP72P5VRbRLxeLxeV90z2uRTYWXhFgotno057OS0DJ331T58wK4+l3e9sRmgDa
fZ443C6Hx850478oOLKvFv7U/m/95TP1dSeNsTppVYsRFRGBwgAudl14h0Slr3naQzTAqH7JCzDa
qbKrQ54o5bN2xn/VtwCYCSmg5/ZLaQOPYG+PY4EtWK9eqECCC/wa+utC0ZVmN4DLc6AWYsA4vgNA
v3k9164xOQAvTiSYoJmIzHLs4HTvvuhmCZozLZvF9D3IA/6AIjdxNlw5XUamXIbiczqnKBS9w5n5
5o/ADQX93T+VG8csdpnI0aMTQNLDRw6u2QgQygBT2Zts7hoz6ylx12PMSJfJ1eBDTtGgiqxDxfu7
vPwipeB6DsxADte/JrZ4jaoXMC3Q+2Y2+oUdruGUbqYfsrNq05fF30tD0pHBwlaAZKlj7c7fjeam
14BWi8Ufhm7le8iw3AAIDZZO4ecfq/PihVvdHNj9V5cEOmrs/z/+Xx4Hr4MRAiDUf/7wYRkGoG2q
K1ika30hFFOb3DZ4zTDipMLaXQP23Flw4Ulhxc0hLBrjwb1glGKb+KhWK9RoKzDttfZtKtZM71Zl
/ZNJM5SbdWZXGjqxhUGcrNrjZ6e7phBsQ8w0+Mr4rRU6ZAvIL08HLEo0DvXN1TSU7x6PfF3/hhqp
obF4FV0u3z9IoMJz1Zng2xz9zWvJkl212YXjRu1di3epedmrbhIUwmJqXLUlzAqzzjjA2qykZnLQ
uZXbzfmxb9rYqvgcKAvbvdUhURhlSherkqqGRq3Qc1QlkiyRpW1uLdPWHTl7fA7cur6yaYuBSAwJ
zU+1uG1YulGotQmeEnHi4S6es189K0l/QSykkDWodp25FnV3PawRNn5EXzwFVsfwSi+GoV0Fh2Ad
kIqoM7TRtql0UO042pHqSIQ/13+IIZtwzdCaZZ4v4VZoY9pCWbZSXZyMsw6ltNZeZd7bS+QReVMg
0EwW3Ie6gSosnp/5uzTWfrOhCVA4HjISIMotGLtrLTKvTTz7dL7tUhX4vmbfolEa7XZ+ModHG/dg
qMFXm1X36VsJmPllPwBtoYhh1cgqvg1TgBharVnTOKzbDVGGz3p0H7x8eJrALC3eWFvrSj0+ay6V
gLCmUFH04jVYcPAraIA6qBvUuqfygf1St1g6HNAWkN/ADxO1utv2JZk6JTtyhGTWH3PSj3x5lguN
yLymbWvGvl72xImpRpwiCIiWemAzLdVYgnu+2sDjZIzM0xVDqykcH3RbNCt+ybqKqrGJ0ZnbSUSE
FCu35QE7yCCpZYqWRoUlvWz9ATGDfUZ3OU9LZLTMeNQKDutSpkMe6h1PVlGGPp8JHVNiBzQniAMg
VtcheCS+2omqXUHG2K/xPNBmxtC5hI+Eem7TuKCNMVJxnZfjgYK4LVTYUM329/n//OCr+CAgLYhW
gxoCwgF++DbkE5Jm4XaeZhaygCiwygDw4jEhAOE8VpJd2+AUEfDeznWEIK+IkKUiYxIqZL16GmT+
rASh8d7Ajxr6QO1puP090+PKJwjB0XS4YNUI+ZP3bCKOLW5v9JEfKqt3gjIh3rE9hx9IQW0/h8B3
/0eQdo1i30GhsgAwuzJC2b5KnCDEjMPYvJYnkFqZ7iQTNbbebLsgEhus3IE3xHlMR6GRSYldBfRz
CrOMKLnFX2YnKPVssIHcLI17UCEJWwiPJ4Iu80I2bvlMPtP4/APGIMNAhMxCtLx4wkK3yw02vkWM
e1NWi7eML9Ecx+VnrbKYrdCTN0m+s0GlmrID6/u4zFT5F14GuVjWDAW+xGIxPoVHQcA/H01uwW0l
n5cIcTF/i/5t/I+1A+FNR/6go9umMgU5AjfMW+KmL/9GWMJ/MoZWtXbq6kxLLtWNQOfSLT6IYvv0
gcB9avKbERgx6w7UU7bgd7NRUsskBxUoO+UL1AXzvRWb1DJmxtk5zBLtd8xuTGwaWxMbnnlErG4t
35B8IVuPx5fSI7kUZTU02RhSqWF1Prm26k7OCHdlPQ8WOshdMeaiqhSbMYH79MIcO8uQdXBhgu1s
kJ8d777IqWcnN/LrAWvTWY+d62UMwP6e8bSihjonT/+Z5g/RUq/SP+BXAuchTgMiV+cqXFClGck+
Sy7bNr5GvlVY7yk8PWVEL7Ga58OTbSiL5PFYaelPO1eQ2f7aZPkfhpfHYDyvo4rjjp3EUeTU/1En
81MtMl3PfYbH1PLCdYDqRCnUYuYNr1/rAFPsBu2atwmQ2LAK9UjsM7W9dZjD9zE4mFF3Cvpy5Rfo
/aussFvTYuZcqEzq2mWzE67HQz28nF6BbrVouBkfeKZqSyogUamH4hPS5veitzut+VVy3Lk9USQq
EtpJIrSgrD9mz0rntakaLrWEKTNoJBzm57RF8YA7dPkOoCsAFYK4AeTMWgdmNN3kuAzdbDY/qNnq
YYx5o4bWR9XZ2EvTN6CyB6zXuGFBc/i+bKTZQLgjMgRICu6DTPkI0dm9ic7tWcCBfKvODDdL+DRQ
5zUk/cMt26vf5dWmoC+EURcVullHY2lJZWw8yuN+C2cne/UQEQQOZ0CQZwN4xJTB/yJfj5Hk7aqw
Y0VnvdE6Y+qLvw9i79r2MS82iAC4xBg2hv5D73gqM4B34uUqNtxA3KCiayWHsRJkfy+Tqo+niJz0
gJEcRYZFSt6SvatiXeyPK1kZ4NplF7uo1AhIop0JhiX2SdW0tOFpXhJfFkDOjzXgItnzYlJuZcCW
YiSKtULxS2xF6AbkvwzifnAsSM2ko1nTJcmy6v3HNurYxpkCHHJQPBCs7zzRZcjeC5pyb+oBySh1
mjWL0xlv3uG9UklCRwQBcFKwzDAQ+H9rMg1g7Lkpqyhi6Tg+blDKaEk1lJ3zFEEOcc6Sx8u7mNg+
zXPxrGam7XZ2r1eVzk37veWU5/9GAifs4EHa0BPs0i5D1yCgCAP2Q8RSsdiIPbdY9w3HKQpd3dxQ
Q6Gcnv0eBHeMUhiGlrgFPaQwB+oFQhDNUStDbyG3rTi9l6+O/69OQLRr+TgLlX7XzCk7uJcbUzMX
XqOWD6pouRo/ThTeOD+Rlz8iJQWInPVrRc3jgLg7qkipmKHg0IBV5omMLsO360iZOdC/IG+QshKR
rxE9o6ohZgh7nmbg1rf6qKgXxZTyC0fbEv1XpPN3OdLPEzk0FWKaaWK7J3/0LhARDPWICw5Y1ioH
txTL6+Fkek2c4U7UrHUIT1h9Num7hgBFTPrXQw0qe+jCXs2LG3A+OCF9vMGHYWZUL2gN1l4J/Vyz
DmPdWR1onxvxU0fsQzZcvvyDfL9n7edkrYTsGmAK2/Q8621WYaZb83VDqEN5nS+FIc90VGtr6LE+
80xzCJP+Xhx23UhLNqilGfZX05/kJ/D0p/yhQpKVmdE6Zrt+NI5inGFeYfA/a0HXAPTQ/OSpd1qa
aBc6IiQFon5snH07F1iWOjygzeGnO2SItp9AoOVJ9gXggx8Jo30F4q35FsKdzi2Yyjqe/KjxXxV3
Yc6VCgudvz+zkt3CEq8rt+/EibrGcJgxxILvDg4yO5nmgAvbAmVn83NCSW/qXCwNlBLRgoVCqZVt
FUYwX899oilGTXpkAiQLYLPGySfMGctQbzU1mdGUuFETaYDBLeekmNxeXCpyVL3SOZ7LHnKMMRp0
94FxztJFuza0R9VAfRW2xcoREyeE9RC+P6iOGUMsKeyc2iK6h5fPHwpjEHzZS+HUBT1CvoEfqAkw
moLsrniST84VQnl5EMotK43A+cPYnjLgwqqgja8/33+DdJRK5SQOF8t2QuK1DP3q8qQobrqJnjEc
60hVgjJuaBbXDMyyvQV9zh6b0tmHcTy0HocCDVrm0+IYk7TviJrJD0fIyQeyFckW2sSQfegWi0vK
geHsejxwE2/t5ly7utCbPU6ecdMF/OcXIgWH3DCZAUld9jbdz9JdEpgP5uN1NXID5v6F4WqqrTJG
o2w9tcZKWTRDzsxlIc9Lg/8M/spibCSeTH+aj9iANAl/OFsM21tj9WlfXu1vaC3u78HCPR1lRw74
dKoaUpFa8rS78vMuH9y1asf/C7RIhAXFARmxmkKbtefGeZaPhCAW3r5NpU99OCWLh/k12BuFNgXW
9f+N4mmD5yehJmzvyuJxPjw1wZZOSQUqSqOZD33ETC/E3XOVtHD4Ax0IhJNi7Oza6zL61OB3xBw+
Va+PHs5/2NnQSdFQeBoGCopBWHSLCgvwreBZGK3yB+XQRxPa6cO9fV64jYIXCyGZ6BRBDde47pxh
eZK8/4S9W/ONpDPmDwgL9VbB1sMQk/eJboHgP8yq7GIl1OPr7k5njySgkPu0x8hG1YpXNZe5FKKf
X3ll4CSgl+LYxC4HoCRCNM+sOH3F3y6AUTrcPdGupnKhKSNYQg7MZlEpOmN/kC/kiRwUQZifWXiQ
noPYQsaAbyXNrg15S80xiXT/3mWwz4wezcqyNl7tny3yiqSRp2PuKorBNzdWh189bbgkgM+SedHX
Jz739gM4MbgUEkGkO58Ef+uomacgi1T3p9iRB4/owDvGQW+EOsaXTHP849JFLFnRczCz8vZZ0EHz
CUZQ5ZVkjbY2EQ8g+tpg1yI9VDYTtlWDIk8BSxDK9E6mN3QE9PlUoRyaio/RgRNMN7u5jU78L7ch
u5Dy6k6rbk24rRXgd9vtC7Cn9+DYKBHCWSdvT1GE2GZBQFN0xRESl+p1sVxBA7rxX1+iRu4dxsz+
IhRyGNxoWlopPJiOaL9DOrwx3UpyY8kA+YuW1Vc1I2axHEEdhzu0N201bPiNlo19Y18WioGNG8rp
BAMpdFyNmfbV5eplex1ZIjtxYGHM+qbjNvpInItHY2xU6JyG+Yu53lENDbQGNnK9mThYTGybSPez
wQRL0n7fzROzFplSY5MiSLlVlRc76qKHoM2OdXjmlhBr4nc3jiH1CLbNS390oxnMMt5cAyzZ/gsB
BPaz30rRcg9KiwWwSrvQuwYxhT03n4Nxuucc2gwgYmaXkhONwz9JXQtn2kTMchTJH5v6PzvlyXnw
Tm2/3v/DfDRnsyyj8x+DDImtg5Mw1JYrwMi8/Z3VvZ7y+9c3CoE95DpIB7ZX4PlmcW6sg0I5lqJe
KCjwntOyHJt++13kB0adOwcuaWTqj3SY4ukcgg0SRJhqtMJcNMF4aZBK9ktMaIq4WP08odtBxxcL
3aQ5uIoFsHSy5uwMLu0xRltq7qoVXn5P0DYmbVvQ4U2xAMtOT7i5044gFoB45n/7JhrLhNW75aI/
vGuLz21JLmrkNEwJAHQdqMyHlHexVQ6Z9QXZT+brCvIjPdlFxwpidcYw8Lmf9zy/MaFZPkclZZAx
YE1C0IokyNcpwtEJD9HEylCAeJEdRjhbEihpBKHTx9odDLJM8IKtbj8g3sSNDuOygauvpQ8q+feq
AHcVHDJCkyipuLhiNEOZOF7Uk0SYuJCsadott0BYrzHXfJDAH+KkmMTGRCl4HYHvERhJNHKdxMpz
BZSPe7hcclziwh7B8OfOIevBh6g+/fBOVJH6wE0A/ntHcgdJtOVCiMe5gW4aAi6tOEAugR8v07y5
NNxeI8wt+3VgVw+Qd5ekwRs6vOo4yogTSpgCt5sOxbGpCl855QIWX8hs8lyX/EnilFJaKX+MFQiO
TV70CLJS4XVHhey+aHWSEy1JqsQw74asEhFFT4SZNG8knANhYXBMQpsfA3zKjyNmQBWCSHqDzXPS
oZ6Inxb8QQt8zI9FMZ8z648Z5TL/lkjnDARny4gda3+4rC9olGgZdg3k6PwdkqieZ3A7vcfhTPwc
EWFQp4tBEwGAc4K8LM8PhTNs4Xa/EEs555NBg1rGIN6u/HP6EkkZKjneWMeww0/BfhPPsDjVhOTD
DTgKWrfhPnjxeUdUmkDGbgJxlNSDr7Z07yI8Fb6AuVX44sFwOF3CAWzMO9KS1MX6MG1xbnasv99l
LRPY7EJes2Sw8M0YEzNFLoiXveRK2ubWDSW8bTsLyWtsmJZrBS83qjo0eP0oG5hGKQsiqRjU2Ayq
BPXxkn/OejZvlgkxDOf5EOv2M2mpwGyeUmiZmT5LX6hXlWAG/V73aINeiTZwr8tTLg5+hAn/tUa1
ptrmXPxVFJJb8DhqMES/HZjxsdx7BJCOn887UaWcdAIQt+kO0RlI21rOPiqoPZmW7QOuriHxRzU8
x1BrwDkVnvlEq8Eve3cQ3gPNYf8nkK99DYM7V0vI4cWFgPOlv6yEym42M0Xz6gcQl8UmGPnpJnsG
7TGQm6W7wJbyvPeCXwtbPg0UH7gS4a+n8ENi6maTswDV9paf5o+ut1bl5E1y7sP8l6SooFLTq2mg
tbyHgCM/5Hjf7GNDSEsj/bBNWXmZeN5Z02RZu+7l0ss1cXBwWND89o7/bQHy5Jc3i+3hbbJC7spK
2xeAn9nMbYS/cCxC18LisPBHt+V5jdbX7zJl1o0rEJPQ172w/AJ3kTiVuisZAIfM3yUIisVendmB
vTx1uf7j71o/g2bQia1z5c29rRzuWXthdXwFOuPSbn3LdQ7OihO83hfJOeIiMsPPk1Q+vqTT+OoK
dS0TX3fvBpr8dgsJ7VmDjWvpGH52HkuGioVucmx3c9OObit2aMg3lAetuXzO1NihqxwKyh4aTw3Y
cGpgfvOau5GTCg4t1/p2s/2sXoJPAstmshhTXaCO6tvsnDip3KoY0hMr2xrHLK/RcveflXaZjf7+
iWhRzg+4Br23AJskKgICSakPufk5QV7VVqrD8Y3/hinLBlgQbK5JoYgvNpRovpbIVTctagyHf53n
jvFe4HWit+vdDbKVMkbkozWIzhPqOr3dPYnBXlFPBN4KYMcdXVvkIJj5+DON/f/R35Js0kRt8ijc
syB7+o9+z/yJTUUZnJgUDkytUk0wqfhGiM28Qswons4PN5Ernpwrn+XZB8jn+mY+2rBf1rVZkOXR
+CS8zghmgDCNYkcA2KMZH08qxD0iY3w9oUNDOeD5olNDtMr1OGu33fRtbGETRGUlsE0o24wRY8SP
pg7X0Yx24opDggj6sMbyeg3sU3atuQvYLwLaWglb5SePngn6v4mWdJaRtnW17kNsSx7n8qVWZSti
bJllpnvKwyBypM+MNFyPypGkMKOk+DcWnW5qFNhAa5x0/jbp54iSsxvBl+Nj6dJNSgQGHTb5/qIO
Xv6OU+pyohaDVWbD0LvTq3wiq2Fzw/taQqsnTbHWrbLwUUqk9nostlP93eLm/NzZL9NrUMUrqyMK
gibjmBtxD3iKFLwkzo77+qqIxTitt7eGedATKqI4W1Ppcx0ly78cB7vuzPvH3BGzUNTYbddT0wel
EvuDg0rlhlackHmBz2b1CNsbL8iizEgvGDcVqqMKrJm/cuBG6MQb5hdI+U9i0MSUPZmnIIUmkkyH
0m1tTq9lN8pRpuG3TeClfBMFJRRtQ7n4Aa7AcCDliOs0L6DJWj1zSGRjgOOI11wyp5/rJBy6DbAH
fvcOAyB/7O5sPf5NcLBl9XVAe8bXoflYWZ9aosWDjrnYXRQiNSqp6UErLHniF3NCnnD6qik42WuP
DfYIDHdLGxmrjgPHDUemPEcfZSO1QYqRUKhGUCB0xPNErUtZRhAOuNOM8aPcvHnobKHysUsiNPL/
0S24wNb6le/Y0B4N2HYGMDDOjH6dK2p+bX9UWNkZebyDQ/moTPdxprZZJ9Nn4RFFQN0rLU1uJM2/
buSZl3Jy2YqHw256rAcSgbWqJQ4R0b0I29IafbJF2fv9QaHlimQbpOhTnz6q76O34B6t1GAvcVie
mPPsfUyfq9G1vqSHLDv8rTicb8Me/cAj2wGE71o74bVLBpyyk+Or8ncGTPwBSEmbPKj781p+t9Pr
KHZXUNkNx0iKJBEoBtdjq/x7W7SWAlmdXCYb1Kx0eVDGFG5V/UHgBvyXRtKG421lzSUlfd8EoIH2
/9tlkYmxbB5VUI3/NmboHEaMwDfo0vZZ8i5dXxo+JF83ehkxdIgF8+psqIckbfON6vXw9k+nUkzB
gq+OnhbAd4gKniAXFxfPNVm4dgjmKURv0puQ+etScJQKS2fbsedBqGzaiXLIlnMCau9HBKp+cxsK
FG/kfYorXPzK0s+e0Pc/7iiXMQh+imKjSWZgiiznyfMvHQmlGiib0wYgrDfW3T6Sfu7dIpRZPIki
1xpHJWhhFVntHhdz8wPYYpSxhwHwsg/wrUFLnaBFHJme+WX6kE0LnqavahmyivqLmuyda1PE4zjo
zeCa55dmEEHvzWfYzPM7oOhWKNBSPIJDHwWu66cAI36PSxYHE9gKJQ+KivENiBDvfZI/JkLq1kJ8
Q+/wEGg+NZg4ct8R3IkzEJo+m9CywMckPIrihOXedODw3wYWKTwW/KhsqQTeHr75mayN6kNLt5XB
knbsrL11JRDWqyzexeNfUWB0HDv5Seqv3umSS52AtLyDX7ev/8AmGCQrLbD0KC+iEF3A/fR3F+ss
f1jhFHgaMb1aFTOcfzEbVAxIIY80mSt49T3wvmg671wKNaZuG9lBZNDewIxc1COuBTedDEQE3WUG
U409UQdaAbZlVzqYZjXYkzfBsmXSEP/q2rhLLqnA5iPjYCmFUjoh+KgzLHgUAzxOB+o4eVISxnSx
TeCseFVhAsQ6QS4lIf9YZlxMJjNKSFIHxEBIS5vsniFTadRs1V/0g4LlP3HzImmiqNsmPyJL6JzI
kUmmUSpaqK9exwzOSlFM4BgYK77A1XWQAI44c9ad+C+BhhrDWrbvf60Q4WwoC2YKbDPPvGMT+8YQ
J4s2AnjwA2jEd5FM6Io/ieU9gNrXpD4qHO2AOkLefRxEcn/z4E1yDMNXwsDcAgrSEMp4Gtz0k6H+
hLGIaPeehGZvdjs8NQp/Mxw8X1nIjbmxOz7/o8+Qh0zsUwCWSzKnXOQj4d9Z6PUZlw3h4UVztT7G
3dWPtHEFPnyfmyG81ONrJdRTK1jCbEBphatOJhyoyuBWdcvwHm0ABPw8OWlDlzzSI4lhOb6NgpFq
Bd1mUkE/j8fnQY7ELLNwcezlA1TFMz1ppQbIQ/dgFSSZfXpJpdqyoFgk1syZ425bPWw/9ohfjGlc
5NMHIa+2/DheeKqD0JMHdnkrB+lgWV4aLgICnQGCUzuQGIrmLeK6xiMYkVeMRZy8Vj/KgMlLP8qk
GJshPVjWeZkgdD3DwRLgMOdgDmD+fbhZSbSpdRfKPwfGNwLQ6PgTo6mSZBM6E9s29xolAL0pHb4U
XrnTHuXY+AgfWHeH10m0TDh5DtLtrY9uDD9lPhnJpHQmwyqKeA/wQIf6RawWG1dtqVtzEHh703vL
2P8phwBUmZJC+vix31DR6tzSSwrNsEiuM7Qigr/T3wy/gqLx7oZ1ZNrv9ocz0bDPDjaZ1vank8ID
alA9HGQ+3DKDkTj9hMcz9h0cNOTK8+CSD34S0B95L7HJEeSLsLU+0o62i0WebiVEl0mU0c+fiZcE
BeM5x4MReDThds/6kgnarPRjnwoJHKuAaDMnfrl/BtjBefXnzpulXpA3hawonE1srmcUqKRQ3dsk
D55/DNZ0ZeleowyYAQjg3ddwNHXddo5uQpDN1a7U0H2xAFkr6sbp0LrN0jIIy09h4dntn7WbV7pP
7UnNve7sMpL/+DGAJ7te+qCu/g5UGC9DYNlKE6Ye75pBuGkqJRLz+Ta/ZM+F+hq1lJfeeBxNY6dW
neVlkQaFYyPyhU18wyMQjk26B0c7c8sQA+6CO0kQYrO68KKrew6juZeXheRJl51hOGUXvkgbkZAG
v3ep6b1CwB+YMCdvgHIHx83QFyJz9QpXHQ34Lj2/Mc8Oy1glTBej51mE5Lv6a1vnDGxui+ovT5qv
XlCaX/AS+7V7rhB9/8muD5Z4DkIN+uIFTke8u3rEIM2iDG2lLidjsjpVYHmUN9ftoT+IK5KMN9k5
PaDkY9HYC7j7i0oXy3Cv7kekSUC9AWLH9srrrI7DPPM9rnbJaSVW752xdInctzQpqOhOyWgteFhy
OGbRp5lqHDAnLrQOarXDgb1yJAFm3HEDt+ckcUrysXG7RGorotfYsRWggJGdQszC1o0hRdcMo2st
AzLOsoGeV1/pP+0JV6opgDrvWSCepF1MvcuphfJmYQD81i0TnVN2KJaSuvoRRMQB1cMJLkcvJjPf
PgowhofL0Er8+AGVvo7Q0dzPIe3I7yoxhaWPBCOPxR/U/DLSGvCiZ8hfXHF1Vx18RWWprAYCkdzr
sYOW7oUVkNEQkvm5fQIIBjx9iijn2Dx2OtpErka86uKU5IebpyRIMXJsD8Q6WYfxrT+oy8a2MTQn
STltfOpwP6unu3Z/9ZeYrEUpvSOUMiYtTYyI6rt1JfCrxRjebsZYhLadkqsr0ZhrTWPAY9e+7JBj
bPxnJgp1fvAz6ZEaig14crWHqRhKdXnpLakCB61o565W//pR8ytojoS6rSUipuMYOAyb1NB9Q+HM
NBKIKpDJ/LBFmi8eZTZD9e/1LOaaLEQJc+xf0BbqFbVkacI9NiA8ODkk1YQH0yGbda9T6hreRGCV
orAVt+NV8sMEbZMEx0AZHSKpIyBhicnAJCr7JEGeCS3GM6Rlvn7d6KhxJ13ajypj6BvCuzIsdNg9
Ynt2y5w8t10n+Vvoby2BaZdnamnMjpYw4Ddfw02HPclyxJEnQqWU4tRAy6yzemlQlBjR4dZTl1hb
0KcIhpVO9/GeVsAabSAj32KNMB83i/lNlvkASS/mFi4qsIekUxIAK2XfN8sz4IlftWjh/ke+iCTb
Nt9ORhAjp/90R3/4pADi9w+1yxnHgZ5l5ucUXaPlcX0i9B95DxjhSHjaussiuW5ZR6D8FfBnEwdC
sCLnJSNYH29S/tw8fmwdclDpUzc8AIGIvwK0dQpOrKsOQhnuWFOS7JdBzr11Hsvki5FRGvGFrWei
LXXN1a6UDD00ya0KZXrJYAj/1t6xxwyOtIMd/ZXMY7Fj9ERUy/+yKKD67+0PVdFqW708rqAXwwxB
uLLzjgLC93CD04ah+eyxBqKMmLanVDXEkemyOVZh1J8GOx0NfdIj1fpHQNWFax60Uz7LA6yxxqmD
QcD/QKCOcBiOH8GrPo5M5uLzSvdnxLiTtsE4HjNYg30vpneniz3AUbBDTi662JHBsExNO+W0dfnF
kEDeoBCbDJc12FTkEh7HcFS0OAlf0BBRbUABFoDRtPUM2z1rIcO0079C9385t3zsRzwD88QX81kn
XaSCI45NiFdWzylPw1BvocEJwf2w3nK1Z7d3c3bB9sMINt8IWLiHBxCgMJRWiTuYExuxUlv/c9OA
DRYw+v1E2HGs5y0iqwkkuausQw8myoEp0Ipgq1JRnzxgN/XvH22k4yR20TlfCGi5oI8cYXUS6CW+
fg74ZyrblAhNhuF41LqjCac55tmGX3FTyxM2Pw11r9ieXtkWgokk7EZ67BVwV5TAH9Ww7ZdDUgpm
FVxJptQI8LJOy7HUCzW63aAn31H8UDMKWm0i8F7o46faARJY9T30yVvfTxKbZx7wp5d2Q6vd5pQD
At23U71B9o+xBIvAh5lohh6kMG/SMReu2QzoJWUI0VZfgMsi+bggyVSohweRTkrPlrL1yxLOmxRY
oeoOnobpWPFFTPD3NQMJJigTa9I7JGhrZLFzt4PPXHPruB8LHnuesqfLzZfxOO3EibDzIYw4a9tc
i/vx2+VruOmWwkDAwbnGA/YVq03YDYUNSXNRsE61D3gA1gm2qQWwa4f05NmCohRsSmf+4vInNTi5
gShVGhUAoyZKn2RGykdwC+qe72oU2pSUc7K46tbM/B1L3MXslCunGIHRrQWRy3frg9ezOFNPnBGE
6JasDv2pdcjc84wOwjgiKQavQ//n9hZKJU1w9BGPDXIS+vzktptPxT4URJxMnuosCAHsT4GIz9LD
5flyNMeIzF0dBERgr45ML3z+l8wHAiW01LIwQKD+GrM5MHg9chc1D7Mv6GUZApK2KbCdohDUqOKT
G0eu9Xb9Qk904njNMTPlTvuyLBfuwgFw8nu7hG4LQ3LmPgnY3s0R3tSQ72bXdFf04TKVy5fvlWZN
LI27goHkV+CVu6eSDWmbMugnGprrpy+PWPQAZucoUjB5wO5zsRY5MIkghJuz/ev2SE+fS8MIhbIP
zSDtYXZc+vjh/9JOaTZdmpirsQ2ej3ynMbC07YSLlkj5BlX8tI8NfZ6QGMI9rSsq1kUm3o0boGd6
/f7HtQHbF8sIXHQRPfauhGqGK76Ks0PPQe/zR7it3ulqeakrgMlbSVonu90GMSGysrF+JE6aKi3E
hWTLcKRyOW/PqWCJ10xAgeSsl0otCESx45N5Q126/99/17qUYgrDVBNLfAqDQINqrMkr9BAEp68J
TUOnAVxXv9TeiN7YuzULL6R7cvw8a3uMA4V+z141z6j/9zwaujAWvEst13pigGHKyVgkzHkt+448
MphOUxjK5W0CCqj4Hkw7N0P6XgNFkOpcuOoL9rOILAmOWm/EeFJU1QWnlURVEgXWLoBBjQtisx+q
2yCrWjH1Z9Q2aWwVSvTg6F0279rrs3FnTxjPl1eQc3YjC0rADdLHXv6Vd6A15keEqZefHENewQ0j
BtIQIBlsXNmcJ19pYtmTX4QrxBaukyvU21MCeIlV4vZBwpChreD8mbVz5y3N9p43Qb2uD4Afnih7
MK9WLHaath+qopT4IDOmNZdsDpTdA83IZEV0fdW+BpRFsht5qruO0fksNRQA3SvR/aMf4fDa4OzU
tPk2sHITbT01oP4tS2bu1fB5kgJd6CIbrsuxUjyAI0n7dv2oDUf1YxEnl7QxV+MSPyNYtNS41BvL
5ePLB9ydRl40niK2+0r2NNrtVOqXNBWQWOlQ/U/xrEjG46hugA+0xLwPpNhCj1BAc80dPKGZip6F
JVOZtdK5OqJXz1/eC1dKYh3YaFa/9abny8dqEGBiAG+p1f+1hR6zwn9TOhmqU9NfkJeY5F7VZH1K
JmY8Y5ArcBeRyQmwn+EERcByLhWSgGTrjTX3ECXIw9DdY1vEqJlObS4wmEuNA3HMKR+TNmzfrZQ9
EIkJjt4BaOQWoVI75uPRD/AIneICWM1MebPHtJchQbx50E7SR20wodFWPhwXhLks2gJUdn1jd/uo
qrbG586t7xHczhiYtGoZj2EV3ki9QUOsEa7hMyoKvZlcjwxue4B6jE1G5XDRx/vPAI18Ew4/JBTc
dQseza3d6nOGeEKiDPBLPwpuGckOjqeoM1kUQvpYl2BZYF1Qgs+G++CItaqA095kaaxUC3xTUpoR
SQ2q8dMDxgjWzB3YyQaMyURM1lJtHPInNDU7ZaHp20i582i6AOwG4lVWgP/QD62BdlYKdUEKJAmG
4ylDOcYTHrDdsKoBYc3f8ywAGannXgDpAeeEdaDZoRHFlvqw3U9cKl7mjBkH8zEsLY3sxp0fwlrZ
SH0uqglBEwC7WMEDYSwAhkCHFM50E4hvlRQOlDdTPIET0hgEKiFNMjQpsyKqApbupNXAmLuJ7ASN
J4W8bo+hPfBXYrBfCUFitm3MOpyzSOyMZB0VZ8kWflDCwznELi7ta9Ai+1PgQRphRo2V6lWIE8cu
4KxnuU8Of0HKz6hBsKGKm34s9m5cNgVWzs8Rw3LFq40u3RZWQ3B0OsqeCZMt01fLeHgVWAVK7Y8K
Dlw/GCVjn4ZMiBZPbINAZA34Wh1c028AxF7awUQVMMGSEh15bGvlLVW8B5mO0PHS4p02PUHl5wqI
beIpi837YKjeRfREEr30BuBkK+n8mrDegd5Pxdh5Mf2U3zrJ6/hzmJ7yZ61yOrpxWwuHBVtc4Ajd
xfyTorf8YN+/vfNYMf49hTAKxhT3YuiswS2LC0EalLgmiXZvx/XtLOH5bZ+mMmh2rJB8AZaTfbH6
HTp3qMRs91NF06lUcderwEbLljDVnH6zlxM+SZ1FLUE5mbbXhR33Vt8nuUjGLGPT4xXEfeOGrc4J
chQk39yMgU9L7XuEa+WVcaOjtdkCUWy2H2H5qu2vM4enOujVJ3emv/IyDWOO6iq85z8FNNI/Eu75
1xUkgxZk2tAqBHhSJ+jE9ZoJhXRVBn8i1hVtUwVg/Wn7Cl/vpZrjQtdUmHqIh6Z0S3WkGc1kQCE+
/vw7YWsXO1cgVwYikQ3yVYUBYyzFRC3jXZTwvBawtO4H9FckBWUjGmfqStPhLO5EOQWc7jJ1V0dk
WuOvSVR1tYBYcN5UltkozaCs+qOrwB+LhJ0hEw5/ijs5Alz6uzyJlaNXWowssnoJJirgNkmNLnMf
ifAjdZLc+G2hDhiEjtFOwwk8qEJLznSqB3dQ5rsS2b2wD1/gSnIEQ119uZHB5lKzjhZ1kWp2evnd
meTXLJb+pK8jTC4bdOZEdD9OFAmr+JwcWHItv8shMBhzTq6m52i//chYtBASzAFV4oDSfnkNZA/8
bROcSBLrCh8/uvlLLeZ77N2xjY9qFvH/CCrZwqijIhwPWGaKLl08uWxJqZfFzYN58Q4V/kG6VkXq
0dD5RXyuTwP0uNldkp1uExTpq/S6cpRYGMSS2lAUBFRly/nEx+p7l1chR0aZXw3BqJNDkF1fmcu6
j0H7V1JhCoykfrm1Sq50XNU8wqw4fHCTx7mxIPRYyJUN2vCkZGIiUg78CGYMRFCbCWiKbAqwkFrT
BEgSHxQhQEtHBmxvJCSPaVUGFMBxjry3gv0QQUps2ykmZi3d0+3NxCmCga/MjfQs92hTqq6PgfxR
vO4gRL3xWL1ezUC8ZJD21h8GXAy3K4jJ/kOHF+QvWI87wTipZGXMz9M+Waq7U720ZKsmbLSScdkJ
ZQGXp9eCeOdUyqGXITiRzvlT4a3XkeSa+R3bNspKKEJcXUgTrpyisvSjtq6VEY2jM3zVIVSO4t15
aEw6LdZWHCavhcLDNxYIklQkSslhXoZhXCA6pskJqcK3CH35eQwx0Tyb5A2RVFhoWd9ovFxYluQb
MaQVpTSXIqjn8RpaJwahjA4zb2ObY5i8kWoQDmPqXKdtuAPP0LcTmE7xkiMwiuzWt4hIcNTGeeo8
GM8pPkEsGBvbHO4xhKm2ysT4X25SHBMeQ4e0ulG+GKdrqduCzet9Jzw3+0q2Dpk8/gsWTMzup5s7
DXWU+s3vgfPCfPO7HySqEsIYicpLjqooBCDCpq62Vkak0RxayDtOQ/ae8wCwilKSeQHl6ghX51um
E4Q6fKoQs6TT/CVUCmnIbOGof7TvuOHsg7+al3wvnCil3mpgSzOWOzp2hdYL3vUazx++EQp4+M1R
jrAeDzNlgiFIZvaR9wo1/kjjVwc50xEkRt8ol7ZXJyfP0JIYuxBUYNuKB0m7ajmlrKeDBMxUnIoK
yDHLwvOzP738Iyp/cgr3rEIPGSP3whYd+MzXkFYsvPwQTGegggAJcvMAdHkHUOubx/44d7IR3t+g
FBYxAfhZmteYBQDTxdHkujInTA+2COqigr437jFQ4lsvQCMo7AmZX8wfYC/RzvX5lkwOiEGRXpDI
MaItr2hnbyMJXvWr5NZRuviHItNrnJvYh8N/PUYLl0C10tFlktmDJGXwWbFpSN2qp+9QoLaO6VV1
a9qov74pADSAz5eN4BIqLmfsRK/tmzV1kjMxXkOCQhwO580xzbQ1OLzIzaX6EgpJYrlFjzfb5txA
EsfAPxqALXbVgUZvIPl0P7NUzvp2I+yM/JTdeuiN2pb4Zskcs+Hop3spqWFN2NaBFYbWaj6yp084
KzqXa9yeUxjjDP0aWKjP5XPoWHMpaQDgrEe3VuDgpNPDudwAXvgLYkqXWApc3e1qnFE2P4CY5tx/
4OA0OYCGPJgA7rG/rYSm/o00QQnpmUQTfPVKYr9hhJlL8ScPF6Dt69QVwgLsZnPu7S8npJq2oGuf
K484BAsC1aL4y6yvlL0tFW82hvuFnOMUe1MsaX2HAhxPdBN1TtSyPRrzcNqbno3W6+JNHgi5vdub
GHFrcMZ4GvaZnLICFnh6O2f5R5OWVj5r4AoBFreK1F3/ZCqe9FAcDOqPySDFm4WxpngCkeCMmwiE
Kk52Q8dSZRVCBWdL+9X91ftp9CfjoC/EgO44cD0zR/5AJyGjCnrR4GdSMCYPyZ308f1PLuNMwR+v
TZb8yPIZkFxsRnsN+HmfbOOJ0O7DKuVQcJnvTz2NJgO2Eac8+g3EuNJKbrObOz1y4dslwm+82oFl
lrYMTJSTDnmp59FTrPg46j7kMfRKVDNPpOv4aFYZ3wSvlo94nKvI43CUNKwaIFKIkawjKhcsVm1E
J5BKCA2lq/B1isX97TTn+jFlJ2rBFfH4k1q8cQ5AIzuUVWMy/3p/MAjfEe47xpCPdGbOU73xf0H5
uyixEZvpKlm/hdmQGjqrE9Bz7oOlmEI7J1M6YgW/ZWIPFzY/UQjCGIUooWIioL/1USo8duw/lTXA
hM7HSkpucEjzR2FrktT5Cer9+8m8I+Dk7YAJmEolTqJkhSzuu66AzBuXX6WMmV2gRNaPHnG6kS1c
7vjVKMWj9lS79iLqWZ6FGxAcvugiPucGqOEMEWX75mgfgrKz0dUA1u4iOWU2Vvhkm67PxJPj9Gs1
cMM8dHBDnRm3FAIkAqlu0GGoUv3BKJ7luniKKRGltKzlokteKXEt6QzqHsWCXKb0zaLAh92medLJ
LVGbEAlSKDIxgbmD0t8eOhyZpVkmpyMqGSxMhOsUZsvOoTuTisKmutqoX9iN9+HDF0xGwRXHudDR
beB06BLWaDpVMXbImaz2rohQqPMXy1PKo3YQdtwl5nkO1HUZFjiN1mH2JGLB2Ic+5AceL+AjH+Sd
Kp5XNO3UT1sIWKzIND9aX+1Oxw8px6NcMsAYLQvFYEVMjVQBlhdyl5QAFjNVWlvmG8l4vLKHVztv
H+StWGjPVycDq+DVkByqxpjlDHiAT2uoasyFHsPBX595s1eeA052mFC67ow0B+HHMLw2dlRlpPqk
+zEyUa51GKw+d47ozcnwfFomFaEfA4ypBW7G8nvJ1ibHqkIXKWRkWyLJTEaYNBUiOTGUKAE75A6c
/Cge4RQLROW/mVH4xRBV+lBuiCyyOpWg+1PL9+fKoVwQjnix5ms+OOUhHoBXI0seLod+f3St1C0B
dARVzb5x5BAKN6Z3kND9YLVuceShNn3svoEWonsm/nBH0quaoUy5MUS8cQeGaazlv/EBqCxbS5jM
5esn1jifceX69H3xdsLxS3Rss7FjD+NPIL1l8Yf7prIorpzBrCjKu8NNbyCGy5X1gEKsJTkBCHyx
QhQxRKsZE3acPM/E5Qp2xqSaNdBHVvA/VvntD57nwXiTnA7JsN1dtTK2L5l6M1bWL/s+q7sURgAe
ZYqNYy2XEOLaKhlgX370Kb7T5Ej+Ll4YMNkp9XpEbakdK5cCoS2+cBaIjPCHnU921ipGn+bWRNxC
yFTaiLYM6GIVzTbe7SzJjh6KmjHQCIAgdAm0dgTBUt/B8Enw+h2QOInG17Xq4Rf9QUhsGuVL6Q82
V+JtRrbrAXc5Wj1F7j+n1ij7lapY4QUW7nfkueClqVhtEV1yeICozcKKsxxeCNgsNhDtgdwDp6X5
x2RtsWbZ3gJv7MVT2fUmn2XyhnfiRhiBdUhcXMeoq37VoPeCjhwEXC/aonIVi7wuvkYX5K/CAy61
yWr5bgqbo+AmxOBZDjwOM9FHSU9pEzYDfN6p+7nvtezeV6W7uNJP6ubv6qq77oNSMB161gZTmwyO
9nyFDYkXdcd7HIbxk0XwR5OnRKbnPhYSsppf+ONGUm+0osmLMbgdB26gOsf9vmFqm+lZqewJSLoC
nCi+1xJCI6dFTzXi1q4+wErPObU6wxDOl/F3Ln7TqRaqAs9ZPlaJXvl7TMA/iYqkMhsxJQ3Ht9bA
sqvpvPprflQkoiqit9gnqxr6pFM2kz+5quGvpGuYTbkTOOe31BZD0lEaYgPEnK4/K6hT9Q8QYzQY
O0j8uAwFH2+E0NyH7q47OMldPPo1QKFXWJxPjnAb0ci6ywVJQ9ZAENko+/QxTb+VFRcKtJot4mi5
Ku5D4tfThLGxBBHycilfFBfVOC9R02SSTxcRwguqJGTmXZ380TRNpb7sucqo/9UgiCc5unox/vg+
fKJB+5ltwrFquRDU9yHdkfybkY24v9ws54Ld2AtRMGyoqDL47J4vTPVFjvMHPr2cWsLXNYDqW0Kv
sBNSBjPoqEOTnPdY+rQs3/dq6q2j6E7TLXUKxBP7Z93ZtgeWvMSptkkGY6ZFT9DTttNev2JQqxxb
tZKZ1UvjToMbvwU5MHTulsWL396DiIRHKo5FIokMV29HjB5Op0XWfVlgkutZ4hF161ZhMFHp5Nh5
9h0qh1Wg03kpQyZuhbJETykfygDuDMZMA5GfVOCjkjUmNwAaHHdZfou5ukI/J50JYl7BRM576mpA
KUdJv9G5rP/9uBweevyq8nZ5cP9+k9TLkhT/j1uy3nopeauGMSCiWgNgXht8kmsPu1KUKZyiBjLA
g4ZZPkqzf90i5JZ09bDF6oQWKnh1MVKG2uhL/uLdYYGZCkJtmhD3TK8T3PCFYlYfJodEWgnTvjit
3P6xpkNKuepM3J3FNDpzu+3j/RIE8KMze/+OUI29E/1DvF9ZXeYeUDtcRSvgFLtHj+FRYiY9u+0l
op2v3P2eIQTaVAWr4wVYEtsmv0AtvwFFRG0pIUUId7cpFztJISlph2wQwEyZdTSbyCmAEpxgjp77
rqwzctkqvDSimZy+29zaFJRGGuPPXaWZ2wdC/mIWSJwSRPgn9hMqYbnlbqxues4km0sIMns0pQPS
i1vwjMgyANF7o4M1ljGkmGudQqwKSYaPDvht30PcuB1cI3i+Nj5K0q91B56q4kEUvs5AUyE85yd2
ckNasbjhxAORyl7EEw2K0tGwaokz43OSJ8SRLzAWCm2+IV9jOBG2996VkxZfktqbGqUIcWS2XZz1
gLGSu94EF2VQhBw9Clm+I0G1Xin4NKH68wvZyLYoLve6qH+GFlLXzZOjbu8huhUuQQOZc3i44LVT
eisdcCQhVe4YCa/nY6QxKI3nYkAi2uCGO4mmfzf4BwzhEx102GtDWY4oN2dWj4uEm1W39GaUXZA+
g7KqmIfeDFi8I6OsWKtiGmLdngJu26TERNFdtYXHT4DdauvtZX+o42G8S3Py/wHyuRR9TSXHEtME
CRE+ena/nCOkJ1joBuRxyj4+4xiYrRRDML/qqIygUtjFG20ba96WeF5n6xAgv598en2pbpboJIS1
0v8BNIn5qrxsEbET3pQX9QrGWyM3Sihi7psoIsIU07+PU+X61NNj70sSFZUdQWovXjGaN7Td2F7L
JiG6QLgW1il7pCGfJ0XHTRgQoz0Nl4P1Cnr3gbQB6jH4l/6VtNDrdgws5oxysNwOGslZbEY99khZ
q1g7aCpxIUHJQlk6Z8Jy3A77N/OERxQTuBZ5fJWqOovTS5/432sXmNY0MCAy+1ezU+yw1RBb2AVF
LZnA/M3YqyEnRfKmPaMSWbB7fNJdGoqM9fDjm9Pju5QiqFPH4LQkULcKCGew++7PSJo2XUzyPZ6c
eKPY4pS/j3JGVvn1lEAD/HVkx1nLV56eXyPxtJmCF4y8Z4CCNW/uyN86cLzbwiU0ygIxJS0nHUc/
M/Agz1lj/ME0c0eaP4bN9FsdsY2fWnL4X6KO/hTEuGGxohGDRsHf7nPr8oDg/yjrQU7WvUBmt8Vz
o4LzolEkjeCKiCvZQB2mD1mS7+xWzu5Wcqg+aywfCwUxCPpKwfkQqdt4np3bFCQGlKcjKhykaiGa
AIEtRqM0Iq5vwQPdjvsKK2GOa+uI2crptyQ7cN23kl1xjvt1cda1fgWSeRfl/+QxwJ3P5AspNEkV
z7hv0YENBF8eM+0WLJn1CevpPFjjidv37em4Qnu83nur4qk74KTSXW4ZwnIO/HP1+HusHr8E4fIp
ecnvoMYyHfMoh5M0Je+NnvK7Nn5YVacOz+9A7shXTPucs2NXVe6PfvrhJWcNyzow8F+Mi2EIG0P9
RnLBjOpIO775qHe1F63RU2YwgQz+uMIuF0bzQtoYlsOUBcV/K4I/YHlozGMcz12NzjLbuX6nfEIu
xFNSiU8s4eBQ/887UNAGtw8+gs7vFVc0V65JXtn8djy2690eiuXwLHsd/1c6HE10U/H5wgqawpME
DQ9weYu1Y5Tt0z5jwcRqVWgiCbM0v470V0Z+fY2qEhQgBs8PobXjqjZMyw8nQQ4PNkoLimLJ5daj
1uE66LrrwuOsF0VcXU66LPODHY6bOEMkQv6JaKAAZVcZHx94og77r4ffQGCjQ35wonqZFJa5mVRI
jGInsp08AIqk4xlRm/vKZAoN4OdHTS4gbZiD2r3GF5XV4Tu2x6oJ1yG3db7eX1YuGyKAGwFvJVXP
YrqyAIvcuAykYk8N/w88ACfH+aSf5RY7+Si1HAImrpG8DIc8KTama1KPp/gtk+4Oakx6+fuPVBr4
lm4kwSENARwkJ//9mIzztZahxhCG1XmbMXCmQ1f9NW3ytDJb29ud3xWVLSN2HCFqZOwwYysAkxFH
mKuTihEu7tNaUUkRQJsCSMdXi3/0jgMwWmw0rWbxAYNTZudQ1K2sYQpQ1JLeZslvI20humgBEiv4
QvlDsMSPBhSfP6+tYXlFPbncuHdl5M2VL0pnk9IIxsJOb7W77QqcTtvfuEcsxS7dFp5KcjWe2vc3
Nz83KT1ffhlhdSPgvxNc2/E0DcXNhFcM+RGB/lOMOx0kWAtpfJf8b/6MX1jaxBMc5lvGf/Gmd2S6
feeIdEqGq7eEH5o+ucT6xz7x+0Pjl0MqxJtaTwl1n1/aBZLZW4BoN50akFTzfZVfm6bhQ/8sVjNf
sE4MVWy89cOsb0woQHv3x7Z/RViwDF4DSYP9t97J11jnKmS6xZpL7L6TRKqWAAK+Xuz68iMp1gih
hjZ8k3b5w+R6fiLvxCqpzmU4yhpTXkdAoIvExgW3Ui4h3io53atT6weAl9sxBtPbLYqN63KA7gz6
XA937ld0yZGlbEb/iv7MjazVghm84YgeGGwEAWnseJ7nxO+Y0l6RkslbDF1fVEm/kgp/EA0k2Yn5
Cz6YKQpzg+uL3Ja2KOi+8P34IhAuJ3PdA7B/zEeXxxlpTl8KssKNUebRatDUw37VKE6teD28BHHN
GMuNub8SW9xBXXSDWK5Decugznz0q2JqIhBcNQ9XrVyaRbPjMQtfVSrpihV4/Fl5/04YKJIV08HL
UVsmBoZN/7U/gdqlfUDX1SGoEVKhRcCT14Rx/JWsocVuB8bZEVgRwOsAl7o1krOEfbdgCUPiF80I
zZOWLzP2SPZ73QD9sBk7su48WMKLAfc8PHAjr6CpvqUiIda4bAQQmxcGmEZJufWoG9VeAcJqdvlT
kGoSyESSU/ualsOH86VcqiqyIIqOQkqwdE0wwKZ/tPKIDIKeIKUNN+S+6ihXOz30s0P6lB5+/3oz
BWw9rmD6yvzGc3CyfGg7J8K61n4DcroZYBrVTz4f0LgmXJHkXCcyk2YC7eYJD1akQWsvnXm38ILK
ttX/ocFgUsLE0R6wYuWMScOZGC/kYuAdiG99hQx5sBYDeWREnC9pwgNI0AhIbFqyEkyF0hN9ekMr
rOpVL1j2NDQZCSpYK44aXrn9k2qwafQex5d3gHXlC5gg5fFvwPtEDYnfO5nJpaRxdVh/nsEYyCV3
4P7rQ7bY481Xe9+a+uNWy0/2zJGTJI8e5CnzPcS4VpxIrBCBjRvu+eKGExxZ8OciEug/Zf2+dfVA
zma8R87nTvnsbaFbrnhrPlh4EPwqrCUUb+br2xtRzO+dWkfwXEwmiI7NoiHzzLaionrEf/kFliOi
VdQuJFgwFzzEnUGpMKH1yVWjoAvcFovkesHINmEZjV5aOrhoS/w5Si038MF9nXf78I5j3tEcxdDi
fqb6nBztKh7oTK2SEXB+iVKZs2hzJS8UpgMbuo0MVWbCptpE9CSgRvBDZUbidS5FRKPrbjeXxsxC
CW7HOr6auXxGaOhdz6C+207fplnI0RlBkzrB9W732//SoYhG3TJ7POG3JomrnJIX9/o3tZWvhdT9
M0fy5AOO2QAzwhOBf7tRN+3tdV+jk8t450CA98pCx1VF00srkAFpH1hO1g+iYfXI0VRVIVDczeGS
CzibT8c0868y2JNvakYsZHm2ojrMMtisEyhaHMG3fiBnYZ0hFLbOvE3Vwu8APOzVdEM/GsbL7aLB
i7oBAkRJRe2C80uTg5IkDrTP0Cc/TaJp1VJlB+0AqLdm1rFusiBsNsfTe3n00xI4Ik/7Fy2oLBJh
gL9tDDo0MUfx26CuEKl7Q7Xh9NUXM9SbndF2rhw3obrxhRw7A4dA4Dj/+T0+1fBovuikQrZ3GQHh
8PkJWB5mkjYv/TaARpgbyMvEYK7KASGmovxfTcyAxRotGPvt9R+a/XiSwvRRjjbR7cTzD5c2HfXG
cZKKvJzyTqLLe5Bx7N/wydsK710ac9N60C3Dseh6wyyffJv8ZOX12zcvnsmkBZ7Hhp1Doo4sNWob
0lyvm4O/JUPV3HDmWEe1x5r72pKyWfVI0qQJi9cYH8/Dl70CPGyeHZ6HqkDB0f8XTZ5hC6NGFXNM
YEEegFgf9UHUQLlaQq2ssb4SlZ+zk3icrimwv4hvZUuWguw0r1fVQ65DmrI0ef4rVdMGM7heTA5c
ErQcR9M+/6zltZVxStKAjaD/IyMNIM/yO8qz+vbxfK3pimzIKpb4QnWZMJmnP1XKDUHxsF3wE7ON
PKgMmPglO/W6+d5GDSp+mNhVE/9gdkH1+saeGT0lG17th9TKR5jHDUXH7eWieA/K6gpRygqxe5/L
f2fbxNITCF80EtvfQzoUbkiyzFHa3RvHYmK1ypSxbKaK5SR1wRs6qEoIEuioKlbJce7DuKhvlWXJ
HBXJy9umjg8lJufcV7Up/rSYQgJzMzzzb1RNHc3TLwVuIz35NWHu81ZwnxhTxCzhNv8GGomR2sK4
uICTWxNKLGj8QePFAFQFE6b2npvHzpXkVfF+t3Rtr8Nv05Ury3Wmxyh1INMk/InD3Kg9lM7JiBm3
YV4b3LtD1vimflSbuQ7RmqVbJaHTnpqMcGbZMwK9pwe7A/nXVokqPeTZ3BQAkU/zKDx0scabISqw
oeHpf6svObYtLJsCGP0Fcn9Y9N+HM7nZlFFl35NfdO1AMLxnqp/kbQkq/4BFvx4TkIEJeGxeFI6p
UvbzSNXrE+T8R1+d2YYgWyr9ebGkGZ37sflhyVRdpdiKckKuy9tvzfbvtIJfrf0z9upn/jMpyq4F
KBxFcievZ9rXD/c4IqB3AdivZcfnKMZXdPHF9jCRNJH5z2tqzVR1lEOrqUwq+vvcjhMHdnBCrNIL
24vzqiyk48hjQ2QAk5FBYbnQe9RzgwBdBv9Y9EJZi+3YPmNmA1CwIpnurtl8Gc2xxD+a7jbPsKmo
QwnELrL5i4K1amhynGZhPXpkcyeVp2ZTQCM9HN9TfpJYBycmEPkesYdZSf4Py+t0Kd/x/4elLfbZ
hH6jRLtd/8ebyj1fdWLuKPJm3ZNPLX4HNnEE/EXn5SrjWTC+CRNSiBX5boivnOIwtWAy3WjdCkQM
56fZi++rxtKe2CG0LERz5zoaxLXrm+gJ1clbbVH77aA5tQrmjf/yK+2G917qhm7x/4R+Eb2f5mIN
99dzl498deikf/CzfDgaz6sbV4NFj+EBoR8RgoDDE7kEAoxl/VGz6cEhIhfvQE/5Kl0g61551cGt
8K51djoA5WGi1qTAIlkbZoU03TD3AgOIIGqTcR2XeOC1WvuEN8cOEvtBD1y9hIlUjXv7jVRfeV6L
1Q/3nI8U668AxBZywfIEf7wDV0QUtyEiPx7fiMEBUfABeMJD98enK6IsnxHYM9cNpnB5QVQp2mkh
SfuKJ5qKHg+eNvju5nCVMSL0dItLLroKBxm1/nPBl0jTZuBbzWjuYUXHar422sDEfK0mRDOACB3I
L1uSI50sRgmK+0jwlfMnhweY+DiTsLhycqo1Tvq42Yj7m8+XtO/IPcgcKMjQ3QgfCbwPuHlmuSMR
y0x22N7HEPR/0wWdmn4XgPzBtqLTYj463Q2ufh0LTtIHG8oe9AB9ML7E6fLeqg88D/8LASyWAJfU
aveG1p31O+3+bDym8mQB//eu3DhPlc4eal6KlHGoPHFgbx0XmQwoW1q4dJhyyaLf9oqpHdpGI9QT
KATfkVJCsjzUr2x87+Pczw3y0cgH5VayASxtVdduiFiycAEB4nn1+uTs1cNNE7/GogmqKLPxykqz
pAuvIoB4BQMkqlDm1UYbJoehVP6H9x5ig3bLti4Pxf9c4iLIkMfVr26I8hsiUkCCQT37+JiwdjJL
BY3pKClIb45jmwVJk/s9qSJOU9rJqDoa15fdTf2G6athMf7wn8s60Dc9N8A5EEtEKLJNo3sl2bgY
t+xSVCHi3YrimsTrhoEoFlZtkk4a/uAs/YPGWumgvW0iiimgAvYzzbtDG1Lt9qsf2QI4Gi3S1eYS
Ma+ekvCSJPxukmcgkDVEZwwAoTEoqbStl6tJQ5SMLGzj5ei0axrymsy5rNon3SXHhoO03qhibUCB
kFSjnsPWPbNNaujmvTkQ2T/ImE2eYXwxRV//0rK5DX3LlQKdxIITeBEC5neu0iQBNLFB1XiJsViS
T5TmYViNSl7hkBK8oAKq64C3hwTT5eqLoEZEFujRX2kvgrmblu5ncPGNRQtZlsGziILoitPtTTa3
hHRNQJilzlTQuxP2raEyz1Y4Rb6ZYYCiDP+FowIVoljaSl8KLvIXQyPPTnMTOiQ5oVb+wd9veUFe
x0nAe0ni4mqWlm4zxx8vheUDVvVVIMhdckXiIFz7+d2vzMf5hQS4XCHA9xvlpr9l5qXal4fliuBj
ChzFqaAl0zYVjSU7BLrjpyQOrwWjOTa5X5K9Z/AQv+MT0ADMTAY99x36MMt5vzBL7fxndjRHsM/B
guuJlqaamXug1tNGoUpfo7QpH3Fu+MW9fFoTtRJTOVxQmJWqtAz4KBf71o2B9GGVFSm7I7egWQmK
pwsm5miwod/dfTtxf6QWEXC0DmWUAz98jgIDQ719iYtYYUL1luM5hFNT8WdWvl0SyRtaJWwP6vSy
+AdUfZDsefmvbsDW9wnlLqqBg6Ua9PnTOh7lh3lvIAHnfZK3BJxBAoAhqNni13acE94XJlrlunyj
cEcZj1XIaDUf9p52HMd/FrUvJlGM+Lwn741RHMOpPTCybEY+HzPGzBQPWTaOyW0xbc70jqK8Z6EM
A9zZ5FdGu7mI6wWcG86SkqhA1QhW6q7YyU/w/pwU90KgLEAZoFaDI3HuqRiK97Xq4akDmV5g5sOL
1YLYLQOMsAdwf5+8sbdNk0TomnLuNuu6IscX6xYZt55lRjmwUtx2cERu2E1CCFyvbVkum5/WdHRE
3uMjea/ki7ENqa5DbNXhKIfwagsdkwj4Syzs+9NIhv/Dtg0RVYfDlsI+VsNR69o/ebyQU8FfRw7o
6wktlXYcO2ImJVdA5OTY5kfOQO+IsKjiqaFMIVPhfH4un4UnlzvWxrEDRTs0Eogb2CZSNqCbwA8D
4TtMOx6JZCe4/jeXFM0Kz04d6xk1+jQX0zbtATgQX4IquoVHXZ2BiaOLnSvSiQpNKV6PdcM45Aqq
FqSRZJPVUwG4cEf0T/d/CSSFk0FIYviSnhpgHwpH5uJ6XV2xdPGOiKqPhQXuuF1HUrXsUwIxlOui
/ZlBHI7OS1WfjILgg56pbGEicyHCHMDbG2ZfzQi/jhEZsC1LhjmMBd0+qZZ4dbUrfA4kxvOv4AGR
K7lwqrSdc16caJgghR6WL6MLJHlDgW5D+4SmK0D22FXNOUEtMMj9zuSjeuf6UE5+byDOk7fdrrKe
aOoFRnMCy30sK1u1V9QCd4P0o1cno8BNQP8HEPJvRDwhV8ls0lPEshLDWOQita3d3Ya+cdHh9iaS
XzH00cQ7rYy1Sq77irPKai15qOEyE1EYBneMDxuURHCYQw/lOhd6fjpmwh49DkqpXx8S4KpPaQtg
FcfgUh5oD2ioaFZEZ1QvaNVwM0mirARTNKTbHeP86p6wQ/82Ulz54s+BbA9HKw1T+MCPN5i5HXur
UifyCM996tQGbVn8GK142ibg/UZUYoYJELqJFHiwYvUOrUagzXRSRxfvG/q/2ykIlUtWMABtsMRl
km4cF1ipgcq1AxTHbSeZRg5aqQUDXbsKrfQz9fOIwOtzJR8WMSCyYkQLTYYrC6B5b7Epp2UzRNt4
IkpdqxW+nBZTef3YL2GnlE6tJT9eSLAZ7yXgKD3AvbGyqX1YsIXqQwf1owrqNWAbzOTnqG6Bhuu7
I4EfAODpzFXayOnDBd6dtAcP4cYXYZSSZHyCNW7j+VnYuXaa6pPrVGUIMtC+qEo2LK1jTHHjRiak
BPabvW4ulUXDEfY1kzElNvAWhQrAoc6/7C6/h7KzY6xsndbgjAAKJuDlvM7XfUlSgaBh66OQxSmp
YtQWJaJqBV7ImcQLKKZyuBbyyH859BoCUieLmxFzVogNIolms5Z40+3d/9GGmSSIBvhOID1rVSr1
YBRjPmVZlphbPMQEx4RBeMGVxUvDC4VVFJZZZ2QhTo9r0VuekN/lsOYjggoTmAmV/KEoHDgfqdRB
xTCModQTTOVJXPOttJUIrohhxFTz8UDOFuzlhXOuqbVjCf5dD+f5XdVqNapVZXcMvwM+QPOyRWlJ
tCGtFqCGd40JoEgyMlHkcM5Q4d+kEdq7hFbDzf6lWKKw602B5A2DSOR8dBkRor5N8Qjk0pJcG0Ds
xOZi1RFVLMjeDjvuK8Ug7Ko/fjwYTzJwRfKKN4PpKkM7RZFsar1Xq5Zn7qlsNkOYRmqYh9CQen9M
MeTqB7drV+9ujzhLVYn09U0YfHDUK2caknAfHtWST7D69AjTeI5qh8M9n6nKywTpu5CMjDBFxmsg
55iLzHiI6WYcG9IoAxC9mcVp5uO9xCEylYfc55eanlYChyAEcjAvTCF/LQrHVZ3YiJNfVCRoasXr
0y8co7TtJY03kcZ9ktxzq1PZ4glQWh3D5VDGXqzK1VfjcyGmTUYbALzhjc+CW59AcW94KXrKKAkJ
44sAtRRuOFAPCRwrpkCPpEI7bOK3AD7iRFdx6c9BPqJLPsuRNZNSTRNLyMv5ycD9q2xGcxhh6/wa
HHBAwfFBNhYlZLRFTqGf6gDmFZOTVUaXQDy3d5TDNDjbe65V4W0IuFO5WZOkYHdYwGZiRO3ocput
EY5HNYJCZPQxhHjaW3DII5qMPJv30IoERP4tCno0kvtQXONxehywguob2BKH1GjdJm59PDMAbL+b
wXI+48k6Vl7WG+THmcfXZ071n5LEkQpQCCPBuf6UrMU5/yy6mc4jQ+Ezqtaqfaf4hkGglw+yfJhP
pyqoD4xn/wNPt2JUJJEuQDJJ56xfweN2EJdNmb/1VCXw8ErgJNR7e4lKhTYOt/cXdeJm/9kqIaGY
SC+Npbv6fQiY8ekVBnZnkmglVyBt7I6Sgsp2vF1oCaaNMPezggynCCi8XXnlxczqQMYzmKP0PhAO
DUFDt2Kvrlpo41NcSPe6lP4YCkdzqXvmos49edYvu0U5sCxXgjANK0beYj6paLOkXBgRyHMP0QFp
xQ40DbxV8La5UzhHvFuYZWsEciHxlCWhia6RXVlMdyq1w/EfPzy5vbTZNcrZ6RVYGmFulQ7Xmx7H
iHTaDNiNrwLaFiXdXXGueFe7fgDZIwN3d3YwdL2j9lWYhxBUWZ/hAR/6lfO0cgcILCoDACO6B2iX
d67fMfnsdgjqV9ynjcpjuKCxZ19mb1ZH8bh+FdmgC85NXI2I+IIX1lL7XyRpmGj4aZk39WKZQ/q+
NDz06dNxcJ+RMLs/d+E0Dvq5CdVG/cu8M+gcQ2thhbyIC12kc/8xfThO1Nj7BqeWh+6cH79qHUht
9DX/YgZn1x9LFeV4ooYjNIhrxpR+5pyo3HGRcrxfOye855EGTNh9V9y3UDPUkKWqfWuYP1BaNGFn
X1yRj2X4Bta+tGG0gWBAmLRRhCnEj5wjvYAXltpRPgfb1CY8cQNEiDDT5zzgMBH9vz7gdx+7KxYp
TzgD/EXXG90ZAxBn2QpPAXfSROHoRx8ifliByvhh1GmOhlE6GdBzVRFgEpIPzAE0CLPzVBODkrvs
AtKRoyTiwYEg4i/+uXoQB1msbKHq7xEnKy89Zmkks8WmfaD2w+6n9cvRxoPNmTXxhB9ziADTpjvA
Dqb4p8il9UrsLBrTJ5jigVargD0CovlrrdWk0TqECtk/gdcXgv+x5f5r/eFf0ukVBWAQpU2xVJ39
AbaAFBdDhMrtp3kTDkae056/CNhQYYDi31SqsBcQ14uaBIXXDdw3shklTyuwT1tMbt4nhsm+TBkn
joIHJTdHRVGQe4XHzO34/flw7PbA8u9Ex0pHY7xyKooFYrGz7irI1ovYohaTkUGFqNge61AAZGNw
HZ6e26ThTsNfJ7JewP6OkHVJN/U1IB+yb40K96IVn8C53DU0XNJjISwe2tL0SVfarE+pi5P/jeMC
ZzngNtS6ui8KenQfhpueB5VSgejSEaw9JGrib0o9aVouhpqmHa/RP5Q+08184SypWiQZltFfVrB2
m7zGjQt1MKPFNzthUM6OiSX9EiDjSvu/qyV4vhEVwkSDD7LWmYNBVCTP5CjsdQSIh3mA890NOJP7
QX7GiKmBbaaFSKXl4o72E6g7uGH6SfojNY+mPAgj/1uMeghEarhYZkNyNTOoaoqpC22GR2vsezFM
MaY2wQXX1U9Ttj1BN7ZecmNMYoSVPQ167OyRDfyiPFHCKaqVi0ski8y8M6pYg000R1gol3caw/D1
b2tOHCQ5s1PiwJwN4V9z7FVHYUWOsnXoji/PmukVFESppEnCIEXBGSwsc+p1JawOKuX+asiEBtZ7
ZL+zf4WgSpOOQmVRcrYfbydVANZEkX2ZwJWxzovBcxIiaydy7JwEkjh/7HfUa3OSIFBleN3OQXJW
/FQzPfYBqyc0/QtNlAB+McJaCd34lSC4NeiAknNnOy3UiQXAM+iajyzhHblkTcW9Q8mi6L9dKJpI
onYfI9FqxK8dMH0aZrInuBqvaLqL4GO/kIj9mTZJZhatrOtdhmFN2qhV50CSBicduuGeMsUXhS+3
cKLSTJAIwKxaKAOKiUVoWKi7OaZ432ocJlvkY61triUft3QS1j5nglSJe+uU/p4WA41CqHQqtJjD
tu222man4H5YqZKlQtJb8Sw75bFssfQCoCPDDn0FL2+ctnMkoKChFGYXImN4HiadW8Oih6wWNMoz
NEkxDziFtoOKoXzOgOH94KmHCqU6Zg/6SG0lohSrmqW9Vm4mRSQ5oLlp8FRWWRJhmyDV/AnJN4Ew
N3dWIbQp1E8JFotQPgyNiW0mZ0lvDsgrW9smUA4zUwonKUM5aBgS/gvmlbil1HbAmMSCptm2yzih
d/MEwLghgTiOmEC2lgAqjbaGFh0u2qCEV27R08jQq5Erur8BPNpWosKkI9002FSSqmbXIUrCe1pc
8wMNBPoLYBKwFosGkz39Isx+p88nHSnAvDfBsgWRRDq1irtX/kZ06iSiegtljS/tqfEZhTizMvUp
kOVrkLpRDZ5shbQzeiHyDWMtAVFk7JjmNQ0dhwv/k9ZN3KJPLnBsV7CjjgrHzvLCh0/w2OJBDO8e
E/qYV1uuHfHrAL6POfpQFwyAdH/r8xMZZmD+9dbkHh+DxFRcD7s22nioITudIOjGY4RaQ3XkUHjw
WTj2XpMwCVeV019LI7JA7gCWqk1EPD9xobhQKO6IoOxOo5VOCInk43iqUdzZlij65h3EVjWZb14J
IIgGCGhpb0uSljIgVndqisR+HnlU2rkbSFnBEVLDkC2iO8iFwzOZYS+zJHXPVWLaLfbTd9ZzyKlQ
wJs1VJgr70lZ29vvXze49CenUQ93/cFB6bsk3smcNdB2Bt+KWbUEYEwp3cbAjz7Z8hu6B+8jfvXU
WIlzmRYReoq2YrmEVenGXpTqRavVXaeUDH0ZT0XKB2BYUnDFPlPYHq7uH2PLgbwLll9dqygGrAbk
ekTcKjjNeFkPOAI7jGUJhg9+vrLCQU9+20qs0sgeNnZT1HQM/iDNDFbkuS23qi5QqXYTNV1cVWgN
rmpmbmZfAPhXwfg5qufd4FyRkNLrWA9tGJvVyjpIPmX54mPKVz/aiJRfcJuQr/U/j+HMn+0zA4ev
xo/wtq9Qr12nO3GOdF7A5bRuGjQ1v17Vm7l/ukAnLdExF/fqgToMLgt9CrMCtxmnWN0fP4BN9J8T
l7mHbpy12SrkqI9nplGJvMcS5tmr0RPAgHJAVjkTBuL4dD+ez3d4BMYBoEFc0x8K3ReR1JDRfSVJ
ya1kaV8Pgichz9zJu8BD3lOKzCl6rgyFu2/+K8QFaPeymSP8bbUixxOL2iEndYoAOVqpTdaqCz+r
2ND6I10v+DMEBPrxykPNGJhUd/UxA6zbtaPWjxBedaYV7wo5/TEiEQ9B5pBXNKFYdM1/P7gpS+FG
3Ta/+nPLvcRdjzudBhIMNQZR+V0MTDAo0bNw/wO71dCfQnd+tBtxcYMDOpBPIPTmgFzwIklbjA9f
z73zrNJaJ0P12de4qSgEQ8xarGBDvYh7yrfaVa/rosrfOFhw2IUMnf9gQ+KX9n+AxbnwP/V6pgsn
kNJ/ius0gsUHzrSmo86a/oKaK8YOYMAjE8gNtMXlMdalmRkOtm37tCup83LmSM7GWjrMtzbE+oIw
wAD3DfobqFg9dw9H+u05ub3ef94ysoPnW1nIn59ETjpQRbA4NWV2KRlOROvdoPFjCb9QYr+SdIHr
3Ll+l1SWmuUNGvEDDT4kXda6/OKVXSY6AQFZoELARUjUj7SFSaDVR3DFFWCNulnqvrjglAFhTeUk
u6tt2SapOHYhlYtOLX3Bq52SQsusmfpHqw0+qtuf8uIp9Ql8MRHgu8xiyWdNVAfJ6HoNduJZDSE+
WB+mmEmKi5+0vkW/YFJbnIoJ0B3qcVvVLB0+LZMKe52hllbL7GT0fzrcsEqDWzsJ+EtyvJHH5x08
d0ScYEf8sUkDEtwnTDGSI0QuEV5CHbbgaD72c75Tdu0dQK67o+FHx9kFH5Ty+Bk2iyvSYt6u0EHZ
OAG5qQ02mNJgJyVclh8wuIvBv9GRSrtYMptNamW+JZDEdInz/kccX6ywEqemJh6GvdfkmHj0l3PQ
saDmI3xvc/PDVvPxB/OdPaEzMMlLMban6CRo131qyV7eQMTjd3TAdaDz1FiaNpajmNCCCT70FvAl
ACdu1fGjo3dHGCcpbgcd6o+psfcira9MMUbxF+IRv2WE9W1KM35/TKBMDqykVROJXJzEKGf9VVos
TVGd0iSBkAnXI5URE3tCU/GUCMfRc/BevMDtaKX3fk9oVYkdlRGGlxEx8P2uehWF6RqK0Oh8QPtR
uI0NiyIeHzoLrbelQnN/Glr3KiKwjgHdz/MB9RSx3HvksjXoKgwOqHPAVGZ1457wYUqG+RBz8y+P
xWB7Ef7Ds4mVpIiPMRxLfYEhiW/RriwGog1oBV0Hs+L7i4MjbvUQvfZIRpBPTt3FjNJwsQySAmxO
h9TYQhqbH3UJXHhJj4gfgq3bDY90Kw9EwkjhuVSg3DUwOqv3kxpPNdPmAK3Kv19F8qBCzsdArSvr
mlKOVt0ZIVH7RSi0qsT/hGg/EL5HyV4sg5l0SXThOuk2sUss6oPQTrpDrdPreVq0MS+keDtMdDid
MaJSbKopgwVbiOmP1zSss3KbvbTzEEs8dA+RXAdTa8FVCp/pKuFrMphrZw3BMezHkAPkeu3PCTAa
XOVpsbbDgelr+Zsl2oSo9ZzYllflQ2lHYxIFFABV2mVpJGhlmClvNNFrNVziSFyGsg1VHU9SA7vU
6LB7mpoWQtA/EJuIc1DG6tZHP7JJhO7yKOqkwwYyJMIz6eVKi9asrHdAkgbvKxFv4KZk66kvGz8O
ogV/5ny5ow1ABFEUVs8hwQcDEWnVFGfCY4vkZuLvhIgzNZqY3sZUurx3Jg6Smh/RmXTXJ82FPUTn
eILLuGSaoqOAvLFiE0G27irCjql6eyhoN2sZeSH5nnNQtasUFgb9sPi3myl9iw91GAzAErySKGuW
sSISVY03rxBK7vYGPGSsFlpgJWzaVfn8NJK5ca2I2rFd3rBKjZpFTWOEMksEiGDqf06o49OrZl/x
3tNU48P+sPm1zDlOVluKOo2XOXWcXfvh3u0drRV9C/yUVGeoCpYJzeNz3XQC4fKcte3wvfJx40z9
QHBunLxShog12d0uAoI1rppgtMJXBP6jPEfmkjOkT1SHgiAMLbPccjXoEuuIUiyrRZBDiSG7n5E+
oCc2jnt9VX+xz2di+Q7yXKcoBbJTj/9va7Df4Mz/XukHPnYClGU4aVBEtbWdAFVaxD/LOzBiXWwE
ON45AEeIEkhTzF2DPhAC6I3vu9oDIqG9pxOKauzjhsQSkBMYVVgaBhiuCsPtwq/hxq5opmJqfOeS
Fwtql2s6K2Gaep4Mgo7XVZfjvomHrO8pBDWFxcDcoxmnDn4SIV9Lgc5LTg+3hv18X1UtfdtLDTKz
d03mtQiL+bNK0Qq4seFTg+Iz9EqQVxgUZXjLQ2Qh7Zoyh2aVlyxMqLjovdX1u/JKJw3AXbJbi0oo
y8drc3hotBy0BX57A7TK+6FvvwzyjyAFGPROHQuiTHv6iomrtKIhFHbM0uHJZ16JKi/QTMBTTA8Y
qQGWmiLe5lmIySkLurKWwtSUhvls4JPurV9IVXXOnt2K15iaKCKL3/iUwSbXcZIiniDHMGGbTKvq
jhErskeMf+UFOD7h70n+UFH43p6vTFz2uw7PvKX8/NB+JuViTulfKxWR9o+fqNhoYacV8c06ektr
gQplqXJDJToJiVOO6893HYP3q0JOxXxhcfuyDKmuDNwsIoQOuiyiR8kgbdlJn8nlAq7DXTPBMCAG
JlbrOq5QFfyNG1Tdnd+n0ZJBS2E6sb98IiT1u73pDQgMcJ9kx21sHpNXdPIE8/m7tRp0UL9oT//e
CXZ8J4KbQEOb/EENeR2slGcTnP9XdDq+6VOxpyESPzVsMFdP3YmGlBGkpUGxGc6E5/sHT+IyOU70
aiiNDfPkoVqEq75p0nJhgldPmCUgVGl935vCow18+CqcfuZf8XnHS108lQwVQc3XOn+r2VkJTbMp
y58py5Iv3VnYqEuGpHi9KXjdJzTlqGjMsFfY8A1fHg67ALIpWglFnsRAh6y9QR1PPkBci8dmHILY
OQpx4pKow+FsOLlv11aiJP+zDo1Gw+/EVXGXu+asX9ghrw6McmJWzIMJQzYeXxAZj53c9DWPjiXr
CjUXnjIY+lA3/5mFRsLlQKbVcxniIQe8zbQ4TcDgjGM8ES5p/uGU+Hp0Vv5FOosbTwYfNFWkZdUZ
dQigCnYzxbZht/hnkBzpM8vdflQMrt7m4Syo2frxuOFKQBmFKB28xSrzHZiQ8wRDRoMmnV9N416C
UF4HEjVL8FtziHFBCwslDf5G5S1I6QsrvYJwXswchg74H1XJqJU8REnsNicFQQIh6LUNuOsV8+EA
XH/IwCoSc096hmGIRq3uDd5rQmkD+xkARZrscjCgOXxXtrC5/dfw47ei1JPk0MppMQKOJ7oXxan2
9fGfyShUOUdxyYwe17N2YAFKSDc4yWcYY8uyOPEP3oGMpCeEqdb9ffJvP958yIi4KD7cPF9U8Yt7
+a3h6WwM5oi/v3Eoj1vHvHfRYvnS5FYxnYxHSdhXR4Z8JZ4L7cbjr4D0aBzZTq5GceWfSe5NXs6s
ketnehLKXpZ/IAmrwshvlleLQBP4Ye32ywrZciN9RyxgdOVDowJxdl5zvEMBscntHVVCK+pvlGe8
qkzN4esOhbMMC7qodcvD/4cMB+QbdjiA04ajtNN/dqNwpUSu9EclVuXcU+IG6s7nCUzCEy3OmVg0
7X3p80xmYNYnV5/nQlVu3XjowYGTolqVNYMIGdWCsUGVzM9DSBndjL1iP9cLCVAIY1Mkw4mM/+hY
dY73Zm6o//e1+ab57S+sCnYfr7tdtybjd3oQmbQ0BXXSBdWpZq8PDSN2vJOq+4ENlM5EESEZVPCt
HKmCsDiwYNbTVrkVODlBuRt9QD4iNFz2wBwO+PSEKV1TIrew14DM/daYzMaFbTQQgVKwftAr/Dzu
Ftce/UOAPCPGStrN5xxH7pKWFnjsgmcgllV7K9uiKvLhH7b52d08dXZIESAUlCoG1+PjCcGoc5CO
9mV5LgQm7HJZgD1fe+5462R1zC4RB5XkdbRnPUELFobcbXcKpW+bpvFQFjS3I9hQ9a3lHcCSakSi
uBvnvR+O2QIHTa34n0+0b+54x5dArr1rjpXz6P7uIRhGkIxk0pTXE9/6C8TlN2rCKk3LcxykVaXi
PY+qSkD4biU56qYxKyaM4sRabGGYi8o1tp3/dUNihN3XLXXhAhtr6fWpfuIlEZtHzUq4x0X5dObw
dNU6ISaJmbJxaMYQWgkIMKd7qQt9lVmlYrFne8gIyXP//57us0SoA66vOqcFSI5dXVcKdcYtIy7t
UDghmTpT7yPJysVzOyvZtW7JTqFNmJ4CXalIJC7cA8IVjn72SZjc1ugA6+l0QYV58Tvm/Lea3Wd8
96XvAAIs93QDVd1XqCHGmpSy+xtnPT8+R4vkCsZHEfxQErTyys/goOVo7jiOssI9vuwVSywoBUGl
9PZp0eBhhbYNMe8qvdR0EU/UhR6yW7zplnk01je6WkldhwETrDLYjWy/XZtf4i1kSDVy/VaTivLH
BZGUYU6ZA7bBUh4Xvv5GGta7zWW4UlF9oXTBh6t34ACujIc+RfpYSmV2yR/Ey/CyPDmu7koKl+Vt
LOY6UCO3TxzuJeJIxeO00+8hMNiO7GGbDrg0hrfjwMXLq8NFWcv2XtNlNcdZixHE9heLVMdUGzo1
P4CN0NtNlPlTWvv2zXfOjPTd4FS96uaJHkRz39KoFKSMM8xS8SJ1c98pB2ipzxkXnGy6VpZ26a0I
zi12A8LKOyQmcZZqgxcHztqDcdOvOeOZD4LcZMYTXGKVdR5WGvKfH7dcQlQLoCypSpV2/qrNV6a6
TreCf91BOyx+xj5wK7EoMnZwlXItmz1jeV3csOtKkpo+/sxLX4sWuHgr88FIfAD0CCIPdL3UqbM1
tb8/Z+qpE/4zLZdmLoNgLhHiuKE5oO25iQ99CFzqKnKat7zWN+dKrRg3o/1u5sN/SOwqyLBMUCi3
eMsH7HwWi8ePqsnm586Y2tW6OtjUBxQxL2yBo2pLE3zv7ftYv/NetBrvh5mu9oJncV88PCMP06BD
Wdu+uQ6FsoNVcwVN8us85IEHwt7cxx2Yaoj22Qq+oQ0AeKkP3Zs/L9bIdHuFVewJwAgaIhPysXt6
og5OVPSwhVH/caJSej1eF1Z2THx877eVyK+4s7hsNNFrqlz7YP9iFZ911WUImdwMoLIOpGbPdEqV
HtgNIe/OxtX7G/BjQLyXxEytacDANw1ggelC+yd1XQPj2lkkxAhIHgUBBWkRaSs1hThwpsg0W8cL
yvjiiRaZB+7b1EhbDMcIa5iuDhC2SiCLrR6jzXDRO6bsAT75hCXAoEOeMzPZ7w6IqFnKqD7zy4aa
0AKTcsDym9eetFBJqolqxZK6pTwX11fKr8Db0t/CUEsQjTMNwfAluANTCP7kLoj9IOqr/jy9tmcE
I6YbmaQ1UAXkpsPr71GgetO+cTEwkm6y4PR+4KHBnhB1Bv0k6uiUj3dy1CSm84FYDBxf+/iydyJB
j6gY812yWiHANLzKaT0vnEQrGnF+WsQ0KoHRLFrRUm+2BO0p1p9GdCrzoOpdL/aTg95cgtQDb4AX
dOSPi4Y/xykGLhQnHOOvx8MI4v+k7RMxVPsc9n7z9vONlWScBxzURaR9bxbzxY59IABZdU9mhBXc
SSLhvWhX9AddDQnj/TjT0z4OwxtBLIzTMRDSjhy1ctgSDLREEisRXed284Jkj+Z9q/LAHnM5TmIj
Jsb//a/57NzyGDk+L1cW8qKBzxf9blPbpD/nG/XQDPELQqivqjSCD37U64FQQ2GbMDVCCu0e3DNS
l8kARTpp9rpWCYafcGL/DumlkRXbjj2EuVM908dPksn1mNTvrA5mr+3MhMe38UcdZateoAKY1BYv
EUhe7SAx1DDv4fQsw3cuEHQNmD/dAFrVdJK0gUoN37yUWadB9x6w4a2rQYPG5Cn9gqgNNPbLJL6B
wIFEF2ZhdNJooOZfs7052YpySOJH+CSIDjPm8UoJDy9pB7dUOtrWpGamcVuJ09Vcn0P6MzLy91qu
3moPngxqJ9ACHdjLk7E2PI5M0VqrabrzGXq+04t6U1yCsuUBfWzvsFjY0WasebCBqN8HhkkQpOSH
kYcyMqXIfbQU3Msn9DLNRPXEnHxVZ5ELcrpa06+drn6pa22juIsC+QPfE63uL9HPxRHFfMaG/niB
rbkT9RAoZjRnwxzUFgMP0j/OIBp5mKDlp18DOQR6jkxR62A4CgFkGy/zGNN5ggfuJ9LHcryD6NE/
rrYNqJaPz2ejX2s51ijWO7Y6RXuOZd6HvDzBSkjjT4Cz2z1ig2s3UUzlfi8whMwH5hMN8bAbnyjo
XlnKZjMUshfxcSz19CdIu2Ei5Kck0CMC1zlQUSsNebWklnt2Zl6JLkfV7Ar5/NbBY8A/jdvnCVE5
hSP90WsSfwqqKYLshyNIzQrZgly8OJzaXxtefMXEPpijxoABWKjMoxJUU0oS0ovG95tsYoxGTCVD
pLwIf4aYAX5gTK+7HkciDQcHENqVWFC0GeCQXa/3wV3r/hAmr7i2WPUyxol3shpiC8r9Hk639FkD
agzvVvxS+sLTG9BuscTEAJXjaTfLWo8Vqz6QMkW2rPoaLPNjCettGcrOzbNeA0JsDtd14KrpFkg/
VQrzE/FWHYKTXwz/QRedp1qqI5O+94FDjJ/rdGOGBJD8bWstjvNUkxKrW4LP7dYYw//Ot9mpP3sW
NrUvwh8x63Lmkx/PY46zIR/yKuN+OcvDEZMxt3EE6FhlLf7JKzWapBhqFiSdd1aq8es4dZRZ2ZgW
svOekMmJZoRilzK4YCo++Cop6VBpOikXp3udEQL7PDsV6ycB/NnBn8wTVOoDbedrG3eJX7DlxiiM
TOSV6xaYbX+OVHqLZ46xkGIb9RMY2iXVLcXSBlejdz9y7N8rSDYZyX0E6b8OrRK61vV/bTglJ7Y+
E8C3yh8vzQ01/vza33sTWRr5ffZ+q5BoJ3AAMUlOXr9m5qOM092WTphInv+VYyrIuDcCrMOt/d5y
EWKfB3EJiyCI23SDfKVv+BFwpnwJZcB6GdYjFYcs8iUunmG7pFxklCBPZBpvUjDjJKZRokZOW0yf
50CrGYKySqx/vLEJ1Gf56lWk5piAkEbOXoYiu+LDs18nUZ7Hbz+jpmw6AEmVdiBjFcguibRT8kqi
XXhA4Tc/A3CvNW1nINo8GwWre4Gq486qicuKJlie+rwM6PPkS/jJMK3lCXu4PY1NAXX5MQRgtspC
A9H2SuawqFAs+W8rLK3Mg1Xxuwqzk4qhtRbbt6PRHqHRHweCSfIxJF03/0uLwWPrRj6jOs7wOMRW
058bQls0xuVoBQmroGBgKYgoYvdyVYGtJUm2oCnwyAPqxYfXRusZMnyC39z6NUSSToB6yLrzzp8w
itFC3nfmb4resS8myiYP+UtT760VqKSlJ+nhT6Nv6qynUDIjwWNA9XHcf8GraxB3/RtNQkMsIZ5f
vdTSiFRMjYWprc0HYtVf4zNkUoxM1MCUteeD5OwyU+alyhFkclyP3oDlEg/03IXfuHFbl3GJgLm/
pBXarcszo4dinFNFsabEGP5CjVsk19ltaH0na+/1Fo9je171SoQssvGBbpt5iHqAEj+SIPlU9thy
Adw+LoyEr+AJTzdwKATaXrlkDfzdfeC7lOXmQ2WXCOviKL9cqxi99jximzJfzy4jQITsCVEZG6Vy
vLmuDrYSJ5CRyl2YUbqH1alp66xlJizvvnVZQYHU+2c5sq+epxDYRyD2wCVFSYB+rPHMGwCZnbom
xa/7sn1EmtGJiBY2vwDanXeqK2liq79TpJY09UFLYoNcemQiRlC1mqfwcfNxThl+xildnSFbEdHN
ZF6JzVS2HvV8pYa2YqzuoN6Hpiy6wqdlb9wB9m0+S7EgxvTFeeM+k6ADWuimffp8H90bBEBJJ43v
9iCrqfV9W3G01/Yfm8cHl2s0ZEXDkm1Q6fwUj6tQnvmPS3L2J4H+Whiwzv9f4oh7iurmp8K9lCge
UYU7GZEj8l5BVtpHlz74F3ChhOh1hH8Igw3XjMk6N7Nifv96kN/erxPmdAl5H8Z2aUq3RbXc56Ay
TQ5aie7mYV4CCx1xwmMVxmFG06NJN1IiB9mLSwgPqaR7Lg9ps/uutOol0NsYPBaurIZ7AqtrUk8c
A80kW81+xZShl+SCXXhjsKerI+1lFagr/D2RpnwrYInHZwWfTn3p8B7E+dG/FDJkn6rDrwykecDl
UacjgvcrhX23S1XfQ4hGjV7CYD8BOz/wGyhuG3yhfliv5YdWHCBWiofpXU9smwstLVpSJqOYI7jx
/xq9ciF64gmLz/3x1eMc5NnwbMjaclCNb/dAfoECu8zJuhVK2OjqWu2BJa/bUaYwZI1V7Eq01B9P
LuQUGCMJ+vjQJIpqbpGffHOK0wGCfFV8j00xiXsdcAhGleNjOBz3TyKBTn7d9fa+fGrSOY3IKJXN
GrJCbJPkspv9cvp7eCrukqKYyvappD7SEnMS/WhXDp7hsHDqQz1UKxDZDGStmVsk+z01oaT1LC2X
oYnOyfkKzHL7h1Fh25VlDuHK65dO5dw2o1okcbEO52bAl91u1kDMhNB2LvWzSAEZv7tyd+7N13Dc
RSU+A9RzOGUrR3zYXMGKcl53WA0zcFtVuKzVK3M9hmYqRFwBHTxRZOZzK0aai+SMpOxw7WmLVpI6
MHm28b/1oXlaJ1ggfHnOgl9OxEvvgFMhEIZ+B7u1A8vGWtGplERyjLMtp9xgZ+aKsdPD9UWMK0fa
nzIcQ+twI52Lu25ZEEKDHIVXrEjQquoUuygLiTZTVKNBy5BLjThhGsD4zdFEVrV9SZNWc9sa0Fo5
jRiSV8umv8methKSrK7GJaAG3t9jwLMOQD63lS+ZHRhJxEQUwkf2pWugeoypJrccTFP04S3gpJUO
YjlJ4miTT1sGENSeoFDfIRilFOKcZXlnCC/2TodXqMHg+7nfxlpHNBazkHJAQufdN9OAl08kaVdk
zdkTsx7luv2ykDoQtCNucVPr8DsVhH9g4AMmIgjC1HWq0bXD726bBtj6+bBapARsF/ClzcUBYgV9
QjWIMNt1VdHQrNdvq8tcUToVJkH2zVwTecFwpsQb6rcXdkEKXwu/qVALI0sAk4rNRk0GKHOAF43N
jP1ONI0WqTiGUYS+w4snEqN1jnYPNMUm/VP2BK0M6ANrjC0/IrJqbP3sGH4jVrth0jYCcZ9KFmpG
xTTV/MTcYlcwxNAJf9FcTnY4vEb+fboZCUC12hXyF933bgkLogoIbZDpxDyT7G5eINkctKbbh9bu
QIX2RVUYZlTpJPUGyEQh1hqGBApW+lOdAdhgqzqW+3WsPtx/WlkVE0Qd21H8s48uU+BWjY2SRo41
ZiMD8QR7r8LwOhmTjPWQbCToVH8Oj/XNJaoSxfyLV7VHZ2rZ0sfl+A+R5gF67X7vIwsXhcLXkZaZ
Q16/2e/vavmNhBJBkcbTC2gav3n6dpaRM1v0jAfY+ObV6VOVywfYdVKmtTsZ1XMm1PsQ+oopPQtW
aNrrABAV8ud1KciEp0gyGfKBkJiZz1R6k5onFiPNX3/23CnTM2yAkVEbJpD016OFoCyCAosdEQCs
wwTZ3yowCNMxkXs0XSfULBuM31Jtdw3ThoMD676uHOnntnAzPD4L66GBo2y7NKd9fM9K7nQZxn99
2nSzB/Onh2tIBYAB/qYRhHO1Ad+W6QepfRRy72Utci8hSWArdlDJ/Ib/VmYM9VcAUrRl9YUh3LN4
gGIm4yYdXm+9KA/VLWDBW13x6bIyNhMD860vKUWLuoW9M8PMyEWGrT42UtgQoX4QPcqcigkvj7b9
vbWXxUFvY0v6YhMiD0lhjvyRgZ1V9kuh1unafF5WgMpG3bZQWh4aBpR/5ISP7K1MZ1z1G7zfgIUq
tRp9g/Jh5/BkGVQ3Knu4mcGSJwkCBVyqVGbijsQTlJMAyUxRys1/cqwT0QDyE4pnTpsa+E67pPbD
ZJojPWQeSKnTM7+Bi2/OWP7FUjWN/BwP3tmE9n6D2EIbG0hRQPXcin/BCJypeN7fhCILtGBdONsu
T2+ynmPfdh0G0RBvKkCtOh6DhKQs7Sx7EToS2X4tXOWnZMQuI+9XoyJMZ0vk88QhKFC0JlVNv8Cl
QjAkha68LngV5w/iviBd2LDn0R6SOqAnKsB/wvDZeOgFCYFu8DXjSLjXDH8Tdk3SIsuujQ8C5sla
8rIV5XQ3Ma7oKlHz/rcBKP5F6qBn95HVjy1Uy23zDB1mbtfzc8oiRVdBiB1fmQWc5GIWtIiwC+XB
JqWhfBDQKOKmL6vryaa0H1xbaRzfWCuRld1/h4ZvvW5et7e9wRIk0hqOq7gYlijhUTZXlGKutiNM
L5LSzC/a9g1Ir8WAWbKoh/PifRHzwldSgPGRwR8QY+LhOLv0bRNtrFcmXINNxqtVbk4greAcjk+A
zKy/giYSYQRcAoyhnqR7/BH3JpWfVz2ybniEb2x3mzZt0GudU9hKH6QtIOXj92nChhgYRFvTQPlh
IwCeG7H9atWI27eKDCVS74g/vWFtYK07DqyIrmdIQ+9niVXT1UG5j49iawH0mKHjRVtvRnl9EFd0
GX9DRbgko6uS8GCnx/oqjL2Z0ptrE+M+JO5FVqK02EtSKaFZ+zu7drmbGaQb7kBb+schxk3/3ixj
WjlxvV1rtOfGYOp72BR83q83dvAMF0Z47LWRyWQccsu7+xb5lXA9YilzIqct7VuN1XPoJSx49Ina
/O4egB9pQn9VGyGhuyOAdJ6jiDUVEhF8dJnFXcVuh+Q5jcRciwJi7C0pk0qO6JkhH6SqXrsSYhX1
VrWKR0QbTKiAMah+iMj9gD7xr+PrtwAmslgKiFTfbDmaYu9r2fAu6HXThUIA3efKhma3MmKZEhmp
CHtcMy/a8ClfvlhAAv79tQDTyKgEVyv9KHNE2BaVXKnv4o59XHHo4Rxj7qZE0daZS24jrDel8FzV
DJyu8rv9PONxJnHeg814LSTGLxN2LP6Ud5ia33sc+gaFmlgZEB5ZiPe7abEgObW2ninC4mEMpN8V
oukK/Q6j+h/jgE5t0+5PIA8HhW+uZzLXAt5ph2w4jEKQWEmP0qSZ+Yv3CWY8teI/2B9EXcFgbsy8
dxtXveZaT5nDiSBCUger0TYNuXZtPXhSAeji2rWssBJS7dIp3OPoYSeTG5dlrMFdEqXOa9B3b6eg
yHTb38Mk8i9mX3IBcphd9A/ZgfNKVvy0DRSJSfGNFOGA4PxhqOUHCeXhwzy+0VF+mCbU8MCAJZmg
SZHdOCJCh9WV4b9fB6XD3uJA7QpSifPvWhgpikado+q305TPnbdDXk1FB1cONuqMcyZcuKwAqRbr
dPjb7ebiTX43b66UfcXrupBrWzBL23uBz9SAf4EYFK40yf85+H732niU3sxBoSx9S3YP8GTBIZFD
ZojbSHujTiG4fxGnVesRQbfs7kb5Wcu35XmZMxzu/JA9Hr/qJ5VclSNYqWd++pKrhC1z6HlCXy6Z
zmMw5Rh6Zr2IpqROjgQT9PI9JMV7FvdEhdGEp9LOpAmuOYON5MrT5cEkmF+Aes6xG4qJ2Yu03T9P
IqC3nKwzHOarttlZFIhMZnIQf5zEyjd2AOmASejiWLX5lOeLcicqEjbtQhXQHtiw+Bu5ggFo33QK
q/tGwrEF/URu8zfXG2Bca4QH+8rn1QmQVDd60zCahDE9jRh/E7Q2ObTxW2ib/y5AMAoOOg3jITtK
0XrUaqOGq0Yuq2ZtnjY9tfvS5ps7Fx8zQlBvSAkDN3V1pgUNXfq1UFjC31JOXA+4ig5DcVVdUAB4
uZ43kQYfDF/9hF9lU9ftgsnz444Cn1ZrfqjR3b5RqkXI15HTs0GWp0rLNnfUa7EY5IsSuNH9fM1H
kqtLeUTJNSqNKmOjIWHKl7TTi5f6bNhyJWMjx1phzqQQNuzCutrUnpxUFhpXYau/FwWviw5FAwpx
VLxJ0oRYYFe/AM7afdgU8sq0/n75Tu3vNp9YXckuMPUy24LbuY+gOMrMS7Q4lYo3f69ExZOhMKb3
j7IgNFSslMM6mKGI/qceitaITq1XwcvHhPPnqBt2lhMoBVduiLNaAzFo4OEJtCMnUcDnh3b/v1ro
YgiqNB9W23gDuf8fMKqe2hJ52f+W4+S9AVGNjH+Rju0rTr18ME7eW9OBhpyLfJZA81SXIrINmSVh
GVV8TgJvWHfBCJYZAJl1hBv8EIwEgajk+xX1g8b69l1XCQlVjvxkIesF1sB3bgBv9xAsLBaGGsTT
f47i8UaAvK5QlSBkblOZc0nMXyOyAw/UXYxSdykNlp18sB7Da7f4BBxHf9+iKbQaTnBB0g5SLGNT
P3eFmp/MuaEv1nVQCmQ8BGt14njm/rBeL9iHWeq/2iJMcCk+kv2a/hKf/uj6+AlytSbKVq9fIR+M
SNDjqK3dwqkInSuZJRcuiX9bwezclJn2UAAb70bLyiPSDJeLWFhjfciic4Qy0jOc6OL+FSU5ZQFA
niyehpAwQlklrbwca5MPVwssQdkjKVai9HcXfUD8oucNEWuoVq566H7nPEdBqIkCMdTjwcTQAXvw
iScotDWHau0gBiKi9Xvd1AbxM81SynYM98OMfg7om1XYkKoivanWIDezwrgV5II0jTO8MwS4CchS
aKRtzsxWtyideePTwm7fG32kbsEWzJm4JLNlo3sP//qBnx9V4GdniCkZMciLkjKX5apvf92cv4Gu
fWLRGLYpOlyJ1RBjGqiU7gmrwvqPqF4or39JUoX7AjAY9P/+yl3HXPldFGiqMOilYwnxdAZPwEnu
QLFTwhtoCw8pb6G7vk7shIZfHGcQUUjnaYuNfpsL5FGX5sXZcusmyO2Hwkx4+OhnOkWYtTYiHFQj
2E4E2ddAxgb1iEs2zS4uYXc8vu/OGCfMs99OMO9OY5jmXgVevKz0CyRpXkS9Bkk79bxYtddxUNnZ
JCi1R05JrVopKgfW7GQvScsS/6FalzhAcM8fG2DnjHgtP1rHLWXplGDVgUeWzBhrUXvYuRTXPrth
tFCrmCLUVhSj9Lwx1uu9Qj3J013veAwwiql3W7rMDzBNPB6XwkYraKYoETPVDf5V6nmPn6fGx4NT
2EwHVImx1fFV/1PER96+hu3y8tceFjrTtVNoSeJi5tH3UUHkPxGFJ3onEBTjORQ4PrsqU44o1lC7
xvvuQ77eEbFHTZNsDnwcR4uK/r0CVF673wb3Em65WwB/Iq20rMrgOuY0WMhVGglLkLuavP+CODS+
xP7jm5rgjT3t9xVQsUs8i0Tyi2xVF22/xJK/6v3FDybu+CBO8vLTLw3fUH+vnNV6KKjFIv895fHy
jB/2SBkf3WpwgeEfWN8FfQ2bYo3hND6oPRMm3SJxCd9P11VuoUONCOS8Bi506mFBcT3SLQbsHcHA
KDLWNn1Jsy2e+QsayTzjP4bfZaAYwMF6OAh7MuaVbpqBC69JVBO6exORGQHtKDVo+UqNVxwEbCRP
fpR+uufHzMw73VyR6+/2+HgDpVuHZ6cHr5/ErsN+oepGVXxGvmy6gfTGFHQs2HAAW0/76H9JwXLj
rdl2tint0k9X9jwiZvKcjguihA0pL2Jz3iqdTi4SuAMGTsxCRFxPC/U7RIkyoXh9HIobP4Xb618J
1IIoZtGlzD9kuTZ7rnlR7zBSHfqRjMh6vnY/kyS+Q47sw5A0mYNdAgnSaMficEQMvNEAacekOz3q
2RuIywZIo0VmchE+32Mqwfk8YZYvDuz33ibY4Wke7+H2Xj0r5MgKX6dsEAtkhMxIgThZJQ69OoIQ
e/CCneLsnnLcBCAjRWhMff16ckHpZYpT+DlpcVCKdmZMl18a+RAnP/HdM2ZL1lZQsW/s38bjPO6F
MKNaDFzcXK+AKh4CnrIgykTPYk8CyqQorsB7F78oF5x6uwLl60r88wsviJeU5NisqoyyuB/LwXD/
YHXh1/t9eozDpm7eiX9+q//H6pT95WSEsmSbeLokU2J8UeniRqnbiSfnN8qJgVVdacG0kLQk7l2y
Nirmsw+oVjeWhEL57p+l9iqwwYM4l4F21oMzYHAsWEvrU1oMYoefufL2HlI3p+qbhCkkt0qyjgaL
3a+sOFoFvWghWuknoRyG/9Bnj+wSGhIF5hT4JdhEYSfIJ2BAD1v5E2LY9SP8hYbF29k5d7ptiZW3
pE2Kq7IGV+e0ro9T/ORMRfkDzVpOztsjNQf3/QC4F/fe/3ZSN2HS1RWH7QeeBnG8UeqJ40On3Qft
sbJux4up7ZjUH6AJW1OB3ams/RooObqFBM3hCfkvZOKtuRoC4saT+VNpcJFs5RP92oJtRrIj9Go5
rZ1IflxcZKiyRItShDgILdrv13HOrxX3icpSqp+LQGcCoaXGQb+UlXZxpzndy0MTgSM6cX9Zocbo
tuXT80XgazyfCX1uTFavvesBlCbGmGCiwDwT3vAu5Gf7fKHNBy0p7qR2/qwamsXGRLy7PFfbVn4G
UxzDhZ4aucv1haw+gEnbeRrbXw1NPI1se4PGSdz8vBxLaIqyumdzXHAuy6AqNco9zQ6ujIA0GE6b
N4WYfoCUYiaGeaoumZdDqZcaGM/E+qhJ5A4CgJBg8jfj6kXQrpJhqpROvzhvYUQfuAlHjke5K6hs
0VrlaWKGlJyms/VNkHX54XHEjOAbDGTrHxlquGSOTKWZQhi4xIaxx3uNzcXKCNsoBVjsy6aYlmzw
cx+L+QZRIjfebSKme+Sx5o3u/xeBATO6uM6V6/MbJeO49hIYSdNrceWeQMkq5vb7z6ldQDW12v06
7MHffwFt8gRzLTyljw/sH+srMKbntgftBPjlqTUaVyVHCbKaUciayaniAW5rW1SWHctcz0qcrh5Z
+tOtEKIiUVKOB8NwPAGUoTcEzs+vrjzlhCPGJ1Sto9W+swgLwBfczTSyR4XZxQzGGOYtUlA61w/K
L7L5s5f23a76SS2fbOdjiDtKzts5xOd5LzdKjNTxqiRl4nBH3+c03wEoZ5iHFdW+OKZRmSxHEqqj
xMzFa9wCwiGbYX5yjsQtX1xvDGG1++2va+v2g29AGqPWx3J8tc7IgLiI1UZytv24uykC+XspuugP
LKBDjLOCR8JcoO8bdIp/zLEPm3W5CmDyFK3OSXLR0Xy8grYiblJteG40oMFxwfPt/eJTPVn3hlV2
SLcCuOSfzkhG6zElp9cjQ4QYb7UG5AVAsCrRVSfgi5E54lBcSeEmAcfhtjXH5eg0wBA3prPk60Z/
A4PKPr1dWX/HixdKWOO2U+xDlqZO9PDsD490PpjgcM/smhxlx8uvdRh/sEOF6g1cqgO1lvyoMwgE
LsHw8N7T/cRgZJg95G5kp2Te2q8P/MQqLo64YU2MelDVcyRxmKvp02qUz0h9Ash5wIT/BmpGSbCu
OYt/WQhtWbcoGxa03hEzlHEkWTSQGqDtLD6HnDnIb8A+bRzPDKVDOjCVw+IirS+iLpF4Z8dKt3sp
mkF34ML5pCuX56eoczKVbYSv+rn0aANkLAfSaD9WAZva2AJfyvmSmGzrU+/+tunjeBe4Rp3K4vmQ
Hhokiz9vcSboJhhE5krxlYbyTW9TBJSx4Aiwf29PIk1tzyJWdairxYoBkBdE9svtOgj/+5lftlo/
G4V5yNhSe2Q8GhVk+HdRjyhfkz9hL/y7QS6z03PziKt0FSy3F2G3gkG0wswCPYi1nKjd+UNOsvnH
HcNGLkNiiPpL7Qtld48xUjg8ZCIIG41dXhBbssWv7YczwYRxrjrsIYyLa9Ltl4JoS4dAmmnxSfCb
fuppkwfmje+4b2mSpVdYY0Am/dCWQlWFlbtxCfk3G/fEXpLHUNO2OiEePRI/l0fuxyv4ZdT5l0lF
TFZGcAjDCfWewWYkDUoyrlX41OV7k/ENwHBP5ohSWP1xTF/5UQryx0leytRwOmWuiRsgC+5ZMhYW
E2mDfbNpEaL3qkr7P/RW6QV2iNgQk4+/jOuLmpvj9FyGD3jYy+ICMeMmX7KaDslbv2IHSbwJoF14
KMNVm6ks50/R7W/dwxOwxH8C3cQax7mMcJS2FEW78cKXZkXRCa8PA1vgT7nqkGP6MgbbuHOSQIW4
Qt+v2wFKUfCL7XoM63wHOxww6nmdHGPgNqPgRi+7XNHho16ZBZxbMSlYU7s0c10ilS1Yr8YLgy1x
zXKnEW0YPwX63x/QwNs7Ars9sourJ4s1IdBkP3NGODSXFT8lSiT6pdpknbhi3G1+RFT1pZNAE6jc
qrGgk3wPADfFFEvLp9xAB66zEo63h2g/yvWVbK7IkBLQaV4j8Ty3pHIJREgiNx+/xcdBhnUibJ/3
0h104NZbkheSCc5DOxpuQisb3Tw58+VYQ6giB8M8BGiqAOiKVZHkxgvcI84ocA+OxT8BfejimwhA
S79198H6ilD12Ea5Kb2ENcPk1REMkmFnRzk4Sty4psWkUvjYPdlxpxqVS29b5OFTIwS2tgNLPRpx
BR+MbTg/AO/HqnVt9sGID0laJotk6kOzN1YVADEGxlwZDcxB5Qq96UbBCFbtsTDblGWu7LDzdgaX
jV/g62Ut1E8WbtAyssKpXwc1moW9nv3TvdXQ/2cqYzD808LfX3k0ipI1wvDIIWg3SkDnsPEzbuXK
eS5ym0rgZGxhSmc9TrqeEI7dOKAd622ncBMNQ57MukUa2lDW3SPtAlZF8AHuqESQUZTbtGESR6Ak
2SL9YdmwmEWHY3GtRJFYPYe1st4MH8pVxZQ8emMAIktKsekJ1Tcf0C0oxMJgnSJHvpYqlgOPNdFL
rLopQW8US/oiH1/EWbTWucjPnhbZ6eqwBLKQGKQCQVgJxqOnwVR2ilgxnPEk4e1LDAPVVxQ15r+p
mlJkuydrG7ytNIWGYsWhCRJxnUNjw7ayELcsUlxGzt4WDIWnj3PzazsOzufgzqS6D/Gn6NPBJn3M
lRH+anElUP2Me2bivzJZFX/mWr/ao45IH0a2chD5mPe+nGRnluyaF6V5kaNOxhtfJVH+XA3ulcoW
ewNGzh031NS8bOanCeqnF66ap51U+AapH3z+Sy1MT7ZJN0Mw42WdeIePNoqFjDD8Qmq8nVQTQtaz
7WbvXAKEIOKyBVW90Z7ZFOayo7jPpJoRfp3DYNshCP14KeSU1NV6imm0Xil5zQhpUapIkw8Ky57K
HhaaYuQDFZl5bdQDVt9yGk12tLa69UBe3agVBVHFl2gmizIY6ofO1Lyr0GpS3gJVL9hLVovBEF0C
RnGQ7hv/ZX2ISD+hUSHqkfszPTboOwDC3FhMuiv0DKj//3ltAxPQt7zrq37PXSI3Ws8uaamXDywB
3oFzzhllGZpoGGQz3maWJrD9YhKyQlq0zHq6/RdTN4lDQ0XdP4ZSC0c5Ls8ZPjhkXXQft1NdazjN
JJOglGDAUKiptrAE/DQGrDISMfJ6r2CtzJ3VpvaiWKC8X54xACosVtcLw6JGMOBX/91M3YXP8ZPi
XMG5Z6v47OI55GoVag2ZlqezCwlFo+ZWCXEMXjV/WIe1QSzXeQoyTTMhi6DoKEVk0wYVFNgmzhka
u4jopn3ZgjmdRJEHVcvLplxJlc4QN5Z9fzoFzFncIMAKHUV0yPK9zDirKyg+0ULRtlR5f0yJHUDF
SJ2HX5chgbhsbWZlIjN3y/boZgwsLSs0BnisIEcWj6g9aICj7M7KtomYJpjxc2b6+y8vZBumg18/
iA57jRPnfVkeM/PeFhNu9QisHYSq7yWauFTRCoaC+VgDunEaHmx1Fz9dLSnmzCnSVEDA9bUsCo3q
VhME2ViVbi6msT3MS3ypRF/Z3RIHyerOrxSUb8IsJAHyfPYw6lPaPhcpCRS81U6aoXF77WW1rM0W
1BwfHjGRP5leU2p7scK1tqDNXRWAAA9HabI8W/nCL93TrODyDky6m9DMEzsB8pTrVeJMxrtt9XM6
I/qHBcfHU1pkGIS3jo8lCcMB2YTWaJUPIdwOnDNHl2fvEutubwnv8dIsebXKrDueukCkUCDEeFWl
RS+ZmlujtvkqwrgQY+jbamFRhrqSLK2CPhZX1Nj6colMNbLpgqc0ZeME0KdycNGSUzT32Y/JcR7g
C+XDAlOcB+HGIZxurG0zvUklqVOKSRqikYvPs2Nc8/0CoRD7tJANFK6TiTAqTsFXdqEASP1Ywqlj
PCO4PTjCuIb4+WKcBWaMDpCIzdCKO1+W5YSBda1FsOBC5MBM+H5QZtdOVYeFQuO7D9pWqNkgnITr
1Y4BmFheVpE6byAeU+H4lxUDMZQ8tG9rZCaX+SPVD1hvamskOtNZ6kFlo6auQJdL8xNUxX75KtuM
gmzHs6oC2KhjTOOsBnmDMcqnpJ2nNCTmgB7w6XKFnMGaiwiRdSi53vufSiZsYxx0e119p+wwal5U
RmH6j39QYrubbCuLuy0W50DzbUeZZ+29cNRQ0+HN9E9gP2hcsZxFvO29jV2WkHxvKBw2oU2F/n5i
NrtzNqGRVhE8bEMTgWAmHJXWs9MpDb+3Dqqdgk973s3jATES3uwb0v9hsrHtghu+NAyRlAD+Ic+N
gdQm8fXgACJecO4O7akDBjDIC1T1T5gJNAXGOiWda15XSmWZFuQay2+AhObXzbgPRnIV9jHgp4qp
YM4YFP5Jpff2DIqZ4uNXFspvfTqUF+xfgG1hFU6Qftb7kldcDnJlu8Rg4tTO3/dyTKkrgBwV5n9l
ABlPptM0FkWa+lbr0onZOK+h0r+fT6JfMGF1NfYNHmK/KNZD31tKelm9ioaqO5BbyZ6IJoj7KUfa
wd3UjhLOmblpn5HFcA7mgNgfZDORKsVMn1DMV2ulGN0HDyXrse5WRQGnYHJIbF0zn45xMBIA8PAx
Lp1xHv7TArUGMj8XaOir1q+1njNG9M8cd4Agf/fHpmzBRz4dtudKNs9DiAENz7up0evTJ1ky0Ekz
UeFSlHW+WsNmSngbcfl2b7jgfB+mzZoEeXf/EjXliu23gtlMdLCuxN+Px2oSsWgkIF/KqWaZ5pa1
uvKs7J6E4Lga7UV1W6y456X4bxygn1toEkjBLo2MwlgVdJgpgP2DZZJs74ftBOofxUad6OH16sqg
l1wzKqIZwutZDstVdLZZ39lugMkGc5VjVUBklagesZLcBGwVKAW6IOiBv4ahqytfs1ms6yXEBa2E
5M+ZzgGheWBoN4wct3fUl731+/p6AhTo08A3cAG70NogTHqIxwh77D1+TAOaa6rV1yqNjHhmiz/U
adMAukAmcmjaaM4OGEQ6rFVY/mzuAvZkceILlS6c8DcuskGuPgGe2DWX0BjoziMW3tEQ6ASZHj8R
o5kGuoTBYOrz3GOatjJHTcE5sAJO0K4HDJeAk234raY3Qn4cMjcvwDMUJO38mxoUsuSnsW7F8tFj
onqTEIdFDgTeUJ13DcaeX8TGOmLpxSmTvcWzDVHsqGLOeIgZTBJ1c2Q3WFJ/hNYuaZrWWIxa9KFV
LV2EsKOou4zdtqpScaiKplP2qY15qB7f7HDTdwZwt2To14M8LqK9BPyYAfL4+cgv7iNuPdLGZyqj
0TWmGFd2kxl4pfFU20Er766QbEloDuUl3SHSS6Vv/+sUIc/ExzPvV089Op6QF+bviSib4kU6m3sG
S2aSndJGipFrIVPA8LiTeS4+nrZ8F6eFM1URQTjX88PpYqbNFnixxMUMYLUJ87u/vAWarLho+Ya7
KqCfHCR1TOZXitx2d9JGXM0AiBDJ6MEZAzOYiNqjmTEXE2Z02jACFscJjkZpLLeIrra/tN8fa0db
6HECnLGSM0FyFSMOFNjbJ7tg3y26KBqWJT935Wdf6ilBVhq0iKmovU4vCIsQpNwDd/eyVhQcoWS2
XFSv0veg2sq5CxopZ1M+cPJM8pqD63sN7Rudq8tX8CWMpylvAVacW0U3Gap5yR44wzDUSMPDMeav
/Tm2wvp4JJSz0KkamFgdb1hvIrtW3yrtZBmD9zwjwN3inktSnq45urdRQg+RyrCJAABPDQh9kVT2
TwDC0FI4wQY7uUowVtyw4NA1TvYZ5j85Yd0eNVJ9pTGAbjEcMIWDgk8rVZ5no0tWgIzfI5VyH4CF
gv7U0C8j0rulatkRAgdd1KPJD8JwZi7NqHrd61RVwOsdkbxsdjz0tSDh9WHiXW9xw//5L4qhbEi3
YkIv5DZLKMy50zPgSjlOzyYZL3CeG4dbn/jEfPRJcbeLSNre9ktL97RDGw6tec9aiR+Jio++hzwe
DcCe5CvuS/700FKpdhqwKAzeb4Dfdg4/Lht2l6agZkhtudC/VSWudCcoYt5weOlDH1tpTZ4Ly3gi
wtGNHOMlBv9KQ6ozw4ZkVSmFF9bMPQPHwTZD/ePpV2YtB2Jnac0GFRmAsyaXvHtOzZ9JMG8cpfnm
2vOCAplT35zU5vd63u+02/+8HMXcVz7L7yi6sBHpEl2mxb4TLdMxVIHcJbZZCdxAv2SbI67M2LH4
EscnPP74UK5CnbfYKuiYnrFlSzx5c0tlP9kke/gw1d8xaCvdalkj64dpkH6xmGCctSiZR5RFWtc6
+NjuWSTxuqetdhe9nDEh7R3s0gdX53CK6ezXCt5Gzz5ZyLE485f+G6EfEmN4FUBSs8pkFUF3rKdE
D8YGKKxzwcjIV+MT60auv6qmfrkihPpPiUWA2+csgKBBYoEA0mmk9j+vgOEY71JkBy0qKLz6jpSQ
KUBnpdmadjb8WDqBYxS+KJ9dKJ6Jd9HeMpQ56dvKsB4qz3UG6kgS25rmejQtvdVCC52tq6SALnI+
TouUVCKyy/EVymkAB5eg2HgH84IrbGSurHpoVx0w6SZy5sythzxT/lpa6UEXrv4OhmpMEs79s7Gw
NXYTn43ryyEhxumJmRtLA6FA/96obp6NSt4/ljP8Lcs7vi0vDmJArOxtJ7/eezIhIQTzDchUY+to
WIikNo4/rHqFjvX1IdbfQM/r9d6ejzAR27z5MCm543iwu1dZ+TcvCdBjGm7WF7FvzZK3J0+VW/rV
zUEGuR2cCKhUctiRJ3H0UcW2adNi3ptLkUeTBnqB1KBgT8dUEIKMGyAhzkYk9IJ+9bfjB1Q38bcM
DxjQN3J185duU3zs9eFKOxwpaUJ4t328nN1FQDxUfxjnzbnNCL3duxHlV1Z6oRflyN78re6BJNUL
pFBRlU0h9fJnUhXEYm4M3ZvJblkH5PQndRGMltGbjgJIjHpsoFU8mnDFIEZgG3Uk0OGpfR+gJsIT
4tP4sMWJbshhUxXnxglfIC/+VyQEPM5H2mt1z4dSgUBxV5oM4W33cs5wcE6Z1fnqFedLiA5NLZMq
KkVdvGFxLCxyZNh5gfSxvFKAw0ecqfS983OGGfhjmoXJ9IV858J0vqEAptz6znPVQ8XPyQzKEfBL
WZCrKO2AYwMhXXUPKLRpNghSOClCjW0U2NxrtYKhgYEr23CyKniJ7Qt2/Q3189ZMyyG7e50mgZuS
yu3wS+J2wGqyX+6E3TcIJ44fMjIsXAVN/51OneMnSXF0JWbuCzBvlEvRw82X4K5GfxdC4A7D7fTL
0iB2187beeTLgWL1jopvQ94ZeaPPa6qf0zfxuHmVPPZmVBmR4/ONnXJ1v6aqx/9SKLFF080ARczk
rJt0Aq50b7g2hBGsDbZL73oLH1rwP+VgoHk3cEgbCj7RwUcMfJ50vYgIWYskoCWKNZsL3f1jyxgR
hD53Y5jAzRMFuT4qdZbWKWTAYmNHHyFE4HGvSDZLJ97eGELKNaJnk8z9n7uXvm+xKCspRKUNkcGz
kK1n6Hr9ncwa4QEpupRkA3hvJCKbbQBZT2W9mtaoOtYX+Kz6h20a0THv6PZsEq9yqgK72VwJ/KcO
4alKY23HJVI6mMNZNtD0BwKaAhUqy571cApDJ/joLEPFewF9uWT9CvorNA2rMLt3kD6Lx5Idc2Kl
Qrzyaa6KDLpGKmHFRRg/BD0Ev77s29Vru3+K7DfOxqB8YJ/pxYWOuLgRkWvdnHQpSMMwvEb7acd6
o1jIz8ksIwG/btjXmb70mN0wRfR+m4GO0sdhRPMF5R0c8ChyFbiPVeXOijSDP+fFBfQ80Ia8S4Qz
TzxHfEQKjXbH2MjWya1b78YFjwMTJa07D6sct71Nk5n/N2EZ0iyF74AOxYJJjMyDDnUjd8WcgLVY
a3ZZ/805FTZAHEdLq9JYrJAbXdS5WirkQjZ6klui36iZ6iiJLhutY/FX6jUXohmCTuBe/ePF+xd8
c3u7OQO1stDsVlq6P4GvNXMUARLzGSQMzkgLCX4YAhnE50u4hAl6TFynQSGUjoCQC50/znWFy/xh
n6d3PdTQ7aDtWZG4YnE0I350O0MZN9WsoQW6zrmCLPOcI9dwhc7GFYhOmLiNOBwD7zhc2jUnmsUr
s2UNG8W2boi2LMe81At8aF16S6XKdaBwuZXxjjdul9fz1aQMaQ7ZfVt2aekyVaKFT9IzdpKvNsWG
4Iw/VxzpuXoKebAgGVDxy7XokB9HpZH7GQyVwNq08MIQnk46kjiw75SjH1vnnIlJixGkgs6n6w32
nmiec1rr89IidHB/J0twXNjPYp4kFJdja3QTPNf1FIfeHhmpUjymGDJlcuGbdeLoPUMDdKv5h8DC
FfV/csokBN4okPek3uKhLqAK+CmGHUJcUEw3BBzkm0NER1c/DVuNSNyObLeMkIcyTRO1DtVOC5xU
yyw7d+7W4nAkhZl1bgj0zCWVIg+cAOQsI3oF18V/U+coT0NueQeIcK1PmkYEhYrdkiwO41yGLMce
vp7VuxIdrHtRhVwiyQDLxkH8Pv9DrA7fq6i8aXHo9+n8A1J5OxrHkDu1vvMxKPswb5bzD8nzu94y
Dios+dM6dWuDBqejB8VvvwwRTmi0nc85909Fv0h0S/iRMkN805cBk3YVwgK/yWQ7v06mGB3KMn6N
+hK0r10eFOuN4S1MmyynESiii4mIjnH5D0hNy0Y0pOQJFKwdFLELKdxRC7y+rfny4gzZcv6ncJho
Lm3JecrPbz3Ttq8m3nntxaZvDfepKpgigvxixZ0RVJquglfHVENwsOKL9pg1f9cMRKbd3Mbm5nT4
3+IVEy3h4/8LYiXwspE2CnwvgwloqXV0iXU0arymWpZJsf0wgxagQ2OOsJdgj9/sfKa6HeBgcolW
Fll00aKDP4APUNTr+OAkroUf3x6SXwMzyW2QFIzGXGBqa43fPvqsmMr9Hx7Gz5TY4wGmaEd/puoD
FlqttxmFwg29YiodxNn4tu+zEGF2Cna+PGYLrj6cHv1YLOpjPDj8ZWu33hTTGo/fzWyj3CTxxwJB
DO7fwXvVOkS4K1IlLeM5Zdr8GAcKGGp5Ibb6haAj5s+fL49TgvH8wM2ZeXMB2nuHFG1ZPIBt9uvc
IxeO5n66xTQZStfYOQG5N3A+xOYLRQyyBjcOMcUizAkgyaAj65GUI7SAa4Fukq0YuqaQB4KmgT9s
f5/XR1dcUMhJEnvyxmH7pPq3zfH312r8MO75qRfZn0cHCK5F/7/RHEUmHXZYGsCZ92hUH9QbR8Xz
esc6aywCCfrnZ7+h6ERiY0qSrvlLS2rj4XEU110uvthy7Bg4KTJ31LoCGZFh5rNe+BXiiMHPkfX3
pHc1JFdM3w42SBz+zYFL9zLKaxstgmnc8We0FE0wLoZ/v3HAWez3CUVlHwjTpnQ+9XM/+zoOHNGQ
3G54LJ1gi392EBbFFDNmluVeAq7O3AEfg7VngRuvv+s4wKjoWksiKJda6448X39KggJ4gPH7aKGX
PtDR41EIrP3OFsd1sdnebkEcLWJ5qymYwSAB6ESKBVRR8tjUJ8igDHFsmhDqz3PTtSq1XCMRUc9Z
j2oaDp/4bLl9/mMnrMn7qibkBuvGmafxSnnBtRxvH8LMNnqhE0uPozL6EbFlH0ZRPB4WDc1Fd+9L
WIwzX/Eo5c6rmd2lTYWWXkILcaRJkBN7r2zIgSKnZq66EirPBOs8gGHW1cL4hgohvW9vMM0SVyKL
Nj+xeCu7tBjFVLFyX/xt6jBFbfhFhj4btFdiBRAjaGKgbGE9MsT2hrXBKbDrc2VCyvwAflBJhJhj
MIPaVyO+jdsWW7S8crgUx/ptNPvHu0W7uWM4L14eipQkklsLqNU2P34gYOy4kRswya8Oiv1hhpYn
XqwxCrsB1QI+DSt4goUzxlB3aCbuPwH9/D03g5134mvPa9vKIZwdupfzVFhzlqcP28tcPX/WTD9b
ml/kms679FYThu5pwAWxxZxuhRWW+8GhKTXWzr8N2KdxEtrY/4GGGT+kyOfI4Au1MPiJmZyj44js
XqHc0ccDyXfQgPp4pln+5ji2xZ0BDXcfv7Km8x0xDprrmgke+09Walfzc5MP7/K+oqkCLBgiwq7Z
Ak/3/X62hzpDx9bNkgoVfuinmCUNvEC+slI5eeBuvxTkxlBxY5qUySu6C+lTf68+xudO/GNXD0dD
HNGqzQLgAcd38VM5yQ1MJ4yx2zYT4NJEo3AwrV/HiA3KRsJCuRvSWxUkya4OOQU6/qW9/+58IAxT
/J1kuGmrKfSgM7lWbB6d++oAsr14FgPTt7X+y5mOe9McM5dd8sBJp3+kdnCJSIHsJTVl/HPm+NIg
8zii4Ogz9fH906f/hR/Gza7LNQDlTTRzazW4DGx6jokTnBQnUIOTRRgG7qAGLyNfE6/JJv4qv4iO
R016TsVVm1vuj2id4Ur98HYM67rZyaG9ylsmm1HSXsPx4hXtCVjucUPpaZs4cWRjrLihjMq+sF0o
CzJrkASnEJFVk02eulPowCErGE3ShqhDcyGuYCMJq9iQUnAbmzaF2I7KwYNgUA8AETik+wqJEfM2
I8GCdSlNyu77LUMRR/6NdKwqZ5PR/4KSzUGX4XNtFlEWqhusEPXxZQtJPJ8FTAtQnQgy4FIcgaMf
yrRAx/03aRSG7cMs0ayDqRaDbFf2r1fDDDWLag0lYJlgt+X3kQ2/K3hgD3BTfH1kZc/la1qCUoRK
eivwTBL9I8bPzP+bFL8PdaxVflFwYNrjMuT3wK6LiLrJYPaxMRkLRnkpoxB1qyM7Pi/RGYcEgpRa
AjZcZJwgs38FSvXuV4p0g5H2ELp4TBkr/dl25iqKhcHoeUjSRXMyJa08v2mUYzDY5+Z7wcnZ7SW/
S8xxGHrSRqkLj6lA5Hl+tA9Sm55rVHJWuoF0k/iN7HDoqcApMZ1NoMvuRVelJejY9FiNuQ9eyerH
cR8pP23upkZoy1MAggxj4LS3oE17z8a0UoolYoAN8anLShsDxhjBtMsGyfluno612bwCoTZyRLj8
LWBByGkXvE4ujDxkaXlk2X26ZTy7zZaj1kwlQUyVyBw+gL/nDfu+pWiAcJ+ZKhbSMB7YTvpinMgl
GyC4injmaMn4LUQa8AhYRL4VRYllvR5HsQwH6YNAdwp0hluN1GnxlQyUZZWYFXdBTDm2ei256qkX
/zKDcf70mRghPGMAbKg/r5hnr0vQ+2TW/D80htcus+w7ChMPgMUucncT0pa0fmtzpDWWx+zkmjLY
wcB26cRJ2CAAjsYCr3ZtMNLbsA2UCagld0VXxMVhy/+th4+nWtoLT5WxT2rcg5BO/xRhtqyrtMMB
P5yzJRngoSAjr4HBOBJZW2YqgiprCPskAop3KNf21nCvdO7TA8Exg1q2txHC6/5r2BN3ePXjEVmh
ZtRtcIkZEpO4fOmjnCXSGTAfCad/VXvAn1n1FzkgVlHyIfiSPUf1KIDEHIi9kpkW2Cxw5s+27f1d
ryp4qoye0+Q9OdKg8vQO+pn+HyQiVpUxkUuhQJYKDP+DotYnngc+iiWt4rTBb7Imqbgjw+V02PBm
Fw/bhDFBtR3b/zaQjz8W943XcPo1qopclelN73sbpTtL4gRuV6ufoE4/aUTBtyuKBLzVlKnoX/6F
P5G5hR9h0MhP8OxTEY/SjdkOPQKf4iwmRmxFsK1vgkioBMKw9k3V9X8FyVZjiv22DZZnZrqCxkVD
IIJIrVh5sMj6cyVYJ+ubtSbaYRLQHgeT4/Gwq2JdwsoofJmFyUWul0y7IRuy7DWh/AY4HbHOptEB
1xGYW+RvTBTot9bylIPkU3NOVelgswZAMJinM5BBHaSVPoQGp/xdUZI/qPda1XJNZBn9Jz+GmkWK
V8EvZsX85W36XO+GRnDRsyDq1fT82DG9WR8pWNU4ZiMxfdNTtMpRP/2h/p0XoB//yXD6qxx9BJKx
vtdfY22g2LjnO7/Pv7IVEefq5+x4j3eCRIe7NqdWOpx6Id3lmmrF8BFCf/QYuhyxtGGN+BCgUpGn
H0upqf1qwgqU510ZZh3dTqZpu5/O4aJ5H4Xb2eFOQ66ZzAERd+JlEuX5iGtyUK+YsIagYPlTN+/N
WsWrbHCJgsyARLm4bdHbCaBu85SqmmtcrfWy8a9sJMmUkBb3s9w1IDCJalmiXMYVz9DaGBhaYGQj
dD1iGZ6eX2AGaMTOfTWvDj2jok/MdFcMjihRNaTBlrhSMSrLbD0bGdcaRc41K1R8cFFJmm0mLhkM
QAPoX5NnjkdsOl6HxhJEDSsq7E3khEXeyHPDfg1qwnI1weiE0V0iuDx8Li8o3qFIPFuGsBe/qpw1
KVTzUcBDninsfr6Amt2QwY3nCX1Fxpd+EFG4rAMrWMd0OB9K8VTO764MwKBmMnMpQeNWoTQZ0ejv
+D/JVvtH8ikv5taRp9ugiqt5UOODCoIV4GZ+VHQPt4vq5lq0zm+o9okedMhE4Vg3Wk+2GhHNRbfz
dlx4av/BhiG9Nvc6fF+hH9XDzjEjyetWgn4geQ4fzzYP4OU6SFqIO9OIi6Rnt2qFRmbjYfE397so
MmwjtNi3PuVTHV3vu/ecd6WoJYRLwj6KR8qhgpzSEy4azI3nlDxhOtLV9bM2nrvt+nIEfZH4yNgc
zRb2MMpiityYjNmvFUaDQPdgLDfFIbXtlST4avoSgL3I2HocU3n2n5r5Ddwv2Z9bc232ntYwYCbg
AnL4r/kZlwoooWi42DLjbPW14x071J0DisQm4SLVX0jvIdwsaQ4lOyKkVDajj7GnHr1N3088N9hD
BVDfsDFZH8IJH53TqlHPQ314UoqNW0wcvA8Ab028p1zOnhD9V1gAmxd0iYWPQXzUIhY31DzpW2rP
zEuuTFjpS2HEz93FZ4IiLH9q/MCewm/l1DSCPMS8pGzC6RXVQLltPN3ZINUCk8GEK8f6IEXEGASQ
/uDj3CrKAJvKg/IktaCUZPdmQVKUPGs5mUw6uGZ5XKJOqA7Z/kM1vH1MHlYPfGXa2gl0m9WsLbXU
KB3NC2KByjlGuhBq4L/BwOFVoAYzImBvzReKp92uzhGbYGHs+o4hmnrOOiQdDIrTI8IP1u1J//90
P6EEjL2z5niMDBmONzPc+EepfATCM8Gpe8BKH4iSfhSMYoYJsRfLN+uKKy9OxbK1n+cMMI9nPmPT
yaKor5eh+QGlONUC9npG6hMLLUPZYMNIWu5NyznjYtjk5EDo9vL4IgKZKLdGqsXZNV6JJ7DS7pCv
CEeFznj0pttKZMNp3RTrnMEkVdask0DYHw8cFnDzC8WN/fwXK/th7NmOKctwbSP6180MI5WKwzgi
BbzMLL/jyU4466YbfbOczdY2wbJ7V1ueWaLYix3zCICFLPKO0z/0mOpRyxyh1huenxqOQ+DXNV9c
xK/+YkpxkefCsFEt+zxHwUqZhVFfZWB1nvGX6zrrTY+ozGbqMesKrtKK3UUqrGxWuRuMjV++82rZ
nnhtbesDvYP65gc090NThBBmi2iLeU4AvIrIoqK7z2puIvY3nIJ7b2q7+P43LV98a8DFtwyOmmB8
wRMm3VSZtnnrJrf44gXl6cbPfAscOe/Puy+zPb44IGbgGc+dAKFXkLryFoZSXsCHxLyFV8tM9zmA
ZIRTUyxNFD9q8L2p8XCqt3M/leP3AnhXdJ3gP9BPy8Uzolbj0W4jcsk+vb8/RAp7Qk0wwrG253Cb
vdSotIcbxEER2mn22El8aEkHHG+nHa5eh5gFJa809+LkfOy5Z3ECFiBlJw/TKr8fVc7JtpYOJQfX
4aIDiPmY7JZTHT3K23kCDtWqe7UkT4whwSAi3wCu1Y+Xfc6G4fGbWExoiM+bc4Xk4FCBdl8LD15L
DJf7CCOp7c/2W4/DDwA0jkdWKiztS5V/4czlhmdlcT2Bpj1YBode47cQzgBH/NhaGBiCrdynvnxN
XkR1iAhzUiEOyMOKmb2Ue4pP8biaBAOEJ4YQXR2EdOALK9anTU9LTTMRNEtM91W/qRD+WAC9Gyo0
p4IdMf/bG5AtPv/jdk8erKg/RWrf0+daLhrZXdqi2jrwlEM/1GR3JR3H3EH+E6KC7LoQDFSq8OE4
/vMK+OuWDD6nFRHhnYy0TgESs6hefGyFo7MMUn7/GHtgFc9dDMfSuyyGbc1GK0+X/C3DhrxtSvx1
wLWM1dzjq6W1Zw7hqtRG4UGIZonIs4K8rij4Cxg1/EBXRlvs6tbtOSuOLWwJAZem7b5BC2cW4++a
+1cyIpC4SDBhk2I0Hk52o5mVFMzzEbViMOrUo1xr3kFvwlgIy8dSRIZa/GC0yY+F38UDpcAQ3sVF
2aUsHKHe1W0zbSXSk1uyZeu/GgL8LRT7NL7cH2ngJa6SdFhHMD9Nv+ZVUK+YT5N+WhfNWsRIvstp
4gNJx0jyaX9O2SnROg2YNNNcHEyyKcKZwzatvvgeO6Y2+qCUMFFoSy/k1LODFKngTy3Wi7HR35Mm
QyC7O+sVAmOMTK0yAiXTbJf7pibl3rWAl7IStXZtdd2Xo5DkQFGZiBJxJ7IZi03xUopZ+VZfUkkN
14wNlaLs+8vlKhT2P8O4Mwo04RvZzavRmNMaKa1/fPQiB8+mq0pqdg4eg8u2ZFqRXPVYl3CRuRXc
PJ3nObKVJYPV6GbxqTZtoARDDRIWAg36e6muGr14r060+JGqeiMu8JOgoWGrYpX8Rs+/ch5LjhoX
PN+MClelVt2Sk3EDnhbeSsebga4I9+Lbea7/Xvk2LSOtYUX5GmiZdDycfRj3KVLdA+3ICDQL8rHf
A3SmQSsJc7RTbQBwURpxLbUcc2jAhU6LQ+UMG31e63nS6hlKy/Xiygpk6ha4ei2VUIwZ4mzG+ykl
soqS0HETEi6rMyDUVXHUdCd6DEn1hAlZW+OI0fU9pPitXZhVW894gqyk0AoFpusQ5rqRl95uUUXf
zfiE+v0SBYArmB37B2jozYkJsXUmQW+/gKKNaiCvdkiidTRUINdLbvghDVeLmn5R4/to43dz/gLa
MKGATOmpb+YJvDLmWBL9gdcyKpnqB0vx6yQiVzswyjdmNGW+hiBOY3pxcMqtTomwINr1e6zZOg7V
Y/jKbVsyyHrcY0EXL+ANQ8M6MijDui0JyhOFLEewlV8cbEPgjBPJubCT7DQ7VI8FxfVUlEG2fbuD
g5UaC0pnRTc0DDKKGckJ1mDTb5eXj6KANaRrM7B7GCNejXNsViBPocfh44q/j3VZQWnyFaHp+EQi
6plwU2Hp9T88HLK0wLQlmXLn3e04Wf7N3IRxdA5YdIgTjLhWLRNCwf/FYicVLCVAAHbcxqhMxvK8
mNhxyFNmoKdZUQ2uuJ/RTzuxzaB9lBIzg5/bqgYt7oVpML0rtGq2jlf5YWYlEuj6dL1Ef6mV6j+L
Aqrxi467vnaFSfcBXvIHKVNwptS5OLzFbTARlJdU/e7CXWbRid9Hh7sHp7b/RSkIH/Oa5Z8Hvx5V
0P2PK81LyCa150guedjs3uKtLQYp1TTYZon5/LVW/5PjnFEvC3VG0Wl7OeWPD7RB8qWEB99FxKmh
A9DTTDbs23Veva2e/9x1ctfrolMp3H2DOGW9CAltGhbrOKorkB0GnLSO7YRvpQzB8np3SjzHUwIw
H02glrlM59LbeqspRipRBLIRfY01D27+SPDGVpHAJEESbciDniGTFbR0knUITU8+V1sWYu22VmJ5
k5rmgOS6X4txa/rvpmiCaS4SGCe5a8VmXV3a8oxhhizYIlArAoJqFhbm5s05fpKHYOi2HsAlRBBl
XRlRBLopZEbczG8rDFWluJQ37mnO+Ju2/VVHnDKNA2VdZmMLPPdzctLx3voSxQmQ0JOhkPrahwUk
V98GtkU7L1jC/DKilo8ubSRJbQVw2nHX3cgEd8isNKTxozj/wQjN9MwzwKok6h/la5M9viIg+ghu
aVLYW/n8MUBcSW6fWql+I09fGks6nC2pKf302iKB1KLPnySOgw0QW+J66YeCZCRJc40Ude5bJ9G1
wSjSo6aQiHLvwlX2+a0ZjEE/FQxSbX0EWDMIeIaQjz7/VRgZEyymZFqBOlYeFvJNMKs1Cp2KHmjk
pdBGuwtsSGfaDSeZvshidfQQRDTjMnrxG3yLQHyQnf1JvzVqAl1mlS3HlDNudRpfeNy+Rl69D4VD
bqVzXHROYdN56uWppyQ+yDkO3SBa3jCoz0f0erFQhDJDs8+BcJcErNNlhqKrU2gdw65C331Ppd7S
cBeSUhCV/LpFR4t2cX8QP1s95MIBqyaM8ZeHqqn1fxDZKmBVaObW+KH4raLwS1NZiHfDUu8Af74N
5DuZ/fhQ+NJ9x1gz5vQNXHtGR82nL/mSiSzZopzd9fnO2HADMZ2Tjia+n6DKkagSvzByb0R48LOw
8K7bd3IdLSI+oQGBm/oeiPJiJToxs2GqI00Fci5KulpjTzbMYM/zGb03Nz1A4w8oeDDJmqJg59Dz
3wazRC/SXvJw0ox7f0z4p7E3v3qZ4I+GauFdIWN3xhq3nekWOm0Pje1SQLVfORFZb3tq2M0Rhsw2
5XSNFbssXNnrbFf7tdANH1mSakAtg7ER8+Pu0mEzrKM+qlHCIujt9DutlyS8ieOuEyTSP5NyUixV
c0jev/vSjqWPNJvw/JEPVJ4Xdde2t/spczAiibPb9jD3cqifDf88egQeoDZZOlTHkyy571omdHbV
RDeCnDA90fcOw8LD9KDSaCgTtG8kv3MsPVCEV6N2+HVzpk1wINdXlpwRs9UxSLw0aDW16MTnnrdA
G3F29ldKyRFSZrzx8JwM5W9eR/YVvPHpGE82Go54b52PMz7HiqshSkvcNj2lvxe97+RY5RjvXzNM
WmfO/wJM9MhEwiPEIKuU8Ojm0j9iQek66jxqUj6GApCVxSSRbso6UVTXf983z+4MSplZfoFTi//7
re71Waus1H7rT28Gq/ir4LrrKwFRABDI4dIH+xbHlV9CPw4Gw+ZavUFJdowtPbVB0PIuWkqpfHIH
wnX/retrvTs9nw2LYkERVD1jm79pKi/Fy0IsPCy2sol0Nkh8xRYGeyG83raauPpbe6RRuiPimTPx
H3bFBDQ5aUJBv8RJ/o+UfhMpZ/gubOZW0VgPMZAnAGtiwR6dtSNvhxXTsaLVO8w0TceC/8HohiMZ
TBTVoDA5lCrNR1VuzXXMYjo5gIemOzWDY5QnCen/Q/7fFY4KwnA27mEq90ZzBEiCXqhT8o+oVy1j
yjvkgK36jy39L6L10dcNVscIbPkDaPSCPT95pla3PzwVJ8+AdEiwQKdp9+iy6jUDouH4VAsFtzCw
51MuHWDxz2Z+8hL7r6lJ6Pc5FCqjRg8Qw5uHfKTvZGaBKs//5xyKJO2V2oQ39HdKoKZZr7gMMiAN
3K2xVMhbdRpKqwztRNt1qBfmAzTA7QiBlX0BeXiXowDRnxsfUr7szKjCiV+3OpsBhH7nKpTdKcCt
ZNBYfP9bJcOy6EyIvv1QrLGicVHjiqYf80m3BEfiDCRH+dXMjsijcwJnhZVMF1d9iLHzjBt3WOAa
nPTli740V02GVFy1k48e3yyTf8mrwcV63ldLdtID1qSFFzxgwsZe6FU/l+AI1olb0KQy1ikcg/Iw
y/i9hOlZTHGhtcEDDfB/mzMz3eEGsOYeYpqZa5H7lGkmyc7JNzwMqmH7+7JREpqBnstX0FR1Yb03
3DZajIuQHhVvsB2AFnmlebRz4pDqUcLC2yGd445bZxiF4ffOrdxveqwnMaic+5gXY5i0i2nOPpwp
/N13Hw0YiQJR80R95M5m2wSmBaK4gZNLRR3xt76jg+N7HBCD0NmQidUlEWjdPE1CRhLPgEU0KSME
oegn2pesmj9zFrn4e8lQmyXitjymB0GtgTzbH25ULLXmEvJ6OZC8xoy1ZqAGAI2XgKOrZDQVaVfs
+VFCcA/q58sMxta+xdL1RiLXpCMZ22uIMUozy5+JgoExe2HZUbL4pl1EUU9sPZJ0206fDv24MMUz
ma/UqKS4pN8vXthylUKhLDAOlmSNiwstMDAdY5rxdorQPFe5KJhrskfzPZlO4YzTu3zrm3niqH5j
YsncnGlalJzdzDy5PcKk6gbF+jxpXerqq7Qxvi1stdQl+ao1gonzi8dNhNeUMmoDXRRI4ND3pcJN
BH77/8FmAE+l1j1fchFcSSFGpnI+jUG/2HnJE1nofWwNBg30Ov8NtYrcBpj9DIRy3TqummDdiDiu
Od47gQABLdo06IBUvOC4Oohl1kTeV6+ZqsBa6Bu/lEGIia9SoN9ucMxkA3dzfKUVtK4/ARPf4ipf
Gc6mSSC/8IKHS0OnlDCyP4k9R9642QoaWVBQgYzK4r9+JToAYoAekCmph29IQUDHjUnlWztC/tp0
vtwxX3SJAm8h6YlqRgoX+3Fo51h62dboH//6D/FHPx67/jnAFbceRuRJ3QfbONHYszRVWq6qDP+j
X5my9p0qeo4erWnNDKnn8d+pnhbkuHi0QKMmiS91UEs+ZWnNVlelpvgp8vYMGR7Xg0e54j4y4ErU
QI2sYtYdqsjKvCcoBxI9s/pw22iEBN0F30CZb3Qo47mBCGYS0Z7aEv2jar/zkME00F4Bgk2XODx2
lt1tONKh9OQC1dN42awKcCAjWiCEYGZV6WlbpghV5DbQWeOGErHF3+X3814uBlq2dVEjZBN8ePga
EnjTy2hHv2ATKQGJgo/mNm9t7+zuaNgtlzBQkaA7MghbG7ejj8K557HUJIBZ1206t5t7AbceHs0r
6fmO+5pO+lX7pi7KMfrCcsbq4qbJeosYNETzjfkHo4rzlqpgPsv0CUMJr8VkR5L1Q6X6J1XIKIoL
g2mQaS3QHyTwAY4fUyZmgp7eUrbird5Epan5FMZKR0Znt7RWyJb0szzAJ8iTaLCV2ZeDAMio3G6M
scC+1NS+rr9G0w6NjC3nbVfh0u8Om0qG+L75GKisqS9qPbuMUKukWaZ6QGF519mNqNvWNTbBP/Hc
zJBfM6kPA4PDW1f2BB/0BhbEghwyT/jeinWg0zXHWgU6zCgskBO9CmotSFN2UFYWh46+p2b4fxln
NQBDL/YqrmfBvLgPrI0EMqD8hcTQ6BG6T37fW55rOxYyo4/GiTQp0TqeJViRWsBrANtQeiXb2I9w
hdVn23URxXlu0EgcQ5pvH1/tPnsyTq+v1L6UNEqCJUOZGS14J9xTKnPj6ftkPcs4niyZwEttaF63
JRiKkgDDl7faxrrFI6C59DXCwlMI4yOis+Y4+f2TAsoBOo/dxxRJ3xasFXn9dfQOXc1xah1Ocwdt
eP2lkrG2nlJh69ERmhVgtp0U4GoboluF0z2x3uMd88B9ghViuAxrRcokBi3M7qYD96EZrkCVYWMs
4MR9tnuZuYIwshoYPNfx+slod5TKG8p2VyW7scpm5UEevVNiAypOPm4XJrPFtMPAgV4zuX+h2+kJ
C3tnd/sknzukHbEV+ctpRDJpQ99VtZIatqq3iL7iLezfXxub3qpcME++cPQzIs9/IuiJzRqy3vNG
k30I4187r101rINdsnHH68AWRpXxdD/usz14rM6Yrtjc/Un/GsopbYngLY6p4lgaasRWzm6jdxr9
dZxydwJntOwTu39pteqpWP/g0jBFdFR5ZgdAOaJqOqtyq6CQ5ecWm8kSpCTWUYM9WNQycopa4+4N
nhkAbe9oslhO88mLm7sgF8Ey0M7xFwddKgIApIL10jEAjKL7fQQmeJ14+VIP1aPdiNcjuwU+N9Rl
3zS9nfwKEYs0WpzDR1PbwFZT7Iv3aXkWdZHERRFdTOlRepHmWrkZNR/WhbK3uw3Gj23D8vwCQ601
gqizNnsobEcmwiJZnp6Tl0bZd3bhTFw23fgOrwlrN+j4/5jrDbgLeqrJgKNOsltIM72eP80QG1wR
MSPY+m3KBIOaZTUnTV6fhIhCmQnkGBKw6Sp+0K8Zu6AVLBqRK+MkzdasrlXCNsbvuofn5yguueW3
dMB7RdL7ab4tKH80PXpDQQA1jw/ulgv0UWtjhoY9aqCfdwMjzgMSJ3bel1cb+y573iGqIRIPtL8z
p8sGfTXT1+2Fuio1FsFcavGx2tRDzB9BG6jY8yI0v7G71HAAgqn+FNmWd6v/D7nre+ZIgHNeHvh/
2sXbKqD8vZVfQmUVhZz7it0ZUCj8k57iFo3ooz8IWRWAR/SptzSn3BGLwA5dn1wfl4ZcfrDGiy7c
FRk7iJmqSRDPc8LDUl8jTqqVQwDHLg0ai0TSBemo6sD25OZpdUz/FDQBko9d3VCcZVtQGD65pjVg
sBTUK515AWYSvD7EvgVgwIwroWFl5ltOiDFR7QRee87CrUoKZCQyJQ4ypcAXiy+LDQk2YnChdvP+
7OrDiNkO5O68d86ddyrpzQ6bWIz+MeUAxpWZ5kYqgQY1iDgPWfn7Rngm0SCqQS3EJuasjSaj+soQ
ptxt4mdSUBY7Cdrz5mJXZwlsCJ1rNzPWmKu0b19tL/Oegh1tksDuAuIJBoUZRsXsOAKfDLKyHVDk
V1ALPkGRtFBjSatoCZAzKN76asbr1Uomw3/DSFs3b4iX+MSWPZ4R35XPA90HBxOAu/9BzILxHO/9
174EbWkfFmL+5Y8RUI7Y0XzZ5gVHEFkZ1WUBukceIvwQQGHfgbJPpM2G8ge0V/cH1pnxwOwgbAiP
WMeIDk7DdM4zijmXCQG1lZL1JCLxfe+RP0qdUMsZWe/4/tZ3Ilm5Dt8vCMuqkNlxpvN+0yjOZ+ZV
PfBtL2nMypg0xN58yTV9qAl/BLv8U2wokh9qaUsdzx5kzKxmDXP5vAc9Dwvnr5w8hRXM1FGad8Jt
uasOQ0JdMlXW7obQPjQzKEG/AWvCn3TQj5KjiNFUTbvhQM1KMg74nftB+nEcSnrv9NsJz8fOfk0P
FxIFaeOBwzMa2NsoARC5VSo/q5og10Fj5vbtkSzkZgftBiMb0jOP3BzlFIoCpnozL2HCfIcy3+RC
c/1hoHB19bMVt0M+O1DfTyxBM+yAdJx4D8HGYbl1UlqcX9IE8OxBEvLVAphmIq1YL3hgbOXE9a0o
3Cokmt2yvYh14wuO3G6ElX3rXDDJVCZKZpzafBtI7R6l+uwcLKH4TMyLLnHjpz2x8YSfWKlY1x8w
VziBvslzxKbFQA/wWIFvjqe4VZc91Nx2W+ILlbW8D5kvlV4J3dpQT+Ys3rd+B2ZgIPOAyr62ma/a
ReBLIuv23X4hz5a9/9NFOO6wAre4xw3LLPVut3AlHkQBkkwOgGl1OIeTuoaVGvVkTj46ZRwLwW6z
2j2WvxNUN/VUETK3kgodWnzXnVFisN5gCpDZ1q9hIsUYTWqymZy8WyDyI1PM7Br1rUZWT0kzCge0
lQt0HMfAd7M+tawun0brO321BkSmkt/3A21BmM5D74dXUIsXczt+NoCNhedecEVTsF4mwN62G9l+
9WbYFtkjrjlbxVEjtekNcfP701+ZqG3pflnkrUZUtJgYWVLgMkXFh5+IEcZzNOX+iFQU284kIpr3
zSVuvHlbT2VvMcvNl43kyef5or8x+4CYKuEtp3QiXqqdpBob1o6AL2ToDi6xHdYAT8DnxtbFCKZS
M9peQTbmjQvcdykwz3XfqyFd4G5LAWREvlCJR0ajmAKu8EXJMA94b6+YGCBsqnWpeeDRZ/+cd6eD
5vdV7qPywCLfirZGmwSEgzw4MMgTLx0FUcPCS6mNstHaagQtTJHtsuM/loQiqcHLE9JATy2NzgM9
y0b0OSA/VHMJ1kRwDGy6Xqvo2OUNUM0PyaAm3i2ahNKW40YIZhgCiRjYufXHgfZD/X06O4zqQLK8
RnovcRd3hY8JObZMJZeM8Kl1KPSazjoCtIBIuyiR85kVQGxfNSzJlBIjeRrwTttHysCfM0P5X3jD
ZDJb7mWlKahI9A3Vim5tYO4oTvkMfWyUGwPB0VK8n31EqKOI2iULF4mupvaAUJ0tX684Oku72Dtq
MphBsTw60as2JoCD8ftWwB8whmYm/6PucSLCoTNTPqMPHJUiN3TrG0rDafA6gwy0o8sB0SUWJ4NW
UF4RKjQKHXOy1tEOXwzPitzt9UxpsuxOpWWxf9Auc4FyX3Y3LqQhJypdEvxG2zVA7dYLjTBJj7HP
0edwmzg7FAkfMDT2Yfo4eAoY9kFixvxj4D3IfxEx6aIM0XBIuHwZtexIUrV6nX8Hcuh1whGd4n3W
MDTwsf5eQQsCxY8uijJLXEDmUs668e0bR98xdl3SaTzwgZVt6g9p2lb7Hz+8vLtBbCvqtZZfxoDN
S7ctrhXYpx9fNs+zp6cgWV1R1jOlCjCnzekAq8SR1hxJeFOF1wdpn940JfajAGKZ7Z1+RajjES4X
H1V+pz4FkkzT8y/QNOdsuXhF4A+5h2ri2oiqEhZpDf1vJut7SVQFZ86JApBzWwk/2TePnNkQasVA
/bKv7+y2fzsuOAWQLfXHOTbaUmFS7x1jh55BwOzka1ECMK6oeIPLx7yU6XSEma0k4gWA7M8tljcw
ZR5fnBbnbIjMnzAa7avv9iEY2GC1b2iINtDoGmcib9bCvZakphx4xtY0l+jPgmaLrGK8TzOki/fA
9Ft7rK/IemSCDfuxO5M8yT0OVJ1xXzTf7V3GMM6CZ7A7kwWEjClE/AmNG4iBDwtr2a6yFH0Ho4IR
f2LuBnLI9Ry4Q1rRwmaGCxXb0wf0HKeLVDKPhVe/Y9AxYGRTEFzKPwzzliTPea5IK3Z6/FeR2QYN
D/l6EQ/fK5zIkvcSq6myl+fNfDTg/Q1+lgpdjbkTvr/XBWMnMm1vACwKiHR1UmG0aWAXqng1w5uv
Cm973GaQCWEcFo8dRi55oQ4x/nwMkPUKvrMjfB1QYpwcNxZSJzvo1azspS4xeuJiK3tTt/dFExDJ
1cA59dMHeD44hFKjFLIyA/PHfWC2Ac8vg9TLBj4iC90+76N89yN0PoWh/dq5MNroR7JjoFcBqtGg
nE7NH/orqQ3RbQM+Eii5PohqOuA7vMagaKmW20wpj3XVuUcBuVzNjt7URVRCW3n1Rrg3syNAfqA9
gfKtqIZOB3xqLaD4yEtBwH6MfXZOLeYA7FXxpU6tNmeMvh5Q979H50U6GRhVL4pXpNfh1om5TzG4
kvb8JGiv+yQyi74DRxT8oYVHm+3E9xNBgWGPxF7jIlFJjf+gp1wPX5bO4k0xwzeRCjdEhzGUo48g
fQkps5L13jyKRpNxVJkKtzNe2xn8E6Bs+6SM646xSeek1SG4WeLwONiZ/UqhnDxEWydH7jKT0YOw
KyCQjEJ5243br14aWQUaAgGAkeTE80V4Yrb69MNUWGPGCGrrc+lE22XiGgrSg6+Rifk6hjbk6iBl
cqfBOC4b/9QxxLIOr5vyNKsbHJq8E+OlACvvkTtEyrg3L/bhOfRn3QJD4rps4VEWkrsK1/Yf0c7B
2uoNoioeT25gsQb/5p3uKvQFKAqlDKQROmECB/a88HlucWIt4bXa+4Yb8g9jS48tsvzH/6If39cQ
fuRIpcOBJvZx55ls9fbgPsFJ/3O6cHCeGmxa4rR1IV6pkBHdHLFmKTQe9ejt8DJ94lm9Nd6XYyKU
hXUNdCsd7SAXbm4yqJsll0wyuQ1fC1h/KOLngJmlgG18eu3kIA6VlpSDOARwC58CRicMZitsLXzv
syzS+axuyYqoDkb1rO7Jt1YfKmzD2P0Au8Jm0CEAiUvXIn7E+gM+y6ggQprpq7B7BUVDQpTU38Lj
aOPfI4EL4iu16ANce9j6r0yoWG+DqVLlp3XUOIeM8sfDrPcdjw1l7WeaFpHt9SQngKtdeGe/qRjY
GnxmBFGDG4tKkF02Pq6yFVZm8TtYtnJyI3p7mOUfnKSIFNw0xcrDAJ0J1DZjIiPNjZWAa5YO0Ao4
JowkAXnjwkw5Jmf0H4mvqs9kgaR/dxJjIm6FqVqUuJ5n49kTztjv1EqOuSNCz/7ZSRmVeHErugMD
BO71Ha6qBR+M3mKkWC0mL5XV2G+2iOKi7WEuWRhDQfZ9xaECxp9AxuFm6tf4rCjsL81Ump4Y1jSc
DhShSvsRll2TJ8L2dMcExEyZ6UBadekWev+u7SR9Qk96i2bdVxh5Y2IzQE7ZYiWaLMD9P1SeBmNO
hlEIUJjCBnEtD8RfJLSQ6Fiq1FN8D4VFJIzao11k+X/8xHEcrmJmbw0qBLNztvffDPFvjVhKJmhz
mNIRHdV0qcSiwBttHu6YcyP6Kx+/AXGuczVqvQnuKyuK2obVJVXTUXROh4G4Y0NtB1lgRK4nddW6
/PCNf2CqZgR3KOfvmkP9UlfnJutyVkZyyXEaB1NCIq2zcRORLwa0nQ/kBgqkkJCnijYICW5CoB9f
ZmVCZyhGZQGemdDK1fiD96ULO3Py+6i2RNVpB9tCRsZLPBYwX8sxRYc1RAIuHS/iZMJjdfM1SeJ0
oG7VDP9ITSmcDgYE9X78oyzGCQw4mm4PgBBEBKGQMiO7MRxS/4z92M7QvimdYYDNkBlgZXgf2jgG
EsuAeWWkO3RdUcYB3c00J0sOgewGFc5/SfX2hO9mJHmPaPhHbh24MYzyT3hFY+lGQ66yUoVHHU5a
no5EN+2a0zrlK91ViYa9DQmwaCzSKb4jneVEO37qW2k2Yxet+s9k1PrNKbMvhUp5Q7RkPDsiwUpy
R/0rVTl8szl8ZZNcU6R+Iq5DmaO6IOMFzy9rDlvlJHJIidG3Xg0tI/TTbQKdDMznz42MIIQlocDg
gJ/Vqp+WsjbvLsvkTl4A6tR9xvRAqiA3hFgfzHRuruggJWCJpVXb5Tt2HvBDqdeYRdriOMjyxAHh
KPBY6eJlIHej/VgESUiQ+1WQKoOf8XlgWSyNGvOZYJPeN+ev/JyiuGd0Y9XrxCcIR8ei+9Qex4g8
t1JJ1ZR+sZ2PfY5B/ppBBIh+M3EIqFmgNGyGI6kbF2JH25fozDUl9rR+b3Vqyd8euo4fvYzqCL+2
87urMU180ikaOd8Ouro8TBL1Rt/s347PH8KT9kIgffvQq5Xs598YmI8POs4IN+lBgAEkSuufR3UE
dB4vVDo3MiAPOjoXLJvSyfssDOrqRJ42BNJb7owy/04xqSD5xOvESwv+qskxQwjDUFP+K9Bazajz
NGnZ0Ye0jEGeMU/bjKY+jo65pr9LMs0iQoaRwFtReF5EYX55FJLgPt3zh8mH3wxjvtG0xnQRSK72
3wT6KUND1os3YRU/pFg97SG03tt0izQ7EEuaKZph3jiNEo/xGh07AekcE8lMQ/DrRFRm8BOp1yyO
reaZQQk+YZlgA3/u0kmFPKl2QTtFcnTBMkbeNDRIDFE/cvNoPTQaAqmpUwv39dmnHLJ6vuSAWp+W
icbUYVrB8iChMeGh8VRwOSANMDDwkOPnlzWAoFUYCDKJPnHFOMKGYuM9kZX/ziGrkdHMjZf4FHx9
rrKnoB5ccBxLM/lb0LLURvgGpb1iS6EbjTsOeM6lBGpUVNNHUV9EWETeYiptxoJTtb9BBuysywOe
fxODFskNpI3BEbsB5JzfeSeHptak8cWa4kiMzh6mHT0NvUlIClGlgItI0IL0hkc8yUd9bAXtCiK3
+r/ViuAoPvDfDWOkUjKSnhz6wsAlzOK/nBV/m9iS5+59G0XxRvUb2q16oljw0PSV797ASDRKKSQ/
7jl+WoZSw/cmJwMMibBsd44kCIrOkiHzLvxIy75brDmS9qT6kmivQeeSF89nz9m4EyL6IjF6qYr9
hRcchLwUKNtuGf46axH/ofxQmS+z2KkFbYgp19X9AvhwW1cT9kw9B7ctwfa1qdMri7vHZZk/SWI2
UcTi3bGHoen9/Q9t405RSm9Y2x0c5g6IVSdX3JUFH1bhCGEX4KRdHgmxSeu5aZVgH27xhCnR/ov8
3zWzHd3CaiA3D86cTxFmiozTwqVfZO7Iz9Sj1V9uHMf/J/B6Tf1Zzh3j4vPMemVUICDbVsf2dk0R
R77lNpcwEBQYwTxpw1criyKPGVH+KEAsRWKD4d2KcSHT6x6iTDDxgu+uivhn/AwIHl7z1BM+xswy
YKXjm9ZJNDXbHM+HmMi1XXje6SuWadnGtc7q5nf38f84PJJAh3UjvU6Yh68oEtEVrJC1WXBgjfpQ
FMnq11aUw89+wIj2bkrjJ4/rirVwsy6EuDADXHspSGstcOpkT29TUSfWHEpp9QT8IwlZOwhYv6RA
PA6xwIAH8jDm8rVgTyW3bbzSHYoA63Bv6G8quKjJdj5uUHFWaHBuTb83AK9GBuV9i3UF5brnhLTF
MT4cqpUBUY8kxyb4IZEaLr+VeTta9e+RDwUaeR/qyUSUnSI2gWvPhLQWLsgkdVjmk+9IndSuc1Wm
HFVsqcQlVmuqCi2jLKT7YSrbv0VOdKhN62zXzadbdIMPrzVN9JJc1Bp+ptlGmLnPIfZKgEExGmgz
VMpYzhNKdJ5/H0P/GpRRXKf/UTlyXUl2xWzuU1cMrYU59aKPe/M29H+vYu/hKzaRa4k6hqTjmzS+
8AnpY3uzCT9eTy9zCI9CITBhIGXuDB4i0AMtyW7mzxRh5LR0fawfGmSEaRVIWGzIsKIzdmcKa87w
m2yyehv+lFoby3AtnVJbaUotQ6mtTNdJT1hSM+752wyTzOgsOKAtHaWl1tB1Fd1cMTfESvhSb4qg
0TmvDGu78u7FuHFMx/v8yVNULHrRAIHkps6XUnm5BFpDUWQ8C6OxZ5zw8DHYKsALleSwWbxyQMb7
tMdCI1C63AdI717u+Glyukl0231V08Dbw+9eAfDm/qZK8HujS1C4mdM+BiNUmi1B6q6Rgvd7rU7V
o6NggLQDRqxmgEpJpGsUvgBum9yyFyizZSGR+DStf27zOtNf6LGUBwqzUI3WM5eZxMT4U+I6Eq/U
wYQ8FdzulFCUJla3Y9Qrepwg5j+X+as7qOERS1iFwD4PT9TzGI0JbOKk9yw83NuQ+xy5EdpCVu2x
rPJAUP9N/wMZ9VyuMzPc/qTZhTXjiMGLT0P8+0Bah/aycbBJNfWoBDAM8KhD9QucXKaCqSTzWxDv
u3nK2CC/h3MZrsZKmypL7Zec0HlEvl6DUWvlSYO91aE3FRyxYiISZllCXSnFeQxJfz+LyWRfAFmc
o/ZJJ+QwOTpqh9gZTswTVIAPY3jN883aBhXALEzNu6lA1lpJkNFeI4O8eKXdteqpvzSiYb+HvTRk
FH4+Mo2xaNAowVMa2Q6/Jv5SW3CwR0Eh/OXVEzBTz2wvDxD0IG72+4FZBHQRMgFuHMOpXwITU/KG
VH4HCF82xrqHJkPriE+YUqJJoL36eDYvil3M/GdNwXyuzLUN/KBT0sjUbOFU09qI6Sf7Z04bBYZg
sqMdF3HcqUlx92Xj/IV/nWHllCx4YTxpZbuJbtik4Yk0T+aBYTDkt+sXpqQ0XgQxj3p73Nmy15tV
Fu4staK2PjODQsy1JPC7FToVVmEC2iDAEZcgzAA2iUVE64h2AgS3jFTPpQ32n2QTmFnI/+8fnDpT
HAwp/nEjZgnbIU+49UjTQGQvJWeg7RVspJ8bNHw4kTnSCnDjOdZtV0Z9v0746pgMAJyncONNuEor
wCXGunxCD2MDFFTLlUi3U44bOnLWf+uHnhoz0XrMPvBzGPSCt2XeeOWD26z1QjXqKQx8r8JWneYs
UtbrUvmXQDizOvnBPLienHKwrO9F3Jm+keiDOaW5RZnzE1afMxj+8XXDV2Y3lrx4lGVdTuGkgATp
GNjssTvLMvzsey9dP6N1UtC8kCcJV+yho7DQfAysAU+ZBDBFrcnGzcQUjy0DH1h6BzXalRKjjOQI
yoe8WTbz69Xk7PIzndWhgvD/a+YYpDNMSeuf/L8MhP//wfl/MWTfH1M6xgs3LhsDPU0bsUIBtANY
DbAZVGTG6GIKGXQa/fEE1AvjeM2SyxZyZbgO9kNqLsQ2qhRUt+JGZxVEW/pTktGBvgpdJ1gUVK91
oAPLSX9Ibylb0HTxUlCgvgpeEEro06L8ta+ZvIcpFlWTQBYOHTZTwLwAkC+I4CSBI3hiY54yfGiT
8WCJwn1M4wCfnmKIKeeptBH+XNNnRfurNrVfpcSl7GZ5XPswuXYfqsffW4W8vMADsXBrx+Q9GtzQ
G8SE+tTLYXaY6o7F3MlLXQoMJ1lgrv9zK6Ak4Yd/WUq34w7T4n9ttYp3U4+gIc5795g+gyxYD9Sk
hYZP3QGfEnPhuynH1/glDS9iDX1YwpvTXCrD4No7eMrjfWpZTtQJY1m/h5Iv1CznTwTDJVLKblc/
cEc3xU+Jh6XUllp3GHTsXkO6UOrs3MhlIDaiGeES7wEhaOyaEYSR1zIhxqddMrmxceTyHFbsCLjd
cLESZsm7DcVXWfKc4l88yjfhduB/1K854HbFjOYW9YfQmG8rK4//ikq/orD7zImKSpT0X54ANNNd
I8b5ms0rMD4rnGfqH/qR0dw08nGJ3yN2HTgIFwjy8SxcuN+4CSO7nokQnxW47lFR5FgwwWB9WPUf
pOwAJzevc2Rho++8Y61nFx0unJ5rq81fE452RhU8p5pMIzfi57oVFv7BkCIjZCdOO4xmcTp5qiOP
XtGYWFSWNUvhgV1AJ41G7pe6KFpdq450Y7m71rvYPFZOBn/Kzpr9HcgOn0bTtqa401X3p76jznvQ
XGkIRfniNfyqrkQxNIjCfD5AY11y95/5v5NAnb9bERIcS7IJEFtsbvu1UaaaL3HamMYsABlfGjh4
aNHtSPpewD5/Ly+MuPxDXQoVMRIsb20y+/z6f5MI26wXXO0leEYyGhktzX2b/P7oJPt2hXRCHNeT
UlZMVgGFhZLFS+poD38OnmtnbptdvLuSxTmr5ibkUzhku5Kodbai1SP9qvKdnbKlithkq3CtQ0/E
tvRdybvBvGYKKkptOYOOoetqlBUs99hq4o3Tz1B9sbMG1kypPUeMxUeMxGP07x9GiUmUsssaa53Q
i10mc4aKjffW/OVjDH2cU/o0rhIbW+DUih6DdHUT3p9GSpmp3jt0q12ywD9pfYBoDtkI9Z3FTlFI
vFSrj8unRa7WE/DMkKFMQwcErQZayvRRPvWmdQczfisdDvm9L8OI74GPv3YFy1YqlODLBpw2eHcS
3//1V5sUuI8iQwR2gWwL3zaBB1UqIvi0VLzFXTERQkcQVV/g42JwC6279TkDGtTH4wVX7iRBqong
EtBhd7Y0aBthDmIC28aUmSIDzV0SK+HhEtgNiWPlUZJ6mKTi4h8lSQxa2y7qlkV/AojfOXNVbG04
5+dli6N8xazsKfZDOvKfJDL4lY3CCJH1WU7XwGZJpAzfZKJz3sBJPSUyyAfaqSh+SCo7jWONxx+E
u15ZO07CS+lQNh6aeFeQxtLRdDnpO0mpe415SnRWwKODyhjdzhttWG489abbUWHmS/llOpz0ZeCZ
AHxIDAGQ7qylYhWOxqEOJ7ObSMBBbTZhtQb+x3jpZPJqO8VXlc3zFPE7TFYmRSeOMhBIgfC7M2HQ
QbYLJR5O0aeALs0jkboiBZtaJbxYyQ6tuH/x5YvfIz+hOScrW8xxxI1veJTw201WnD1ueuImX/M1
nXHJxwxXeo0h0vaabYgfrhU8tOJcQAq26tH+3ZasFWBXd2A4iii9DE+FHWcAxWimiFhQSTx09baN
BUhlJok6UK+opWHhH0g9M6PymLjJDH1KMNQfBu5OD/4ghh0jw7LDymwWh0yu7VwzIdrtTUhnMCfx
KwuDnosqGLzKM3VlZj1AQCxpcvSv1fltQJCkokl5OZHY2qYcx+gr9gfBvDYQcYstSrG4QPxWtu4o
poWW1NVF9Xuj/NTbDDWFUv+diRnIZjghsiN59CYL4mIzd6VtQvGvfYkX4/VEVAnOwzmvNuTzcnUb
bLpKJ7b3cQVoez1QuymSHZeGXS5Ma4fQdjEY31G5IusZMC8UdLU1HG9gCjCtAtRumWnP8jOalzKY
WVwIMCzP/rjFh1WjO/uBUDhKzZDZRh6A2iBd/PicVI0ZM5VSzsHEEHPO2oyWTiXSpi9v38mjQ9uM
hZPKwgfhLrcthibpAD5xEvA5TVWU94ABF1lse93uCSW0Sc9OPLmIaz4Qpbsxmw8gYUnEFdwoax/k
eafUpEaU4yNUSsgTSgimuzf4/URqfxcGnzsRo4TeelFTL9fEabwcSFOKuErdEY6RgVUiznRiDJ1L
Le5jOK8iIxTzfFYihdNBP1c3VnyZP8wDPwib/XypEvQ0iQl6n1dzQOudktP7kLXAw2BbZ9XfiRtJ
iMADa4jrevArcSndr0v9itn0NGWOYv8Q9UVbMqJLyYqhacVSy6zy5ZCFAvBDN19QD7yhhKP7Sp+0
DUedsQw4YHsiC65Cf+W4Yyx1bWOYF2N7wdn+TpRwQ4dk+GnXpwuJjraUAEo0Y9E9xJYtbQa6/s2s
P4bhiJtyL3OZebYXheWqNr/Sdm4NJ13xqWmIwAo5KlYxNfPFvikWOnj1D0vbWLR3ePd40xbKVBxb
Sw5zLbmLHO/EQxf3IChOeOMwSE0AIJP34k1VCgbhZoKYM8IGlM6yjkpRONPQuQefgoKoBn292RaA
wqHauahJwON+cqaqcqKtiwgRXRj3CpIv6Oo3oted8Oy5NlGUGfNJ/zOOcNKv7+OeCjTl/bLSZsJE
NEdeX5S9iKHxtN/JbkrsD3xpAMrocBUnguBbjDt+/bbQ4ko7wYsjIh4r993hoVI1NB0CzvpUh+GZ
HnyLg5MQpNclJFXOyeG6rAGGUxQDo0sN9TbQ7DR7Ox5YsmUArY7DtYqGvrsErPaLRFScHxVGP3Wh
tJEfsqaXbHZNdgd4JgzXb4gogU7KJcSy+h4T5tV/xXjvMrxbuBwhoDk3PVJgPeTkOulWDuX4AUwl
pT6O2FTi1ZZzHeoEc4umpNBfZa1tg45Sbk9aOd2s4DBs7C7hIYXO2zJzESg42cGwZyitZNtBUzWP
RxZx5gxjSd9kJrvCTIwL3oLLDyExWITLw6R7znbseAdTbbvnq9KDD3lmj+27jPTdoI0wJHGaPkRN
tuUrpVoikbgdJl5D1o7xllI6Q0ZaU25h09oyYK3p7BFCrDBy1dszmQjXRAz8ra4H5u7W4Gp89U7Y
9mhbKhKDHfOPpxfVFa/2k5AZ5x9vGaswvaVRlylIFYRUdUdc6xs/y9yCKuA59x13efBVrGWT/FyC
/K2x/0AYs/DJeJa50gEw5vnoW04rXElEI5bxKgHQs6oPc/8zQqSFglzNy2i7jYPJa4U4NpKzCpzh
WLsr0ulTCBXrVQPL18e0m2JDUUSLgag04VMlZ8mgnwRV6YafIZKhIZby9olyc5VK+hdznSTMHKNX
Ru56ClIktl4cLhweTj85vmFLq9NNFgYRPYygvTQllB7jWCeuS+8uMDgrdr/K14egVZg3AD4lm1e5
5iLMgOJyB/ACEETmbLs7ZcxNlZFD8MeCZWlx4CUpkbBruqCiLMWAI1dLxHVd5GafZJHq83ou0CFf
z+DZ79tMulS+TuQJBFkR1cLHAbUP0cBrH+QIhpViNE4DQfnoSFtioLrSb4mKXJdb5Ki+ltefdKTo
1etpZyIVr69x4gsfXwiYcQ/2skk/Ev6ils97kEZPb2dappQM2mS2UvISPqvo76XgseGJLmoNiECj
r9hTKoPOwqO5n0cRiE3m8DxFL9byaILW++SnMEBsKJ+0SW69hOnlkvQkJlS7rYQ7DnbHvvjAX+bj
++hFPiSFBUopzzbbI4vbdnZhlJjcCtAlRsIR3LHsMnnxQmJkspqdYj+YK/mMN8f3hF/i994DTq1t
kyZKjFaabDSlokpKhFY7wo3jPEN6m43dlOattOfVvf6SHZgAFg/RnBE4OgCHj7zhFmH4JLdCAlmG
34zGIHcZnfVX6Cfl9zh1p4hdiBTWC8oqY4eP1JdxBTGMKrICN1LF0egtnezdnVKLKjP8zBweTf1w
J/bI0eEJYySBZXxZ0fiAEEUtEfDPlpgBLdwEAOY9r0HvBP413iinoo39qxBl5jEU51ayW0vtrZfv
2HhxmMfsq8Goa05WMofYHmHOXRjF2fl2LiMz1YoXPOSbKoBfjRrEsSJItNAOLFNG5cJSSFSwjAHZ
MHwEi1JwT4gkGEdaJYSh0hVQL461/uzEbcXH+GMIP7iqyNjXTg3b5cE1MBtejv68P0MFzhR4LUFE
1V8C2kcjam+gk/MRdr5fJirsByqv44oc1v0gy+Pa6xTR9qOb1Adf1RC6FWOBlX8KhiGSr+1kmJdz
DcALuynxbNArXdKwRTxPoZDM+wSRLyrvIjVDAQTAXYHrwyBfqkNPfFDUR8BsnioKHkFV9ptLKyIR
VgdvKWcXUIYygyaiRw6VjAOBrDgD5POvS/VYkOjBUfBED6R45in5wYeegJZ8Lblu51zIq8CteeM+
UR/qEMTF8j7f7b1MINeHsW7IE7tz8uhxTcZ1lWN5A4mTftIbetD0Q5qaDYHNpKZIvPLq7H6uYjMR
fRJMPBqQKxmh8fHfzVT3fo4EsFJEG3R8b4H3Cnra0jfww1cJfNVK3khpwX+xTIfX2H8X3QnnSE3d
Lr4zXW8fv9LdPvNcqowB3YLyyj3Se0Aqp+OtVPna6G0hegL66Bf+FNHO9TaRXxLNHaDAotgE9Tck
wItVQVGLH0wwM14S22C6noFAFpl2b84t5WSMdtMkEFFBPN082I5xp3wS3Ejsb6EqKFE1cvCrmUq1
M5BG2yN2BpoUQI8SUvQhy7j1E235l9poMtttpvfQlorTFhUkJk+ggKRr/+YXrbznouEzL/car3iV
ZST8syOJ7jnkDp/4AOST0eciJ+lVQj7rhAX+mPIsidw1JdVggOkUoFZnWN8YXPFkyO1c7Oi2l79y
xgmtN/xXFJNxZM3IrFa7QKjrMrpVRpYOCiygFVy1+WbOqH3vmG6tTuG5BN1ieBt/srlB4uNnk1uv
NvNuqP9WqqcQNsyFIHGFeygXlm7EeUom/usP8/VGIPhNB17He4wXWxg04JKK2WF40cWaFEufs/wb
2M3xfp8cdUz2Bi0SIiInowtR575Kcl8uylQBropIXchfQ/v/gX5nCXdTh3wXwCiaqWlGEVy5m7J1
JmWa8f5ifpDvZSNF1vz5QGWWt8WecM1uecls88ZXR02Yb9aaG9eqHrPkJEi9VbY+9j6tAIxPIJDp
RkAsRsYm7ZhnwW7hSsQzyyZjXdp0y+6os/tImV10Ddgy03m5iBBatWRUyLsqxvw9943RNe2mlWRX
/yyNiXYdAp7yL3HWK3rUzQFLqoeWDHeetXZcHhpoHFedYa/qlrSdfNSXN6jvgE94wrgCbymlZW0P
5+SMit+kfzKqc6fwmZhlC8IaAShKVHOVvFidd6Djg84ndHMpAfCN6aGARikVGH1T8hmQjjgHhaV3
NRUzrYUMF1wrei25X9vjD69VyRzDLCxi0S5kk+SKtcjGHpTnFteqOSph5Acdse6M8/oYTqKcofgC
yKcxMFdJlPgXe7MncfCGD2AzRobpZEoUgquelLNp/OE4N+av6J42CpFVC36Hkq64raH6k49AistG
Y8A3pOaib57T54wBeJlNLTWXX7rLQvxcMNRx6nJcfEFnAV2x0N6kWZyDIjGu52bjOcYuvF73sdqj
Pk3jWMYA50xhMc/Cy4oJsOBV8kUBYfpsM0Iq4pgz9KAN6/wrUyud3j6qPCPa4SUhmUjHR0ho+oD3
mbyboTbqzKd+5FKwQIKtEw3JTEhcJokFw14sLTD9W1Suh57KaGFetyh5BlbteTrfcf6oN9O+FB7D
VYjr6GmctGPhhUpz2An+jxqGHlz4JzcBjoksRs/cQ3ldhRaSmigolLPeRIAx+F5lsEuc0gx1ADGr
yggYfNWD3Ll0wCbvwG5e2ZePCWWnmoGF9zSMef7tkI5d1wh6zwtbN+N432ymKC3xToaaHNYVk42V
MCWDeRoW4AAp0lkFil4UapVl6lP58uf/WPmixdGOyDZIfHGMEqmqtS1sKUzww6VKHAGMiRdayOQF
YauRvx3W8CGj+pK1aFsuJiN+yxXgJAuf6KJ/ujEi1KTNCqWixlnOx3txDk37jZfdnHcKIiKxktdq
2KHEIuBL29TVMMZ2ZdVFVhD9WkouFJSmTLM9x3dU7uicHQ0qcv8toAoxZ8+RR7vlWjpCr97k0uYd
dCHDT3jcyft6QE2ZRqW7GvklZnN4Bq4MIIL4qvWAiAT4soUE72Q3LwKsXdnaJla1ZaBp9PpR/UjD
ZVC+H2TsXMxMQNUvLv+OwkI39rzTxT5n+BMtNbIaioWDuSV8+6tcDDFDb4JYd1kFK3ZooZDiDOaV
rubTHZNg/ynyMEcS0jmBb/m/zsj1pQ8BjCV+l0rjWbjmONP/KZFTVVOo4sQlWJn4fjvwtgDa9hsD
TXLzgp8ZU45V4Sk0SSkcqxE6+NPm+zhirkxPFj4Byrd5y/H4f2LZ2hd5wwueW1pUbl9PqUdLquQX
taKjOj5SwbAcyOeVinuxmsbP7lW0woJp2AB2aGhgdYT+vNb1zgs+xZD8Cj3QBhtBqQsG1XMf5qTc
RPAux/oCTW6uudM4quvjAy4ZkVQzcpLOFTj1ozriysS2Uz3YFff4TLKiBabitnS2oNmjgQPdbxOG
M8u7mzEQzgWYeKZFOQFs//i3J13tgNW52dBFrdmx08Yf8edIJev9fMy+N+vAMjZrJoX/w0UHCkhu
OPfbvz/m3TCPuHMjWPOKLG2UXVQJVbiTaitRNSyjwApVRJpGWdjIylei72NBzEb9ogPuTddDoMR8
pysFjX8u/iSXxgg6kCjO1hYXTc0bLpeMA+kBo4cdfx2r0z0srnRYG53KzJwL29TE7LpK4bR1ygfz
CdM4aCKYaQJQoBnYTfXA5lGgju5djN5LR3DgmLWIkWVr8dIvFEM8fLSfi55iE5Wf66A/k5RdkxKO
/W9OCqAqf9vJE4bVMg45xmIwVn3z/R8T4kxSG1Svh43nFHVEyGO8nyqA/iaagpetxAsiwqakt5sm
3rakDgvAoGYLMGIJnkRk7iP1RuHFd8MOj20O5xCAJK0KuyNB2uCb07qpQiTQDYQkwag5gIuh0ZbF
H+5++jy/77JMvquNq9ktyaDjXNsGSXMQValdYh/EQZvAPaonvd5p3oi5kiaDAfdluZ4+ly+4Jm+I
PB6iguQK/cyOkUN9MWaPlh0vH8VD3EdJ8RBXvaCcdrFL3y3Mbm2QDKiQpnN7t/41+pfFE+2c0/Qm
r9ePZeNagx5DTM8LBgHj7IFvr8ozJRdUBiOVN82FK1RRUE5o6ryarQ61bKh6lY5hnKBzPEC5FJwl
Ytkf4BI6uUBVTz55t4A88lmyOrwc2sMXlMz67mqyoIz9998IvvqrJOl55HPh9tQhtXqTxIcMPRZ6
oB/oZTGYwjPnh4nXCK36QB3+HfYkXirVVX9dF4bc6DerACPB+BO3P0wJ0dQjlIjBwzwBeNymmGtU
9Dl1O2W6k3SvcRb/xaMXQZE+psEZqw6qvmJXEWPx9mDKOD58G0GKTBzROom6klsaaikcknHp96Ww
jK346Ntd9PF5RRZ/pCb67DSbjiEiNdAAxmzNhgLio+XZYZHe0LYsUvlxyyFUKbR4EPgYkfit2LYd
0oIr7ZF459+I0+iXRwvvSLEU3JzAVjq8BHk0z5YfkzIggfAojo7+p+X44ngNR1ZWcaoQwsPkOrRn
kdMcyqtc16PlhZAfjBszTllbaBG5mp8y+IUZ3/T3/sA/mn/vO5Y7p+rjt9mpqkqpopplp80Di/M1
DqSWtMW7K9IKkRqN/qIZhO5mIjwaUi0nVw7MxFgik53B1Cz+c8FptSecGSxkhnmXv3Rpi2vVrJAo
qfyTRZ4Psg5R0+cK3/rHT/pBuD3uEBcsHjB3oCiaVcKy64Ku75NNcMS4dx2fdleDsOAHxhal2xYS
lqORvTsaJlqXrhEZ8ONs+i1wXYE6fmat/p8x2/Zpx1Q1vlESv1NHHIkKeSWlb1I8Pqd4IjSWttZ7
IWDt38VmSSF+Gi7fSCAYNIzEEOGNJGFRYCggAWIB/WTRG6dIzrO8wjI+5hBEQABTr3GsWyYicNE9
jAF2IZL3UYOhDATtx1+CgceuLNdbHijq0kh6DayrNfLeKw9M0Kf9/2yiRzo0ucYO4xSHgGBqh3zD
c8vf5e9k8RRpLR6wOAYLKNZ2d29upNfnn8jgnVF26hHV5j8rPLthW2s3VTwwFAKfoTyL81puh+Ik
QlQffwhnCk5BVUENN1nZnUNQaWtkhdRRdYOZ3wfAC0LLEvsBeWgnB4egrlhVMJNryq8LDlzIao0W
tkPzh2XYfdab+45z+rS+eJpeSrmJru3gj74o+z6fkCKnKztCV/+y4eCT+ixMiy3FMbRYKnR7FcqJ
i531nrGZYRpw22rk9mgqSLUGDCXSIum2u2tshkLT8O82hAXuw7Wa1Hj1l03Aqh1PNuFgGjEOSB3E
JFGUgM53usUNb4ZICbT2kZ1ptQ4E/fkwcyE6ttjyvcD1XJTXGausNPzya8ELivwia05kuuXQY/2z
riCiAssEv09sdGiSJ+eRQLDUBoZn3yzPsevaZ3z2jxh2UlTVK6fXAu1BnV3pBuLISMzH+vc3CT1/
x6BLBhJYg7mcdFh/fECQWULAUqI3XsOTont4dBGn0RYi0JFePApwQf/T+VjQI58dIfHjyMVPvrRX
J1LYrZKrbrfZZGZi8MF8MjzhnIskxZMpHYTk7gqvf2/Hn8ZVTxxQkw/dTtPsHUJxzhQ05RBYIBKf
2ekgjk7bdf9nI2E7enYvDexwFdEriKUdrpdFXjMUY4elW5373hgU5oj6KifSitUPZFKYIxTqyQln
T3+ln+Nq+tL0xMdrYixb0cb4BEv25NTAA1q/NFHHXXL9KwGVplzBnrC/hdfB4x3KMVOjbvhx8Hxl
EBFN6CiqiUF0lfEREt6K3KzSOJcvoDJ3tZpsHYar0xvMeI2xvKGybxHeaiJgmXMFmcSlafz8QFN2
8XsPDUhdspzPT5Yhiyr66WNQBtVE13TUOKLSorgspkJNJIpS1jrBQoYV/nIl98W6i+lTTj+USF+z
Xsq1fs4oCO6M2qX/ZsalqpJlI36m3Tm1ICBP/p/gzfPtO0sx4kpj3zz+Y92qh+5mdYkkITCdfQnQ
v09780civT56Lnuhw5DDLkOoX+B+yrYzxFKi4L0rgwzixzr95mHAunSS9ycM5LzG9HXn5qs4TM+k
tNJo+Z9SNLCsVrNMc7nDC0PKXYLBOpVNXKe84FFBN6pmbRkW7IDEM4/bivI1Sfc5u2vn6pBuhDiv
dG6rzpTFMdNgyxjTrc6zsTnPuehwI/bFj9qqVXOiged8QQV2SHGOiuzs0VO6phzXWSPQDjUs+dIk
ObKHXGuda630guiKT3ylPVAF7bcsHle8/1fnWORSB2kupLPQSBkDr7kuWo9O3D9h8E/zrZrBdptJ
pUD6SEaty2OHpvSGKTlbDArkeQOdqVEAbn4K1g/lE/rIqSx7baq7k6KVmQBM5Rs7v2+wJReG3uMR
O26lwFjWwN1rL4EYgth3x/OJh2w+f86AsrqpXdSRZXChv+16/NXMi+/xK2Oec0Eeq1Hi+SaEyLxS
20zv9kgpq+qMQRDm1T39uChKwuXW/gcnDC8kGzVCgODZjDeHSYrPOfaS8Xm0l2rc7aDBTkAVvKir
KdQxQ5DSOaf0qnkCANmOQfvrHqAfF1CB6CKjelb1ywNhkudrH9qDMDc3gptkQ4LYpgGzLVoFaBRT
BOrQ1eEdFdBzyQ7pr31GneGbnRhW95Z5Sg0swM+9f6WMeuidb+c3TqO57NO+aSrUqzhT8mP0A8gQ
m4xSHMluFo6fjWwj9u7kn4p+fMNgcEi/2mp4pZ9VoFzUm8OP69T/tUKUCNEzQ3Bf4BH4mIoAaq5S
HgbK7C1QwUZ6vNL8qtTXnOO0g67nV5fsN6a+W1f9gudyOH/xqM6IgtTjahNR2o0AXKO+bEpSSpoe
BVMur1q9XuvQC1RQwSVOcivl4f9TrbTYziW8AbvM/UeqIC3oG+ryTee44DnmrVgFK9nvoo+XoIRG
NJZYp61lpa36WHtV5s+xlvhQwLwui/8/liDjqswK4v38n5WglHMz1vYjiYhqIE1K+wL5cxxrLJLt
yZO9SAkvVqIRnvqUa3KSyv77JdHBNAcyQbV7syE2RlPj00VIpbS+19FJu6khFz4kJNyWA5JNK30m
QK5gkI7gmo2s5CiN2eMhXUbbahMUsPXYROEDwbesKpHATiqca9LSk4egGBXJU/XWaBk+i/jNyUoh
qa+PPYgS0uhgl1pGqVNoOmgPVdITWYzPVzwrwUk7fC85J2S5S2ponIc/IYzjzhHvrm07cUnYvw4u
UUwSA1nGGKT0pkgF0tnSm0TPq8Hw9FjbQh25sUlrW4SNLShbCXe4a2mogw66MQXIFJgX1CYVUtk0
5T7y5F5AkpW8bJai4JjYIvEivxtUmclhbXiKQpEFI03y07KTPgnM5ISSgws1pSnCYhNY5WVOijj0
PV0PVQtKVvVW8fjUAdcvd2w9+hM2RqUlwupnKRspzhPIyEZpwJguugUDmDWnmpZXbdMNESEsd9Wi
ZdQmaJaK+SU4v4yAxLrfY4W8TLk1AT9LMHsK0qLMeZRxRklXPwxIulVtCpKl3CQm5e/Uj8EiAkcf
Xxk3hO5sDZ18SeG2e7IHMbyv00WZMi5BUrxdPIhEapsvGycWN4uwbFrXFRrZ13nNgcJrnD5MqPqY
W9fSbRIrvDgDTGYFBPhvQbzRMmjkYn1wbIVZ+LXtr6B1nDa1ymO7Ncxdhj61o1U8dv1/BuF0fbsK
G5ZsGhryMUxG63zhk7KAjelAp2o30+d2FjXmIbgguaEZ0x1z9I7Xf1AKuC63B+IQppAmrlL0ZlbV
jQuSjJXl+uDlvzi/N0tV3KcxA9V6h2APJCZrWVl4YT3fqvsAGhIR4LZJGvV4ijb14/4/cwt226R5
VJq6MZkhUldH+aGzkkQ03mZk+B/ij2irFFXCJwIE8QkeSwF46W1LEPOJi5M59/RYUFVHj5JEF3TE
dpPzYdHweN/cRg4HZMyq1zP7QWIprgwQWw+9bIa6mvEVqq4Of3sKOqRmLTo8pD5VHMid3+xMUSGa
poSrC2bGsc2xdl6Mbir+JT/uChgrL8MTv5RG6zEAR9LmcVxYrJy4zmkSLoEAGyqcYauD/q8iScBx
T+CVjrrvSZjjZvtkVBpZsFIvDhOXH93s2TPK2lA65JXOKBTGWo8NdiCL76b3gqpCQsr//JN/FXsZ
z8t4X6CMKjpresQ13KySChuxjMTqFzXqmje3FMqiRfKLbmk49R4w9yQ5eeaktfsZ4WRGMnjBmber
MLO2iUAJIHblhdOd80595rwy9C0GIM1L+SOS9h+lJ34dYJuqHqv7DskEBXN9wF6hX42IYptq/6IP
X5oWf4zOF91Imx4MjJDIW4k18y7ElJJLQ17zIy8yOhU55CbqXZxOiY2HU/PWslixWKKJ09/YhlEX
yM6U4DwMj7aeoH4yUrCe2B9E7StQuOxdy3bS1akZOGgqbJ/4ZEeUL3FtfjbtR5+jf6bj3jUo/2HK
9bO+n2UVgooR2Kd21y41qQSaDQHcEZYjU5IdCgPonZ9qQ2nvLG3T0SPZbeVmQVwFRh91OG1MjP/g
0vWBfuZozS6IXQDfQislMJ9EBywB3z0L5wMGOeeuLYjpNsGVjgyYV0a5co1TSBgJ3d2m91hHhUkh
7tPh4iW1KBVqFHA7v4Gi9c4W4HTscnPKmSEKZhbocZRxPFQNAJRDZwWTfLOht/239hf4TBevhRoB
kfj0jawByqi1Uq6i9znISVIe2nwm43pZseO0ceOnGs1pwVheqQyzEelOAVWzj2Jn2xu+jRssryL/
XD3yKv4yvk06LNNCqE5E59jH0e/47pZRUpb56fy9L4isgsURkebKXiJXoSY+6F9lmd/zbLo1dQL8
a5QLYdQlApK5geUxyM/gF9CW59RrQY/idxKDZ1UQweoFyMbAjxSCDX0sCrgi77LRVsAcTyUuurZJ
1oLsIhyYRxfXgbGvU9TnPLoufWnHVLGTd8/78oYyeZBDR8xl4gxNd/Ue1gMdBtldZZJbp4r8E94T
4x3PcfnDAbkO35zDdHtKAi826I0YDucugCV93HoSFdLNJqE2WoQQdUoviIzalBvz8NN4l8IhDZEt
99CW7dcS+oKjpszwRjcD72zn1M8z2fkscp/gTdSVmUmPC07olrywxXjS/Xdftze7eBmECmdeub38
X1Lxthi7pUz4UsNvXeWxqHqRm/K1xm00iIa6lZJQ8c1TmfHZQQ8pBHtTn9vcWRiCn5Co9ei1Y8xt
O9RSjoipLWD58/C1kV2vOdOUivHdQLnvpbwil0fnTCl8lifMa/9Not1Tj7Mchu4SpyYtjQln7knC
KdQo5clHlFd7ckfGPiAZTtFj0e+nXMc7QHXNu/GV5sID0L1XB27nvmtF+gyfKEFMnq7vz9qKnRaP
ZFGmn4Q6qs0rQjnnhaHZZjBur13uUVGsSCWJ1wxGwPgepOPSZBrzOp5NjTDofKCheIPFCGLA3g31
Abf89Ifh2iJz3ZuZ1TKSQUuirGf/dNL/W3mFgxdKeJCWQP7FROtYN3M06L7OJn20mAXmnebenace
jwC3I9kbgsXNo/GIe0aFEXgoRECs1jngc76vDXe3JNdbKQhZ5zLPiOIvNxyrNRa9Odms5UKuKxJQ
bliT1eY4A3FUaJhxWaVoyut8LtWngnECV+er5rlHDcKtVI3A8IQ9yA+KtbpREOjP+aL+0jaCbMXr
OJiAAVSTzl8u4i9HyL4qdI2Ip4/AG6DgsX81WYwxD4cdwx+cxk3qOF35t0ShZ+dFf82YALTkenkO
VDiBsPaqqU5BdBhhWHggAVnqI/1RIcXNptifMBB7CCrjrF4U/YzVcw5fyWV9FkP1MNJ35Inon4n7
hGdqC8Ha+4+ApTXJs9GzE27A8RXrMKX/GxNY/ohtViW7Fm2Xeyz1h7GsnqY4v5bZkZG/AE+Ea2jO
zdH+KflKNcSAdIumuJhwL2JyMlKzlnviVAvGkbwKFdJzAVgVhxdCvzW12pfdoS5e4TMBU1PKduDi
w8BgMfRMZmknSgQOw+O0K5DrzW0PrXqIgmVlRJZ4a6O1cM/vgqoRK7gw0RSqKy7KqVkZxkop42bo
oC/fp6T2M04JSZ9PxMZqlreXWg/tK1ILjBAwPvgug6otJkckA6uT+FJ5wtH+GDzhAOSitUvrkrzN
B6ZruCEqsTD1J0E+h3Dp3Iou4dAg7QW8U8sUNZKT9Y11lCg+5mttzRIhuag1gkKmwZDezbs49Uuo
1amvYxPoediDdeS0Zx59Yut5qu/Y4IqD2S20w9cDpvhPszxnCCgNDU5j0QANHJUWRjVlLb0DX08K
xLC4EMhLUsJDoQWK0NB6lKBDowpQnz0dVDIx2oL9oOupK+LFvBzCLliKJUl6ImwIejy21yOP+ulo
VvIfE6GiUcwGc4Fp452A4asaE/GyHzfsx2nv9d7pLuBC3pn1G+ejGR2jk5rIG3nwRnu3Se7p+TXQ
CrMmu+DgMrry/dAJcdwh1eQHfIns1Qiy7MiAid4JMfLqlx3iq1c8xa62ncWAxajKb0R5cM8aaY5u
FvbZdRAwC+w/3D4gcDlfquKGJul1Hs0SNFASpkyysOCjTquHwCKDXV3gQ/gdxNrFmTxaaNeNeKbi
w/K1DvPz3EHulp1dGy9wiqRfrhw5+nFgLIimtkC6mJY5VmdDgfc+jPvS9fNghQo2muVMCSEwD4lU
6RlJ1waeBsa6nSaDvFHx3tzVIzgn5g7j/7JBH+rqknu4NFc7Bs/+rhTVCd+dYdn6uTRK2tbEJsgi
YcUa/ffcD9tVhcMHIfs4vmsMh/S0hOBBLOgZ8S6dzVqsI2CKxsvVItKot+v7pmVEL7kjIWwYxV4s
Rb8QNxw6PITpCdOAhFaCzg629Xl0lAkdp6MG3d6nJKMSY29OMI7LzG8tJvay+utoosy0bTSpgSdm
3WcrEUfcbsMX24ZwrpOFcAvJx2M+7uEBoKoAWDoOy3yiUkN82zA54eK7BVeYk19r9qQrr4Pvn4vB
5tFhznk67yziYgBOLsjpfQZZSbmGaaJ7PlM50RZXUipaUkp+SkNuUkJICrWII74d+Fp6FkHZ6cgv
UVVLnrLtbu/5BPocBSCO1Dai2+aNnG+u7X9fBDxvsnnG6PLlpUj6MtGg3i+hlDUFbMD+snlJjLJY
cHRMCA0XKN97d9TWs+cHttPsXQa65kiypT1bhpkK0HLvlAMQujs+OUJ7OiQvstDTIrcr1lf6oofC
74rU4lB7ciayvZPcdUkBQTa/inJiWW5mgM2nSoP+WxTwRdSsxsXQ/d2pELNhEVzvjGJepXCFGuf5
EU0eS10kOJAbt+trULv21gJXKwW+OJCP23nzf/CB3XE2c5ahjFfakcx2baQTWWa0f6+Vz8TxaAfM
zvyjWTPzQExAh9gs9N6g7PVbyCvxkj5C1ew4CsfYMce65VItyPaBF+uYlnCyBdy3wN2rnNeLz0+T
ZLLe8dmz6gp2RW+ukBwBboZw9bgFF7GRpYU8QJ20wckaH8j1lAz3XKr+Zb8qNi/RkoNvpgWdGxBJ
9LB33omvbyEkiijqXaHflI8S/G0wIjuz79YcwQdDr7cWM9IY8vPlRyqPYZ+5/np9hzCkhDuvO2Q6
4hfaN6VU79wWWiJHQ2YZtqNmMeHwKI3/N4pJo1lhJqxadniASI+ic+xZhpws51TPzjeQ5kODOh/n
bszBghcIF5j2aQSMgtvwOVvBZBJhdHyK5w8xltJFt0gL7+mXbvWFcYgreUsGb5baEyML1ybfdoWk
HSOSyXUyN11AuMWOLKDbqF+TVE2aJCBcBmhP3LlCU/F5YR1eyRv+gxgbHIgjWjzKGv2i8fxaGFvl
rrdA8p7sU0VJ7fjcZ0rnt2dNoM68I9cKNDaXcS+WtVCVQ9XO6n9qlD3xxej9vAxRBkbYT0gGhb6O
GD+fiNxkQ6Dl9g4DsCDRmm6y+kqJLOvjVVmRtMi8c0GRZFkOSlZYM/P8zhLx1jNWtPtwiRWN+wDT
wd/5SDh0jCeoxUOdmML8U++wG+mRbzEUvZIctCGve9x7hxCfw4ZbIY+qWLeE2TT9GwMqKtWRiAbE
64jDpcwBXiTt7nMC/djqp7onp/NCilr3+Kf1kMg0cd+df65vyefL9Z2+wO7hsw8X8Ixn6CoGnKhq
LO8/Ot5v1/dbMxwhQe7I2XAHehCw5zkSpttWePnSigRxIpjGQ9uQuKcCI5WcA4rYrdAH2AFd+uGq
VzXn9seOD726Y6vYuyTX0uA9q8CqTw7dhyHakiXDOJqGDnQN7eUwRggg2fzEtNUmK3CS+sErs03d
qnzG1f9Z6hHvSkA1kp2NAmSAGdcasmYRAQN8agDZ0n/npNEXQcLRktvcTUBvdgHjMUZKDkzrNQJO
Ttk/SmwfO53ksMdxt6Qln0io86jWCEPv6cVPb4lujeuOnWSADslf5wKJKxOHdDo4dXHFUa/E3Y1k
l4YvY2DlzX9VS/kpVkE7xVnlHYUaGgH2q2Mf+cSCIOef6cv2sKioLMC9C4CChf2vSaLePXn/cDzA
9klaiq/I2KRBXmC3tQ05OMMXW4UEmle7LJmfMNExww+B8cE8hi4JPQ+DMrNqFaWBwJAGFjnO+Myx
9h67pKEokxvqEN06DRxLvAFiKz5rR70Aq2JOkuDB1zh70Sqa6y4Cd9Dxj78436ubdhwax/RcTZIc
4GZHhEmOt3UM+weG5UtMSUxy+Lw1S/ihB4E1IcwvIWygUW0xfDXbJc+szuZfNrW2+tZkGB0U1eGB
k7E1EVJJZwjUlhEDaN6sd7k4hBD3bBbMc+iJ+7CsZ+3XW7MG86xOxGugcjWxOXMlqmEw6Uov5BGD
9ybUGNkldce64Y19nv5dn/tzJPKbyt1UT7xQoS0XgRq3LZUhdohls6GJwB9eqYLFLubdO9dXSwfQ
IFKa5p6/xelLTcyrVQlcYg8/Vd3Wuan6JgyaNUpzIlY04vXJy9ZzHcB6ydejX8X/BF4F+3a/GUK6
mMZII5IdSy4f3tUqHmYGOQN0oiFNgL9dfpZckeNWvlpEo6U7ksNznKtQbN/PCqqfV0Q4qEIk9aBP
EmWZdC++/UG1BgJVcTEx2HpQ8iF5/V2KEZ0z2LjCXRO0LCmsY/p/2xsrmHpylTa8V8CPCiXm5JXb
kJ1azzMYRrFCw2U43e99GHBNc8DvZJFNbZdSlWQJC2zhgG47kUFlf0sF9rxvHMrtFf8DYjMojUnn
aX10iTC9JzCOrGs3gGjMOAGcHrCUbw9KQMdTNpSlvD7zzdhkC3kU6vfZLRh4wrRbf6t9Iq4EZlYj
yhfjip4gkI2PV1A/2Lam/IilTY3FPmUsGDiiSOgqKh8u+RXjMGKqjb3HVXyk+pEXU/1Fsw+fooia
9/jG5YPatfWEG7cq+5UGqrCdJurNVaoTVcFszN/HNcmp+UDl4AX0pX71015GBV01gPTH7anNehcn
R5RDSM4dVNh9plsGT1QlaueWM2GOPDX0vMJGOneB7Xks8AxlnYVlMy/deXrVl9dkW8Fx7NGiu5wS
xhUsOjRXCMdDxmXuhxQrRreJF1C4ztqaRHU5rx0A9bEs4tVLu+et2tN/LB4/vUKxEhmsLHZL61D8
+dVv2eWF03FjUnOPSi/MKoYBdQzxmgBCX52wuaZ2PtEm6JofG3GEFnM7ZY2g5U2NEcbuHpH+9h4n
z5fs31l+hllexJFrVQD/B9Sjc2Ol8WpghbYvNNar1SdALOv6EwdAxPAC5snTC9Ko/hfaIdjxsPH/
0AhXmK98Kxe5JHpj1giN2ZLGBr08kLjMUY5wr1qWNtgv+a13RgS/NeFe+8AIO6OZE9J+8wBr9agS
ZwIfZ0njsMi1jvWqVc0l95M+lI9TgG8jdNY+XuCYh1vmwVhnlPFHZm8tQvQzkTBjN8Ff34+F689e
GN/z3FoI0EKR/yHlL/Tf3KUuldM5cm1T9V4U/Q0SvLKP0EK4GBjfEpsrpfIPas1CJe/ir5p/4lJh
vzGb/vwLTbtFweQ7YRFlC5dfi3Ol/yzcXrtG/saCQgoZH+vrG+19IESN3iVniQHE2rdXZgYCFvM0
eYLL0qUVcOtC1EURce7YK8vPXBPj6J4QUnVrx6BQLCOwnBya8c4AN5b8B1OdN0xS6M+WvdAYHvmC
HJTxjvxvnDAtU8nKmd8KE/p7HxMWodNypn8JdZhFlDuLYeSUPrYY2CucUfnBp8ZCWU5fqZ7osms5
wNbOerz9Vx1IMcaexV2UIAF668MbWB3u3k2CoF77DlsJS+tnlzUyZs7rgIhNpTFX3sVOKVoVgEqO
GpGaPiTTqGDP4vS989nSoB0r4Z+Glufe/f+7Rp+ESOHWqRwVs8Oga5IscPWDJA6KG2Eha0K3xuri
8Hr6B+tfudN03Z/uUU9/sSyDR2YBKaJgEK3tXw2ieuekPFjSi7mCFVoVGXAAmLWTlLH1trZs6k7D
+Q+KZwmr9B13Y+Qte6SMaL/ozXOLEUcFwb9JVNcZ0XRYc9lAsz4bZquel3P3TDwIk+GrHQM0dm1N
FP6SWBlIyT36o0Bc4rwvnUzTP8wai7U+JwI/VOEs5s0rFXs3xIrZHHIgrEavlmxtMHMgAp+l0quK
6NPzzzMt9RD4OmPMluTZwv3YDW6tFcE8F2zFxr5rbokBbkoRtUERWuoyNeMg0k28enl9A0mEmL/v
JZEB1gUxAzIkCyFFMZf8kFMLq8katCDTfNYkdeOsF1JciGsLCPSgHU4vYTrlxdYcG8oCpETjFDSM
KuQNWrNoohn0g4RGfjb9p78FZOmLV4UtGFoXXfW5B8XXMZ6DBbqi9tj3TG1OYcBUuMxS6soLkvZh
YrSS9uhR7liI/OiNPHwc+hyRwQGLyoUfbg8lTgRv5pTnOXH6oqN3CEiL+bVFXlgpJUhD/uE6Ozux
/q515ho/bwvB49vdJ+S3xn22jSq7NUFzxeYAM4acOfZYuAh0Ti+Qk31qCj77Mh5BSzMGy7rEVnWa
zN6f6xeDwYQ3w/doYNd8IkqNiHAaRfJwFUKVdPoMXPkqYFi/+6thfnCIcODgy+3YZG8L+EDj5G0e
E/4mCde+iROkVAe3JbV0Ceip02RqvXJfkYRibYdlIzEGHO7KFHuP/BBm/PLzpFrCO3JlQ7Ixce7l
bpCG7ZjMzz3Pvxa6QUbL25HH3Wi/S046quhcgmMxhLM0AJZJwNBDDlVjXeiScO30uHfO27g+lH6q
N7+KnCgxi42R1s7bBkhLCWNqTYZrHNDsw7wqeSfAhTkG8su70qic8LryaOLPnkWZPnKoaEbvvu/u
C2ETK1KeLFPaA3ybK40t58M/pHpQalKAejaPM+Mb/YcxqM/FWcX9DXuYiA7MN2aNr2yp3sEot/RF
epxz9PQH07+21EM1QLsqVllwh660K4O+JI7wHuJ8ScsYYVLsIf3owkNwg/1czpZuzg3KrlB3ehJ9
MfjANdBosbR8pT7YAI+bPUhR0g0eTMcZc/kFuidupmt6VXE+MaRSAUDzFeOlSpwjx6/p0vgY8m3D
CJ1Lb67IWlC3XAA2n3rljvzZw8k+bATb91fFOJfsYfs9aQD/fHoHOsr14PupbUjpUprfJhpaghzj
0ndoB2dxwQURFhSOrW8DxObPUiqAmLly2fwJY7h43RB5aYBN8ZSHS2KBuROlmAKZSgb/aspURCP8
k0yJ7v7ng+ktb/w1w7IfueHZanOuKU61wSuJ/kS/WP0dWEREAke6iD63TEHp/ngaeG/PU1adOFuq
21zd9nEzS69/AlSN4YwLxQCzmwRzxLVnjysxyVkW3LPcSn4rRc29IHJ+j6GvNZeB68xtlIw+yjPw
y0AClzIer+kdXZmC68WZ7mRkGkq4mnYRjEkaqpZ0C7IRAKLBcoeqpM98IZoMiFNJOT/JEePb8fSl
2iDFyfANvvrV+lJzFR0dcC8u5ESC1Y4Dao6S5nYP+sgQYlMzgueou4HZ/YwVCg/BAMcNMpAMEMa6
YZjUkru3m965N+OwnEHx01SZst+J/tFMkciqiPJExO8GR50VfWxwuu0uL5GkS0ieSfK9hxjX0SLz
hfSzTKr/nHrYJLpLmJcc3A8C4O1rhqEbJW1Ln3m6ovXOcTWOEA4b1E1aAUVVgngORiYsx8abG7tp
HitHaTIHO5PkxApZ4DfVBlRAvhtS/kcjNATT16bXc+kvG3JbTRhVsQLu6foIJxMWkKuVdUJ02e/D
87icm+Bpo+f6qB5sM4PK7USmshJsCYcRp1i7HLEKY/R031smu1GKPPMkri7rdNSTwzReg+ntxnAF
UQytOmJlEk08OoIrkmB7pvU5Da+bZqnF4Eyz89ZnF/w3UOn//1GwN3RSywJCnhaJDU+q3XnQ+4yD
pp+k9A4i0yfu21bcd+OchaAN+68XvjqMsEydrP7TxKDg3bcIKC+C/kUp8xHcY90JVn9U4iMlHaHa
1bCU5BkKf6X/SvA7IJU9UsEP5gZVBRTQnKWpjBtRMVpdoR0Bvq9DZaw3NcPYGqvk73vkcHYXvHxk
BRY3mE5lkdYqsJVGYsRBuJOHKEGgRmJ5pAe8hE0HVHEsBs2qJuj9cJ/XdMJMzNgMHeXs2RaSi25F
WwbYMqwtmCf5gIW00f6fKS+7IZiUWXm+eIIWklWis7qWi0OCkNA0eXgBJs0BrcN6jLUKqjTe/y+0
eR/T3CcpngKl0mhnGuEej/HeRAazqRC8hJMhKPqYgVB2IKCWjEJaWHHNUhYiDtNXwl1awE7ve2fE
ZQczSn0zonI/lzPvEUrUtm34T2alQZpyJYC5GSf7Z2t0prOEoE7snlydygkmcKNdtrcEYfpuYTJE
T9flj9B5V4uWHNVGoWgyT3e9J2H0mqiBD5mWxvk+wUVnGZHFwo3L9iV8yJn0WtwSnc7JYStIvTNp
v2ZuP/6fe63AtUfOMJa7XeTpMxtsqR9bO4LU320XEzgrR3i7r3BXsbYoKwcCCa3Io3fX5wu0r9BB
dzFMQ0sxAumfoO5BFMq9M+uSy/zbgHV9ZgoryX8cgGL7nyhC07aXl7pNdCIR1LiaPuiryWcx5QPJ
DqqrKe1AuB6XJZTLo3sARbCukZZoE5T6qwj7LmufmOld3bKteLuji4jVpBQgj5z2xg0aAyBDo5I3
gk7fpW7/mKpNMuhsh0e/T8NFQG+8HkT92w+6qkbMXFP2D3iwASIXJxWNrg5c6awXcB1pcvT/Wk3y
mlQj0cBke2o0eyFuyfRFBTGxTr+OmwxDX3KoiuFfpl6F7tRL2V7c8dhMZLdke0Rd2PBDF1KyR5T/
gxbAWOWfER+JNGIQ1Ygzwq2y3VYdWzQCIP/JH3cLWZbYId+jsP+3om+tZaHYWgE8fM4iL2u3cLDd
FgNGY04W+rVNBtSFLqzd4KiYMc5TV3L3wJPy9jWwhhldxu0m9sfezYSZgYV38kQueeKqwxjVQDvj
ssM19nh5JrdOB2jX4hMFZ2KH3pJwm4T151k1XgQTeKz8IYpBIgCZkTYdMezdQoIhlQzjdBzddy6w
7DNNFw/OfWOL0xCew03POwgj7vuPySuro7GjQfyN0OlE0ow6bp9ZN1XAcVgYkuwT6DGHZfLLMusn
3cX1w3Hj9vATeo8nptgiXcOEy4itZwycufR/I0uMsfsjJtcp+Z2A0Psy+QWsyepbHfW7HLJoKblf
57RTIokeypBuKbplMgqUq0aaIkWb0pEQ/EcoOz/wBqtaRVM+dhU0SIQ/10Uz8F/5tI25FcsQ7m41
nO1tHoNWsN9/GdOGsnFhchaknIgfG1/I7CQNldapTvGAZ7ow9ZMwwWNA48biDqpN+pNkiToTwvvU
4Aowx/Bz3pzFi+gORDE2BSfWmUqH1xD94txyCl5eVg1UDe/TpPmN6akN31vGP5HH1v79A3GKzePl
Wp8L0W49OdMB0WtF1R+z7/GTc7SR0SYomWMFa/kVvEabWQCNZIK07iLDLR5tyCTpBoGfCCU28qAt
SbvBs636iS4bowNnIIDfXN/No531WLWcD9Re1OKVmD+nLd9AQ4GJiBmGEbxWioGvMpxbELLD5dH0
Ifkzmb2vEBNpXqcNjlt4WzdeeKOEYdqmV5RuPusKN3akXbG7NckBFLDoLDXCcJWwPiCnciJB2vfP
8HIR/FE9abRoz+5bPYKjfL/GLh9r+ixXUoyP+Ij+ffYlmUtgxlAOPJq6iPI6Zv/zSUbVQDrgiieW
o+iSfORdSwjbR3yaaMrmTlUaVgVrz92NfRFvUDm/ailCNwgsbOlx2Pq1GP5h6GIoebyVIl4ntmWF
GAKXQzULA4x5nrNkJYRsFFVdZIwSDM37OGFuTC4wzEoP6pFcBkPSve+hhqQDQKPD8e7WUcTKjV5/
ahada19j94VIilIOViq+SDcyW6uBLumkfWh8mA2sPYci1OXfFk6xl3DAREx9w06QmrDGKKKeZn4+
0DcCHjz8l0P/jtntIaIpySMx9nom4Ha7Me5QW9+kTGrWcVzFAS46ELQNyiIBHUD8SHcG0QLr2DBG
zMVVDo8lyxA1rxhHi9OQPUD5V1Od0sCwyudvsnQfh4u5AKmdF20Z0iBjfK+hoZz/sPSKDckPEREj
tXk3TTNrP8pCfpJ+Cog5z3T/XpUN9B2bwVk1xgewW4RHZ7ICteSwMQ2iNtKbuzo4VXV2JDeTTmgT
hcucnFa3KLdxgEmiT2tp1/2EirVg0NJg5FMbo147WnxvVvaArIIBvyuRhdOd+4VqXnMostxBvmvB
BOfNa6Ue9wc4wdEOnUnIEQhMzyx8B6QQU37glKcvVS/PmKKm8OF+79wwTQW8w3IDLxp/mQA5jd/h
h1bNCiDOkaG9SOO7GOHXYEML4uLVqgGSsqeF7V42sO0NTD3Lnrzy6u8gv4tON6UUEjXDjxUzGB1c
p0Xmt/QsE/MdTHyGdK0YP74L8pBVvE+pUk0kmeHGIKNCdrQxxZFI8YN7ROqKiv3DGSAmfi1RsE/o
EE0afq8kCWIpLvEwdqu2Lq3he9wppgvDgAYcTSlHjNEix8yG0PQDtKCZ8qzb1+7dAx3vM+sYVDt4
hJdivF1P1Qo15/NtYl+rb0AMYVhzH17ajSIqsNeFB4RL4nkRSJDudrLrLgZd/7GtPO+Hu+pWwq6n
RzdNN/4hyfRUyRLu+z56877a+jBk8wzh9wfqrQS+AJmWth+X6LqPctm0MqQv5OlTctEiKl7QQrDw
CLzwv2ZDNyr0pxIBOzn5um6LIS/VNKSIdEfnrrFvYOsmGA6Uf4wl5MzVTS4D+BTLxJT3DELgcUt0
e7r6xu1kTu8T43J7pGptV8wXyN0aQsnw5Is90lpRxanG9fXZLIuwMcD9sTrAE79w5VkNufPqCUSV
bimRlYk51eFe7mN9YFzA64QtTHX9Jd4V6A+s8NUGoq46L4M5Po0Ws25huNP9y7zsasCeLQaZR8+Z
Fl00uPvA1iR3fCfXANw58Zwf7drcqSGFHJSiH2LeF1pSROxKvPDSrFPeDZuv0ie2WeMLkLgjACS2
bh8zRR8fMeb0W3Ud431m7/Uk3yMazUyv3v37YvWH16uj01iymX49bBamh3xO5Gw0iJg9y6PP6GUa
VjM94PUs+5dp5K/qUqSVy6nUC1U+p/1nnmnD97aTSCd1DdQl9mw6ddSOUrYEfXtez2dx+FERkwXv
GrQaLh2my36cTU/W80a2bKiSCQugSLFUBhMqNJ0BiKWyF6B4vmQptvT9/nzcAWS4/iNDTz5FgtIZ
5ajOdb5rkcdUOgzVefMbJlLDEcMmab8lO6zaC2eFcsCwWl4MDeU/Tz6lhrf55KZ4ON0SdvXrN3x8
05k5hQxjT2az87x4NYOs3nu+3CfMsxZjqef1guC374R5FFecYB6adNPsck0wx2zF1vZCrG8FMeEz
6NYWF+FNBXvb9NIELrjYW/MO0liwA1tU88HTUHF8L3U1aacrjIsZRAOnCHEV+NykQhVQ2cszsKzC
CmxIO0plftRIoF0xKiffkIN2ScG4VwKOi9fiGlPTqMaBChNVG6FpZmGqWCVWsjTnxE/NkfP+bppS
JQTxUoCt5nzKpCKEL6YfgKLBC7Za2WEFXfgRbMKoBL3QEWyZhn9iObFbl8hIFHrHBjgBrcxvCz7i
Opb52VQnogW1sSxvyba9rhDlrpAmkcuX6f5A76+Vx5appZZBzlRWqdgBBTUSwRraRnriZCtf1sYB
NILkoOtgWCXzcC5Staf0CMGyS0HhBXUhJuxWm4mNoEclqLoOpLwyvMOP/wEMGbi2DmDZYUmIjTBj
AHJPSlY1pqcHmS6wd/46Akx7u+aqQoTCxtAT0Jjd12jjkx0G8Z1grr61fdKGsVSWup56mRuZFMCu
ZvzjJpTL6Z22BCyWhM3HdkkTDgNC73akPtOFpS9fav8GXve8InaraKwsdrM/3rULZlU73TmqbNtZ
vE5CP5KZz1xPNxd1nhd3mKcQSahNBC3wkAKXYco9+katn/wd9zp3aylw7qB6RIqDhMlZRw7nKTRu
IhmlkX6valXtDbwHY2SvPYc3YVqpzno0G3jNxge/40Ti/GmFWv6GMgfBgSRl4eKvLWBB+P7cOHKu
pOpgGg+BxnCCh2lUBNng59Rx7UUiTk81+Hy33gJhvxrmCz+ICiYik+sO6MsGkwoGn2raQu5cJpKV
tCGgx0BweiEFrJ3hB6iJHiSRtI33373RSSpDIHvviSfcoolvXvdD9BuSQ1m2Zxm5Dw37zDbdPK+e
c9modr/7kL8Yj0bJ2A99xQNpkyPlLKsLV1sJQhg94gegZlmG28BFWPJP5KoWq802uqUvynOvoy6H
FxOYzDteDw8UpxJF/hCJ0N7OtD2GKh5+iXerhRbaOZ3HGw4i6rS+MC/3T6ddtn/gS04Ii0gEyp0j
tXkO3o7qNguJcCt1zu5zz72Ex7PBrti0A1drnqziXJqrAHbcGcqRifPiDTZvrOIixP1dh6+AMPHG
ybWdh6LVhNun9gquOf/ZVlW7+6jnckl20558vlGWKVa/vzwD2f/VTXpgViWshL86OQpcBh2rp4Ip
l0/nLZa4X4lNGDE2T2Qmxf5WdzVBMbH85/GhMdwkOI/aHvIJlnxSZwpxb8BoGa8RIZedga3681cV
q5t7q5XCWtnkxwxSfXIiheWLK9ZOh2h6L3og/efU9sRaNU1B8yjeVbKnBIpKJXeH2FQIQP9sXW7U
ilIv7LTfDZZVft3oV+bx0TznCQJxwkcUq55NX0K79MTBpMtDl8w/ZKlmfdfFHQpea6SLGJ/Bif7Z
LX6OEhUEA7uGjHeUIfCtqgvs5EraIgeZtlid7KNaWvdK4lZ61KPGV3VquYaLBE4bxslsKICEYexN
7uCck8YWKzKwmdHrAwKWdNppof5dMjtxbY5RZvsqTzgTxn+re1LG+tPy6s2208XaaCO1f9IeEBwI
iC/zuZaLB9odZ2WnSRMebujpv/XE7yP+xb1r69wbKL+1IiLtySymrrOsc/Zk486SlJN3v6/vcFIY
dhPoJrd5XJxRbLLi3f7pFhgDDugyyyhYITV4d/M+kKeIrURcctG75kzUib1649qtNXQYs0ZxGUwG
KRQUscAzcldFmmTvzvzhQgIZ3h0YKKGHflxl09adQC0ZGjQ84k2OsVV11LMTeeIXgwsG2bAEq7Hy
izcFfgPAMwehqrsZD4GS76jwybF8u/uE1m+ow2CMs472dO01VLdn1SYESVi2EuNTK3q5KhnqetJy
TZUVKELkmAbjE9rlhQtw/7MW+1sfimMgO+QSZLn08BXeIPVxByVQ//8AN6K1GlqjUenFHO1jbjMG
dNaTj2zU3ZaN64RVpa8mG6XoVnnhNCHLEIal1lSbfbwLFM6VGZbfjkvJIJDqNnYh/HVUyteNpAQ1
TECj+bFGknvVi0RWEtVtdHrLGNf7bjR5DdrhzAHO913JqXdCTUDIXJPlhOsCXTVQquP2VUUOB/oF
Bq67xAglMw1GmdWbAGsyZnA3Y2WXsSbBwflBgaJpA6hpBwakacVyk2dWI+Yo0wql3IVR9vg7wk7L
JCLKPEufvGS8PECwyDvM1dabT/dNUNlf5G4CitN7zM6kU3u826Aozn6wY2jNXz6GikYwn0i0Y1ao
QnGbQ3wXXOV4O+VbIIFYkUGudUsjCKlU/4d3Z33S7SMHWLKuPEM0jWrnW/34+/WQadab7fJRiYeG
a9DjMp+Kh6Lpu71Yhm/mwGk6lSs07hFcaaas41kyCCDy/+Y44gcP3gzsOpnB0gA9XGjP7QRednIl
SMpBJ72BY3+DmN/9ztVTR+Z0ihtPVIe07eYeZBKcf7PQbe9IBdPBdhSnDbVhGR9NvXveirnBtB0q
5Ge251frMyvkyqEx5J/+glNDSUg2utUCiN8GhvMqw0hcg62Wu6hdn3qUHWOUXnToYOLGO2SzZcdT
z3wiZ9sz5mQjGfBm54l7QdSumLLOmHnabSZXrvHtm0/F3YSEAu9gtkayrmCFNxHkOuUkGuDTcpbE
ijSEcTImuxaUuzi1tQGqH/y3LFIt0c2vfX/8xRv/dLC6H+Jl8a+hZhMcRvc4vH9WHjmP61VTCAlj
ELf4Z+V6VZWcytGO02FT+augS8ZBMhcbIrM/FyzJkjmTnHyLTB8w8yRDZVxFPdUT7GSc7p6ZmopZ
33INZtjFMQexylsajP85gc0jZjWheAs3rxKiLuF/kWbaCePzd4aJUBt/vRXEjgOMCUHZCysVkhSW
UAlfONwJdxdWlyBTPTZlBhV+lA2r27GKM24KVSuKgRgWcCDy+9/GabUTjrYjMTZtw1OSObsPXjqF
pWDpUaezYNuUWm4lf4EP2f5/d5j/G4H3X3hoIo/mkdGnqkYJ5biWHpxdZEIcTcY+eSuKcUM8SZyz
FqIiwFQfPsx0e2ARSC/enPXCuwV7ndAh+f4ZX1+mqfwDD9m3XtrX8e2ldze0H+x8fseu4dQNKHtm
P8xRktep9OYVqe5alyF6suSbCxTLBouKVFNjTzPemJZO/C2xK88zJC/LcOvy5z3OOlphUDsLvrFa
e8nNdpOLBkuh/mQGc3F4Qx11tN5l7Tibu50Y96YnM1XMzdZBeMqHV+MlkdQbvtusDycdOFaV33+m
PighZSn4i66PqQzuG+Pu4mODP5YlIlLRzSXnUs52jo4XdyPPkGTKu2Pchwh5OYDgS4dICdqgjKPk
TIzUv7fhWJ0cZszaNbyIO1Hkhq6CYYBZ9xoNMshECinzSlFfv7Bsj5oJD3lmCTC0F2l8jt5G6qzk
LEpnfrxO7ghJ7Jk45Ggh4offrjjmyYAK9PT9DmzunMDBlCsUslO+fPA3UBnkGjhjJuLlbvlaiVY5
pG53tG9ll9BQ/+Qiz35z6uqf5NJPifQ24HwnvQ93TI0ySZWWgGpv08/x4mMyBrV+86aWdEPCu+J1
AdQEIUO1AYPKgVkqvA9GeeHF/Rj6MOVfHHPyDThHuQ2/NCJq8qpSsNW84mtDgiUTtPWeiKdGFc7f
/Zbg5rwUhNuPLqPZ6aH5NUrp/V2mTRReLdUjJXbceVIsmnM74H3Uf8xWEVb33LGZ9rYH0zFvC2E7
eJUC0yuxJmC3xx8vkhvwgN3G6kB/F025jIHwWHVciT+ivLryof5PiRe7ThWyVrr+x7rKu/bIjYPE
ydNWb0IyCStuFSHUcftATCl085OXt7IXonkiZZp52L4p6dCAXj95+vFUj6WQGM5p9gGRBwoUrWw0
suZXmqPmE74w/CY01LGzf1K7rT24aJ6lIuw6QIQP5lsGSF2lC1sZP0rCpoW7O2O5D51TtkdT+J4v
xiBJy4/c12ukDEvNEVt7t3HACRF2X2RGCYAqPf7WX6zQ4XQu6L63V1G8OqyqXaUVanxCNmecBpb0
NNPOLirEWIpG9S4gYO2RjgVHCoHHKhHaf7V/A8YcJhf+EBaSEc+I4YidZ6vzH7Yb8Q0KfBiVfhLR
YBJiDMbdRaf17YiqDItj0oXlEoEWZmemnshSNJgtMp+Z2C7GJidfDbybW81phWw1EcOzs8McL7iz
D4GmDbwNRKo2MnRwCyRB+Nn4ioAdyeRjmLTKt60+druYQ1NUX801zsMKuaHNCElqZuOCmxImcFIJ
3lA/XTHFpEf4BXQXRWF+LpCwKyIK0m8RTCKHD+Lv72k8QCkOo7dZWA9MpbYh2xtBREcVEaadUiTC
SpUMl2rgbQw5DVVOYHEEKBXwoqSX8g1oADh+nTuhLBisVxy36OfeBP5rhMOE43yRqDI7vtVIjgq+
AbVymtV3S5b8MPPYCH2pBC36gxDGyGt0wdeoNzxxTmkvDfFKD1dH8gjYJ+MVzKotwuc8WfDiJg6V
94UnPdBoZ+jXUCB2GJl5/ksnsCcHflh8MJI9D+2gw9f5VAxhH7rP0zgOq09PsgplDhZrncruz708
gPOOyej335Eycfxmos7/110t/x2q2itsZlssmSD0D8zhkVY3kT5sDCKew3GUoJqZMlxCXaew6LGH
vQCnrQebwVNWLwKOjtiNAR9Z4Pucd2lI2/J9VdAa0Nf5yY9+SzR7pigSz0WhvWoyW7WYrZVwyJVU
QujSObWTauqbL01MvOIZcS1LC6QdoTP2OrG78BgrVHphN38w7H6ehaVe04CA96LeiVRYZ4tdK1wE
tPyYK13t6C3iMjr6DdO8eBbG8F271baa2/lUtZ/2XX2+juwngwdqE3QhGjzD9TRoofigUXr3SmQE
y2L3aKDTBc6aA0XZzB2pBBeZgdvHChmP8c0TPWyLNNGuQUCYtW7ARlfdpZAF1gG6SNln1xddLqar
cgnNUdbbK1Tg7J5a/ygiI1Q/pBr6PW+IVrGtkBr5jYcU9ebdJgpXmKWEfxiJlMQe72ZwEF9n9R85
G2kAhCa3u+J3QkEOUe1DyS8x8wxTckBOiqaudNJLKVxA1tZGtJsQqFb3mZzPIc6Dvjz3rvuvFi6S
hYkUCq4LgMjBPRHsmOrzuonr/rcVGM5qs+8oRbevFEP5OSRZh1BxRwEJl/elLaAgaca7JMrG/ZJd
Qx7kvGisNttwj32v1ewEE/SZfvxkI7D0Q/aro2Mtt+iDmjLRWHRTmJZpsSn7CLNcFPJzRZKr7tKc
he7RMBCZ9BS9WBHRDfX/YTGiiE8uJXQFKlMvSpaE1v57NnxlkdMTw78t8ZQ+QZPn8QKLWbzdYC7R
bv4Lm9Iqvmn7YKexiBo6AyaD7WwQShbTqD+dOijewOK/dL8n4YpnGIIsRrRcl4NOZv901Z42clPt
pWoVpCswr3ncdp85/MoFrvue9QbdB1zaSr4NGwPnhXVuLdXZcJSFaDbCcFy1pvmh7pf7CWq/uHku
aYdmB1VGLGzUeGs6+YAqJ5cjxrPBi+2U9slsSQqkV6yXxYDMIgB48Nuz+/aJtH8DIj40KHKbJwoW
h+KIBicupN/4MaZLogwD3Sajjz244AIIWUdhMWLQX8ubAmwV6fRy8bJD3nTrc61UYBQvjJd9zqBQ
YiJsg5VBMKQatO7rOZGzn479PhmQPxVghJ1nqeRr24NHKBOao1MrTmVA5tR7Y+zNIdSpygKEGWj/
2alY5RwaxDI/7SaoASEVaNNJIVw/QI1xBXek6lkPy55WEdh7gAOwgfuZ7D+lUQ2kVOeocbQWUcDs
TgSdhIXabqvXrtGrpxIEql/5/qFGcd7Ib+wXqbl7xSXJuANA/jiIx/+E/yaeLZJxD+ar8pJk5ZHz
oV16rTOUlfFTFNIxc4MnnQkep6v3e2KJ5reNFrzuhInrJ23GxqxuhD6S4ARRtkIwx4f8uCFZknR9
AQ3Rc34ejUtcUPj1rY0I5DK9twxlzxcdsUhM0RuKh+R0pw1SYvd3HQZ0/RJ+zKQ9OH4v1DGF0Pms
AtuTwMX0s7fBrA9mL65gRgJ29J/eCaL0i+uemhJUZHPfpc2VkXibe8eUUFDpvo+JzTXd9z+TCoKX
AMhD7ZaEju6HX77npGqKw7oRll4I0ttZS9GeNBZ2ZdsILkiKghu1nBLMYjA9b6k6HdexJhZkKoqy
i6U2DZ4dcQOCOAQRcbZ4j+aZ5ytmrKGcYG12RuDaID4HlFZUkgG8Fxrlz03b9SFFbvtjZMY8Y5Gb
EDAJiwhWVXbAiarH6nYuzfzcdCq+KDVAWelbQFMVJym29qYuN52xnTSCDl3bph8WErqLD+eo3f1F
2wlqJyDCh0XIfLI3ZVnE/yp9fmh9ryaMDCxtk2jCePl9wd+V953V0Bc24JBBtQzJEYejuYoUvxp8
k/2MDh8JJ00FxNESYBo22l70xqfS6bguM4DmA938MKvoYSdnKHfoFkL4Xa/edxDeyhKIZ1G50K7C
UZBI3PpAwAILPoMVkEE9ALYcXhM/zxT11+wNdPL81ZsDKbejOe2JYi+VDbs40NkpGotax2nI21ur
o4Rugto9B5VCAxBtfJSsjU9T6Y8tTkCW+yYmoXLtRlg1bTSgXkZrqzDjr8OgSHYYeBahiaiXmJ3+
VFLBj0ON83I9HP2zz0CWsZu3YZoXRlb9SgxGxYn7/BrrVduqKqs+O4k7LHeT/uUvEQlhTZij4FhN
7E0XHebpmEpr7zkdpzm0pm+6GpNwuhqJY+Vo/ahe/zjZKzjiFo60UlYInOfd66UMyn1UmYc/Vsb7
4StwFoRADk4smvwf8yDEBTahv6p83xOj7BcP9TWwfAt1uc3LPsTv2KubzRODQLovSx0Gz52Gmf+f
lmNAbIFbZwpeobrJGAJOLYj/vY3zagZ6Ti30PG0MykLbRfrl7qbu/P98FdBAuHMnEddzh9MHttx+
v2Z3o1iOYkAXQ2whvIO6VUzILJvpIQekr/d3sxO9CImzpp+EtMMA1zl1BrTzcct0Jd6bwrmoiKz9
nXvdvPxVbhRSOzN1F6ZubMoIovTdwB5xD16+5CKOM6XCj+Ts+7GH0+8mAdeSqPeoVuUpIpKTue2K
muIM+FVXIsmnvDKY/n8ttPK9SEv86LAnBbgjOdJaqkkuoRvJqVKAO7AWVnyVKDcP5o4RhAYIg0Y1
ej7SxLwYfiXZxWiepZjL3JHiilHee47Ll3hAf/1eHgYRBLAz9vhJN74E1X/2KDBO6MJsV9qBlxr1
2GWepbC2TI4a1dT5oIuoY7LwQS6l9+I5uuNtClBtqBqou7QmU6h7sTQsL+gp5flIx6bdWW2jZfJa
ofdjUJgLPnq/mTPCiAiFr1QI+39zrZLjp7PiI/jeoJQB+WPVxgyDKnrqcKF/ijKAr0+dYIZRZ0fR
kFKc7rgEuWtrmKdWMY7GINzSdCsEQhBj4Y+v8a7o6FjmCH2erBQVDrOgvkoJIZ27vKnTKTARlSXH
3jEQnTWHqHUidI0UvugNBpqw13YZNUMnhPbiG3ghWCiBRYNx+fw1hVrvFIkxgUOtUZgBbj/gFOEN
3jRk+HgtJejonzLo1hx2Wub/fPWMqyfQi87Bs2ec7HteRvU2GCpy7Eihjne/Z3nimFihhyG0/6pd
1PR1wXmEdfLpAiF7eCrbTwgKGuVBmlrm33s458/wCIpA1ExZW3G6vQ/pgnFpkMKyf14oUD5o1EiV
DEfnz2aefXkpv3xIPZhlTY6voGvtG0AO64KaBDiHNdXoeV1M9r/rzrUqu5rfgUeW5hDDiG2D0VMV
m+h4jratl9lilV5Rn9IjG4O2QF8og5CJqahDCrmEdS7o1lR+hu3QQpFsdFUYTrq0uJOMK/AgD6sA
i+vxy5MIAglYquJv2+SSkIIi1YHNabqgv8sG1q0O6y+Opr6kOXvMzj92zVt1eqrmOz9aaxFHT151
GIbBzaKZvDXCfryxoGtYKwrcQclTxzPUq+WNrqYbaNGNWGMKiA9EWsB/LYdh1oTPf/wot661oYIS
8jQnsFAJGhWtBZHggrdFLJReZYkKPjeFwVQkxCC/okMFfr6enw62/hd307aNLS1OsLEKrGIfwfrU
7Y6b40b6uUA8iIjWE5f29X2jMFcXELViH0jkXhCLivHY0P9ydw1Q2+uhdbYxAIzD2NUoIzzwYoNO
tqnmiN6Tk4mfWwkrYprog8i/vknRr5Opi6USXlYl3Qu1yki64Z//MMoubu3Z0KvZCYaDtaSmXZPc
4CujUV7eABsS80e8TsYr0O+e9PEdo/Zj519BaozUZDotbRRJrOXF9N8AzzqPg9lmlA/AvhXhtuHZ
ZLNYUgBCEoItcG0EAJWAR+JO1rjMmtGfMVk6qL1+xtnX3nSCCv7vB2QRgR1+TtmwLJgeiXAwfnSu
xu6XhkZB7eY/IAmIHyNWzIGgT8iFqHeEhCM/hFx+H/rduzLaxGZK1NVBeY8cizwqm1lu6WYSY9yP
TW5zDKUpX4VQa6cNVQ/bJqR+ciACdRSEZO3NkBQ+PD/GQTfbntLE4Lfk70pC8nwmDkJiu69eHFKB
GyozadW5z9HNN9mxvZCihf3z9Sm0m9XyqbhbjFSGYLiErhRj5sSseusq0ZcJEMZRYdzWhyaugD0H
h/ve2hnbVRJHfPFHjcLLaDDm8+KOJf0UmvnwkQNbAyyKPUNDdc/IIoxhbwRs5S0rkxf+EOGoMFQR
cqJUK0ai8MvyFEFY1pg90up+7ftd8sZxQBYybN7gNzG8PgkuQwGfPFtCoY5tYiYKHWlYrWc+EecP
HolOvLDlwu2gZ5YmpG+/60d+Dac+JyLD4A0r4UvjcD1itTJ48Enu5SQHCOia99ww8WFRgPP8xfNk
anyUL9mLy9++mWg6MxB5kpumKJ/8IvoxZd5/1HSOMA7CiFfUZSUBUPleYLXdkJ6vT1jfSFpxf+ja
hoULit4xbKDMQN8ADVGxP5Xa3MTDONtUiYuIHubQ3PPIzSOniG/wCsSXJZfuMGMq5dfHRfYHfyh9
Jyr3eYioI6hmrX3MFsOpX7pzN0zPw5Z82K3mvBAJOM+YZNGUY+FT/jr9CF0YtltiDy/a3tF5RDI0
BlcoVJC7+xIrK1wpllPCP+2wR/wbbqDcIUHe4VM1Oi45Zwchx6P2eUGvrW/2wjX/d5R/Wh0bifLR
qcWkJWXQYaEVdmzo982bzpDgc5RZaJ+7xFzw+ZtWwlzPn/mlwkc5loIOYd97msdS+EypXmuwz1/9
UD944CUc7C3Z7O3nVa+fQa1ak7PhVZ5vC7MpPUkt4sDFaLFRb2JklOMlq/+sQeYLn89ptTL6J7M0
mZXOTJbdkAINhdNE+3nK8TgCYI6rEPCxxtF2SYXh9+npjKhqjOHu5SZyGf3I0JnQtBvbbNzPolN0
yfnFWn9+pGk+WrSemo0rQ8q2kaoE3+WqxYMr4l+BNJh0oiq19mGPmIfQmJEd9AvzIhTpD7K78CpG
kWlxHqa31IPj82lWtdMHAg8DAXeZenT7s5j1qWBKtRAKc8Z+3rHjlx0KgDv0Rg9RRiY7UAqF26cz
cal4gHI5+iZLr5zgLnbRxfF3aKWo6BmylWjIAM936kM3tU7wOSdGYrJt4TrBH5Ow/kDDu//BInu+
2+dBA2Wtmdgdi3jjZQi6tA+fSxeT9qV4DipdV49r992jO+Lak4LQkzM/9M/RVp/N4A/EA7wbtToU
9u8WV7O19rSq1f4vNfSZiWexaOjwQo+mBvCF5MRSX7IpF6OhzyPqZXboySr726mxGBaKdxr//E+F
zZNx3HsevtBR3O7qVXngah+ZXejYK9PstAG1TdXqYs/b5T+eQRu/b0bHgrbbQagu3ElYhTY0evVn
eRXQEd8JQdwcWxr3h42OxA7TGDOxj9o8D++lJq4BbhLsYpUEMCcqDQqSA3hPMDjsd7ib9igPP30W
czksRTSB40bdNKxOJfH96KXpPwc/X67HFNt43Ew5OpG3DKMemcmo8nMrW8vIA/VDQG7rZIIVMDrI
rnBFmTkPOqyARwX/Q0w7LGdsebetC6xsPg0J14kqFCl+ok1rocgXD46bgDCYVGhthwgJrRaJcipV
witqkwyddItIw6CAjRKFZ9pIk6oXxTqMNOFyKtGmOj0dTRmYTNPR2bnUUC3lLURmDnHFNk5PioI/
m4sfQRvwjQ4n+xOxFs3jSHDnJSjjTVzRPFvehpIGU5IaV+ivjn//l7+TI5MrB9Od3bASqd5zsFAk
Lvk7EgeTxKKYIV6A6nqROFo6yK3zGIwvXeYYMJEklG0IEYQAHFWFIwImSr89PrLQkkE05Xf5U7aw
vHYU+rkUBYonmOGxgzIoXtL0IlZ/vcHQGDJ6XSc8FO0T8G/1xNCRvLl/6fK6MCybRsP7ZD/iuRGS
IOj1fZcPE2up8LNxjrq6HyJaFUDqqcUWZhGBOUPzn+QaaG3vgpauE+5Z1oFrLGlHxJQuLu0xq+a+
q5wHH7i9vpNGQa+hq/WCOHKNUNB02Tqh4UO9WaRNW9pYwIX0UpwG8vPUx4Z8M+GsOiYDWi2qzzMU
4jsdN3iETOtSsD2CxL3snzG65Zew2BruDI+qwgOl7dxvcGQAeRY8Gylzoawfy1PcTdqCIbG9EdGF
CJWGv8SahZ2M0wtt1kkNg2ljbr99cUG4QZC/34aJx1Xzj3oWqRR8DtNSLXA8bTw2dOn7AKeiTuQy
xLt7uGZiFInWs/fNSZBrcyAtCbR0Xnqr7Ews/5DQUKAsafLqh2akJAUliMx5X/9xTQQFeVsUN5qF
6yk01D+O1GtqDzit2pJw6qXhRGnT085lWincIl8Nq2EZTDrMBPsiVWhRSZOIcKVou6lLEuUnVp5c
u9clcInp43dxB4mLvwX9Nge1AQU2ov+FJ7USkxGIHaqIjqVLarrQq/wCMXaAdA7iclaqX6zx2sZ1
6WvLYda7qJA+43Iq0cnyE52oe77dgXEar7DdmJ6c8O05KThq+GsAJAfbCc2JYCe/ZHZf2/t59Bqb
0u27T4V63nQbKzooBWCQTSOvOP6w+XIrQONdTNfiwInOI+gDhtsUGuf8a2KIL9Q+W3gF21uzOtlm
UewiyTIeLNxvfHOMXSppz8bBLMKmVhfvwUlW5ocDXixN4KbM0+BBsABXjRNroDTUHGDYETW8xCUV
01lcQC0OMWVRS4FWbkaBkplJiglV6NIFGEtPQJ+rmXnEoqC1qZ8ddKw0hZhZ2GdKhxHf5ErZYdCe
2Cp/1UjD3P+ZnAJSCQRrBOB978clZpho/fWKvV38CwUD5V0iyZeh8K/yal+UZzpTNBMfINuPOxAR
D/QV/M6aHYalwcnnj8J9Wb2ho2MpEsS/t9Q3qdrMOhLa9LP1F1uXnzyjGEz6xQZsslJLmuWvEJv1
VhhKuzxt7TF3Ojgrk2/Xp/7irUNTgCoW6MDD13vJFmdlMkG4Eo/lpuLkMM1eKea2Um1g32BNnh8L
UJPKisg8o1qvXv5Lun4dReRAvUv9LVXczHox7WW37ybJaLqzKuPmC89gFmWl9MR+mojGHBj5z7Fu
gdboZTX1moa615JdHk4T2kXemTFyPhu2u5wckpauaw9zPuWpCAl4NK+4NMAlvIIoZG1ANBVdJIFq
+yR98xBmw7OHi2fJHg20p9Y7acT92P2yOwHUq7EC9F2aOY7ZytjYejoi8T9OcBdbMB1ogtPTpcrz
v8P5Z5a/dpG4zGvcfUpN4ixpyrUHF6TzgNCFpAJHpanbN4g9vUBrlYLt30ge+9ip45wYCygJvu2l
PNXkd/4IvFmqQPwuouBz0bJPuqwRcA+t4hJgQWTbDCFFfTKnAiOJ9HlXMS3vSK4Hgq54bNisaP9Y
su3euDQFs9tE+8swHd+TKDopupDJCStBnsj17HW9ZL45O0fiNUYYIhaKlwvx41w7SMoEQkmToW2f
Zs2IYV+oTUq5pkFPvCwpqPTBy7y8xUF9zBy9rsg1QNgTk8BkDTlgpNoGNTrdpkvMk1z+wgsv+cFT
AW5UyGH/6yK+HQbjveMmPlBEb7Vxs956518gntBrcj5HlHd2vrxYhfOfbht7k+U11WN2EnLGRSx+
gJ8qj22Eqav0ksJMSzMSHEFNxTcpzl4Ct/JZQtNTmkZjnCrkNzfJuL7XfWwN7JPHEHbDJrP9E5Rt
MhZynbs0t/xOsTvFWFasEB7zlgdyEZqNIGY8AVGy7HG6udQosQklCLWRQvZ/b1SHgMaS9+nRfZlA
40hBTzMEthsfSswfA9PPh7ioBZBoGzBhFGJUAd26Wm66FKSv85pV5VYuJQW7s8vNLqqn2WMM0pP6
hrY6RHJ7OVcay1q38Oh4p5LvMyqmGf4u6eAsyJpWV15MwPy1G+cDUUBgwlmgN+77kkD59GLMd9Wv
BptIzOz1GvaAQ95ON/fuSbO4v7sGx2FhkVCL7M6AS1yR08/3WeaF5DarF0fknFleiRzf2vkW0weE
abdFGcPHX33BWm9iroUXxt3gRfVRT1J/6vC0hu62aA6/E1Re7zkJ5bDhdyA4x1Gf20MInNLaQ0N7
+AfKgeC/Ewzl+HGNGpo9viH8qKsb1sS27kkCxLrTkykPq6Dkl899Av8q1mB1vKZjnM4KS3b+z+uv
w7kMLQxMAEIIQfUEjDJJ085eZDlJWF792l5ftEiO1Ww9mkK1bQ5RisTI/M4DByliVk2R/8OUv5rq
GuLcb2DIYhN8eV+KURVpmmZtrR2K5fTm/ohoJnjLYZ+mVsRZr+mYvG3K1y6lY87A0bHbE9Aqo89c
Sx5DwU7QuML9uIiipxOYCcuTBB4W+qfB4cGzkkZfbH8DHI2Y/iXDVKgMwKfsbD0NmO13G83H3BS2
aET9F2hCBdNjNavQ6naXIBGBf673iPfxEQgUL1zO8nqvEf7PLxmesmJvfQUHd0SUQE/BRIUjBwU8
EWETRFTeeQrf2QUMHxvxsqNGi2Rd63td2fY0vbJAoFETyao7jntfaQNgR6BD8qUbiCyxT0pGMc0Y
I5futot3/4aXs/gjcBy9uv6gMcbT+nOifSLN+Y2RBO2N1837CHPqRiGUzA0Gj+ntv7Yh69ql4dfX
laUMhkRRSHDyQ+Bl6zsjK5cvPJEYGSBA3u1bhSA6IOoYyH6FoM/GmcEUioA4YUTJiNSimMQRM7XT
BN6QODiyi0E2idO3+blHGPs2TLYw3zexgYQBkhX2/s4lntPZ0WdLJ4xW+pRqAVIUk8DQD2e/R+0J
u1eDg7MFrcsxh11Ejwu3XGzknww6k53ZO63HzrJADrgdwpkyroEo1fRAMnRFUTktCQKrH4tXFLnQ
nCm8pg/OtSbKFH8P2JkoQzrUnd3g7UsqzWokzljLIB8wSeAb7dHzMYSCYf1C648LiptyA+yP++Sn
iSD2ymG0B7yCPLxA3OptL7/1NQHCtOwJNvtCoXuXIjv2vfmlLP+qAf8usEyJYNiVPNtV6T0OrEWo
Q02FlNJAKfqkYA88C17sOYTV/fEvZYueRChfb7NSv1Yzj0D8x4qc14GSLsFQ38yFoG71AFTNDmoF
TxnaYJlQYI+y0xU7vTWy2Mzs6DCtJIANwjIorDQjKT6A9+HSFWordZzixP1dOlilDKWj612oL50q
+kmeyncSrCMMvwrOKYVS1lD4HLcHvtgs618cFNxw7tQSvq1mgz1tZv86WsauzBsBr85ZpZ+ciNlM
P2LdccE2tD7YpBtWLUM11A4Re/T69QymOdqI7/1J8+jHLyGPhU2bMj5jGl+rT5tiNHSawgdbmGfI
ZRY4sLWfzb43WCDX1+CCrlNiZ4XzKV0hUhqn+UukArMRsE1kIczsJ4biOtzkOppIyEzUuhRuJZG5
sZ13RlZy6k6ZNIiVbH6f2spzljGgJ+PepYpbDiy2vkAw63J+8f4smRsbYcULyKazXRwRjhLenQ5K
jzHq94HjAHPa9tfa6zzymtjKcKQNERpgnkeNoIEnQKC2JOoVtOIMiU3rRydaBTP3Gv5WNP29WnyM
QDODeJMgxj6N02XBrIuNemkDIja1GXRGtHOlPl1wmEwtwzN99UmlYWJxrSm2jqYYGIguQebnz7Bu
XlXFgXFOHEQTnb47ZhMBaR50sFa5DcSgfWg/vhoT2qOStGZG1GZ2VwS3CSwREI3rzV67ooF6ROZS
MJYDdasSzFpimVmw20yccdvmlPVV7ecV6w7Kf69SxY9Hk1Sdn8FByC5Gs2tPwt5aiQjOrJ1zVJUq
zerTcQdoVl4IeVLUbOGBKLfilJuOSJu0Pji5GsGQFi0Wps3UCFhxaXbo/duDZOEa7UPmbXfa6Sxs
hbD1EleLf48RW5iOMmiCj8pugL4JexZ4AFvAh+UMvYN59Gd31plMZRno/GvX4s2N5+/hD0atMBwA
uDTttANbIcrfgfeE6wJt8F3W0Yl/35pTxGtR1v+6qLQTm78uV6UWVtn/IzF12D3AOP1hFy7FdJG0
NQdlaYlU+a0SBeSAz+2wTPHqEXp+nXKKElfUcvHVsypbRpVr40g3KWTh4phAwfU1Fg21Lx2MZAo6
QEQDvJa4NzLkvBM52Gvls4rpLOTq3iHgYMFY5qq56V6oOZnEl9xp7N/a1ppS79ABWKWRaRq7cdGr
x5lzqKKHM5D5q5T9ArnPyDst5bVJ3QyMDx6GcApP3g/dxkMMRo8Y/+JRVRjJ+MP2XC16uwZmtK3S
ZYV5te6IELZdHXXw5K9HBl1fvRbHVVLZDCxLXLjzPGNZ8DFMn4XBxhC9SwwFmATpnUrv5JE+LJBs
YI/Dzw4FgaGqcp8OKqgGPe1ljPQQJWjFAXyXTOz68XncDwJZEa7/rG/+8xRKsRTKgm0NEKMCEzE5
fM3sHbLBd52gqpPvIM/luKp4w5ItImqYy5JkCWc3+907DI9waIhBJcVC20LcRhoQKvuE7gzKQh6u
nsR9wnEIaNDLuNudanf97rPXidPoBx+29uoE54FVGTVAgLlhRJum0AiU/bmMvoX24rD63VDBrD6h
E5cFJg6NDMeWlg2Nt2vNHZjxv5SBRiV4BSteF3/j9qmR/d0ubxt1UWgODomqHLrWmUYjlOUbSwyg
GFoloyJoepc8TzpHHukQbxLlz8c3nezkjQsT9V3v1Uonl+dqinGQjD6pDg7nBfW/TA0lNrQazj4y
bwd/q+LWInVg2dF4mJvdwq3/L3AYR7R0KWKRU2xA0DKscj9ZUlE80tHn6lCsy6tI+9hqwCPY5VLc
dS1dJAiDOx49vcJR7gfw7hJ070BL7ytP0u345ORqldscvX0tbTbYPFjlye27osKbj6hmXntQJwa8
FpNn6x44IXTFTe8Nlzwb8RNXY+NIr4rfBexBjEi1j1WZcs/MOzQGVHO8F0MYNB6RN9wviSGlNdco
7BuihC87fY3lPm1gCaHI6cjze42F0UxJK7mDahJ0+EfEJZrbCwH2lTFDuGRfz4WxoTLRBPQK1gob
R9DZyCjjEbrH+/iN60/+dWFejPB07k3uKaDYd0YCoEWR0mwtcM5kE4LE1SWPuZjvsvjy7OlKHMrK
FN4ilHKOkS0d5pztOPwz6WLw/064zT8A5yzI/S4mTx4b047o0F87nFyhT7/stHyV9689Y4wZbIAK
Vj2acS+R4wEIbU0pt5jTvyhCd7u3nGLUbi2TPevLHrfLUZWzl2z4uDGzl++8fR2SxR37TBsugOXq
R1Z3ciixHNuriubVJHJrAA/ak5fpJCm9xd56qGRDpVPygMt/ptnaeImxhVd/tUTPTeWHF1xijhNY
ivTZRTkBA67DmCtpTpzN8q+gv/rPSoBqRx/s/lNwlXJG/kMC7K+61WAiZP2LKXdO5+mCZ7saSkMG
e+sFNwl0GRFBWiTKYXDparlUpUylItfBXoEU9GhbkWj/z4Z9jmkHHM86ucyZks3eAK6XpcSeXC6D
+xr4547VCrtCXPa5B+5UITN+1J5BISObCIfiRvndpxIqMG+kvvt6GhPcnxW6ChlhvTfYP3DPi0dA
WqXeo6kCIoi5O8+H3+m3g3U2WACErfh9ZqlvezS1/aVZT2Ly/Z1UfhK5KKFXQsQq/6aKCJxiSeBx
5IcrWH47MGbfMjeZoquhc/jBVCw/UaovsBMKhgWGQS/4tFGr4ZfcIB1nnACZAbxRF0hXh3qML68/
qNHZJYRLG7G5WJVVUmAHvG9DuKOsND/PjP0LD6GFv/Gi/6i7EsFqfiDPxZHC9ZqkOsW6qnmy993o
z1DWLIlpFf7vloMQG7QGU1DesgNfw4xsUusClY6FaDgX0Aa+FJ3mjxOggfNcegf/7D9Bid2WL/d+
rKSwB7mnnHMn353gbx2kJiUln6fOemhlSw6O/ptKK+rdvDPnj5++5Smny9AiTvnF8niQirArWvqm
DzqPLZs+cF8fmDf02plYEiDH5pa4vt/M4OvHaygnCKiyM+H04YWhuGXwbHLQxZp4ulsX3A7U9GAV
cel0S3UQueytF1naYADn+WImCbH8w0Pi6saL1Ycc7RTmwmxDt6Ya0a1SkBAZIHe9ubhoZ003LowC
yL6QOpSBzVIMbYV/1KgiTFWdf9rRK+gYLjc8tEL8647HQjl84+AVVwwGZ2a+Jkwa50GLT06M4EEr
qQUqZPQm+qtD/1ADKKTz3J2CflpRu7/nHFzsP8Mx4W5OWRyR8Hwcb9UqszW2Ug+8P6WOFybPGiQK
ynD5K0UNhlYpcQzikabOF1V5OkizKG27Nl8Gm6b+a8payc+hBojYBDjj0hLfNbCF/YAknI84sizM
qWKwv02H7rpnuoP3w4B5YfUHtqCP7LIsj86KzWu+FHixPnV1Qs5yXiiitmIkrWpBLx+PvhcBWYGg
PMnXryGgxiUPJnCWevKFOEHNxlE00oZ2nIasrtGPpKUKVgubNyM7t88x3res3i30/Z0xAzW2chgh
kpibbgHbRgYnRYQGphQM7hHaSSVr7jBsWGvEFM4lGkS8CvHaIHxoPp+Iaov3oAG+mXq2w1m5Uvsd
gfkS+A3g0U3izbeVvLQEUVTbRV0eXoyLE1ZfySHnDH4SYBlEB5yC7egF20v9cjNlRpEkxmsPvX2j
0twVxt+Ffc5z3pN4trGsNag6AbFY8Os7BvO3EEIz3oICOQNCemByEGlmb/twOOLrymfYN+TROugP
unDl1SqZrHwZpXUy3Lb9RTiQabegktogoag+ufRi2F0Izi+4ZPMY/18O485UjUz6V4HXJjbodb89
5mCfygZL6m7yDAjFn1okleo0MXMcM776RSNKrgVR4qDR73VWKHjzKmEQhHcJ2BrGj/zXixn24Rf7
JYR0qOzReuFvh4OikYtXMqYBblpjucSHCjhg3nlNGi9BnNC80W+u1BIcm4b/Tlo0YNtb8aNjjSQC
El1/NZ3IFAQrdIeU5NSvF6PjYDQKBCyXO1PE3Q6zeA3IoubpkYfuA18S+oKckOyZ9CPe4w+HKgMF
er5I23HxMQT+VAAwkFxJJ46X0sS317FheKEo6fYW/HPHw85lIk7+e79uAhdPV1UzCAr1BKhFXc1c
25uAdSpbPSj04vYa2Huc/EWPkKM1XLrYOGi+THYOO2mrmTiWkHc89wP1VSt8k0j0GyeceJd6YWl1
yK0v+AaEBUBH43hjJSPUKotvO3HphR1F+fX0E7fz6tsMqiRkCINJFwOvVK6TRchu1CNTV6+zBxNW
G6eO408fT5/QgB50C6jzG0B4CGW8kfv35VN9twR34MLf4rKvhT9FyWBkwRO9YDS+V7LuKYeqw5Gx
MOvuR0TAyHMojNB4mFaJ8w2NtxuIePWLCTn3MhSZvGjPpVBP9yKXgjqxPLalc83HJ5JmIIREI+BW
9AGcWhmy3mmT/lBH6is2oAJQ8EcmPnpNHnMeFVp8jGX/laPcOHkWuyMOa1Lp4YO44JQvvk4CPnq3
+c6Z+c4g9p3/ode19dY6jcHmE2IuOr1eFPP3/LlMor/5gneAytn8l3ax4ocM5TuooxquNo1hoWnV
2+SJbNpdtt9VpU2hjn75gGxuKetsQMZA1DvLERL/WHK8EnehZClGH/5JO+i763CpLpExNpsF27v5
ys7c8UD4wPBUszR5Cu3xYn4wysoZkZ6GIpekleD9B4E0SrNxvMgaKvigdHPmEr9tDq7RN3ClTd9T
x+OHQBDAGYx/hU9kESRNoVoS2fF2ZnoBAaLg2g1wJXESV4GBBF2gjHQAySR+EKq2QSVwJc2qoSEO
yxzXvqiM37OIwQPindaOPWNVWLjkjsWV0fWIwdbu5evPGjL9mwFY0sjczAmSgs16yyBfG0tp2F0a
1fN6eieSc0SBa/bQZKIO/DOWMLKI7X6G12IVzE227PxholxJqJF7khb6IVtJ+jwDj4WYHjc0rwJm
0DI3KumTtLcj0WxzxSzNThEx7KT1m8xFWG3D0SUU8fzYai97MIexhoONgKSTEVVHKlP8m2fgvE7V
MFRr+oyW5Fp5wbCHo8P3Tl9tJ9v+0vCuMTVVS1wQyR0ybMiRP6ua22k8pp0dlgZc29+7J5CUkMhL
V125kw6sYh+mn0QAxq5po+cJOu6qkJm6W7FPi5R8tEuqEXSFq1EwCfaumPCGJnfQ2Fwi5+eNIcKg
nX9RwjjddiOayIQmaCiSopAcX9zXs1glzhPEL9bwuOYbN6Q8XpF0pq7ujlz2sZRXVKvFH/Zkmpwd
E2FP9XO4/w6Ja434ETCm0Ic5BXDWqziFTuFYB0kg9/0ry5JwP9nfHQ2FKBLFKCYqBQ8KOhIiGl2z
WjGEfsxyzyV2ivBQPRcpxS7/3VK/xFPVue/7dIOP00cgVQl/pColyE9L7qv+A1cIYT290gIxPB72
s196oyGCTbJIldOD6u70BW4UMRjCc2XQi06tzBOOQgMbHy0hxaHVTYVE5ej05e81rJHgUOUttAy6
G7TUCP0AYNWcUiGQfPjOr4FMgvzQG2rIO2318VBqOhtk1AB+uwcrhNpuu+OVVuYXx8qokb3uzjbn
Y4ooff3Qcj6ZdjyBScxGdAlM6sEkTUoHvtxLRcWnGEaMo3M8IhwwH86W2q4inN9aMdYrC+LL3Oqy
ExXMde8anZGx1Xa/Z87nSKOLxbLHJbbdUZiXi2Kfec/f5zbV+kLpFGbUypOjWn8ZPCMguqQ08NPQ
BM8SVvwvfLj4ui0nZ15tEreIi1DIctS9bFLm7Qr2BHw79GYhtplS7BH+Mu7SBD1nF6ILnIEob9RU
op0aquBsB4k/5PRUzRlmmcxmxWtBPadfoliwvPE3u7khbipPEmelIe2e/gglCLc1Cd5ub+YSERZb
xcOcsFzNISoLxRilexGwNt4gpTkOD46oUnAQZr9BJHRFDmuB8dYYuw7z2pjKFi77HXiM8OcTdJ31
Usk14LLVoVW4OaNLbX5QWSsu1wbhZnxpdbUMP5ebCatSa10AIWTe3lVEN53l9yxpFa0Ge4eZ1fbU
f9zp5pxr75dtADCA3YG9OMn6eyaXYciDWlBfl6LDRCrR+5Xm5oOoHXY/mfZCmNfAsobZEIySzaQX
S0NyDHdrzxlb7Lg/H9PqZrtPZe9cEvzvyJUI7p6SwmpwLpl73KYJjrCqU9UlDTdUI/QNEJVMpxVa
WXWyXTxAq71IaD7/0Gr9jy4fukBBCO8ayGfq3zDvcK9AqSySjqku0BxaJjqRA4/f+BU6hztlmlZO
7I85gb/vyWPpozwlzbCfCVWg6hjubS0vKg+KnUHzSvzqaEm1zqogjPIeOONyFrlideKvKVFbPrl7
FItXsDZuD4tEN/3kPpkWPw7z9/wHFdclchgYlxkvycdTaWX0wrDsBEGvczEEjgA/7eq9MRhXzMHZ
TmyUyp9jaD0TEnndJZZ8xv3GQSVOk3DWZgRsQXo/63V5T5xQ5nHTJWsOORvvjI4RPfYp5F8M7Hos
O7prmkzDI3B96REEluR1L8QG1sDaFrhQcEETDEtvdidwEEP7oOe7x6tZPvrJB3mWtpoXuTCoYKgi
eI9T0M/3QMVL9RpI3aH4vqkkcf+MWnY3oD/+V/piWqX3g2B7DNScslKygFzLDlIZ9mBDHLITj5z/
q+RMC7ecewyHaFRxhGuH6EtbWY+4ImF8iNSb+8ueyQzKs3xSVDUonvcwTLx3WCVUdxhLJyqGmLIv
5gX60UxrxnyHKXyBiqUCCbVzJuJZJ+YTwvBUqCZvd1jhIDVCFGG4iQB1NpjbIDY8fi9Jgl5+IDmI
TPLNyiTCTIqwLkzMbznzSCtOl5nOw/dCJ9SR6fAI+G8A8nxwSss/n4w1F6VipKHYCk3xpzHXks/J
iyi0bUF5bM57kmB4t/SErDQp9yjODJ0QQZu6y0ZSSKrcSnBFBNTUPxn+OKhC9jHYU3KmglEkgXM5
qmOUyNaRIrTZlote+ufp4qCc853Mtz9rb/Lia+VuaiZy7XGkkBQTnnpLJ1f5LV/zgKRxEV9McWWF
MgBQ9ZatQ/q0j3zC+vnb31KgC5Lu/w6yMt/3NqqqVwQtwMXjLxxpeOaspGoYFHZSFd4W/BKuWyiN
P3vgS4Ld+mXVvxLgDmhje1qifWZunfWfPQVMG2VdUm+DOB4eCDcYYXAIGhQj1sWEL0IJWhOou/6K
FgeVSNhVc9BZan5vcWqzLmnPdBVi4UBw9PNc+PgkTFSvk5CDY1LKJn6F8y0kxjj2io1TRRy4340v
KhLqr2dSHkDDPjeQPm7zklzgymkS5dt7aIZQcG97jdqnQuWOCBgo0wdrhutarKzwCrHodBuKpXmo
rDxe0Gor+GOw3LZuatvIKHNYM5KBLch+pd25LsTvYSYksUuPo7zrta8seGRwFuWVdlNBya1ze8gw
rSyPsV2n69QfAcffyukhmfAqiqOdTnJZtDLJTXauu3QBNZA4Bf3EBaXeSYXqJlOryT9Ye/aS4SLv
61aVAEJlYM0C5uU+9wkW2QkCXKnqc5J3kfhiIMwteHP9uFfZn7st4DoF/AQmqxy2KuzDv1YffTc4
C7GkMc0octQMAQI5Y8q9x3v3j/UVvoVyq8ybr+C1PlWgYyomrSN6+LmPEij/im0M04xEChYOyYpL
qr/JtNm0Dh4fU90ygxOZ7/quGV54qREmzvst2/4ZtRzHaFc/yOgFPcys2iMRV6gjYMG/iv1ldqJh
0vAk3bJkLeO/1aVy+quMvP9wwqdaqHOxnOw/BduiHfP7Z0/iH61/65NKwg4MvHZlUdhGQBZCBVN7
fHRmVgzzbR9BML+g/eTpQOhcErw+UF/Lf30i4ZKlxlF4+7Pxq7PWa4T70X7B3n3dnCCn2z1a1diX
v9umkhdKaPEKRXwovlloNnO6NfaJ5D7eQtueEBwHyhdw723p5wPMvOPppOHXbUQZiBGtIu6Yj13p
fQ2sCSMbk/ykhmy8EPoE+oIjwC+vf/QAIDLv6Q56Oe2MDKwSLb20jcxrHzRQarjjxzMUWtDU8KrZ
NN4WS2awRWUnEWKgmuIXNsa4XIG92LUM62vFYMdviZPw2EIqO7oJkoZ2U3JcQPUo/ptls1XBbuI9
D09cui3pVhVRZr4qgxbj2oFjdkGT3MYFRnf4qGVP5jdghOhmOY+Vhr6Hei4n8sNDn8lpYEPkIoLi
P/qrV7eww7XTYeFYLmOD+v4rP6zPajG1aTMY4UDyB5J+9gahFeJU+VFTwdnEzsAycRcEyIa7DoQA
/CuGcDxKjnev50v0TLh6ld6/Gyc5c7ZOu9r11HegCOFM+2GDj/q6AC2tIQJhtRXoqwbZH1x6OkxX
vGQ5QVOdgAfjmPhkP7+hZXBVRRCryywGio2TEMvt8eBZ7bQCSeEcOR4SjmtH57iaaXfEITlP5vJ4
FLYSkol8+iR2Wj64otLDRFPN7fLqWMNBVOHPZs7XpdgR1Q7T0EjnWX/WDLLHbs5chpjNG81hjwSX
/SP+XZwOSmRkwFngmuEcjedxTQ6rE9SWvV/RnArJMRWimn1q65EYbR2AD4pRZZM349c0LOtJw7QP
xpiDr0oBIpFP8CU3p/77gwUaDcfxoIPaiQbz+FCfbUPU0fq0liKBEl8BC4xDm2xex4yz1wLZkui9
xcFSkSKr4R9oExSWTVKTRG/kP/jdAKb5e4J74uwLUyYUpjEegGwk2HdlJbqu3RYywgRXVKUZWtSH
I4yFDT7AeNbELiPmWBZcKTxTW3WYVRosPN83Ea0hBh7fGUhWFhnttzjxTRVUkEBM+J+SDWqUQevA
AU41mRxjvG6oTLou/TG4IOBZWJ29FPywWV6kKz7BrHC2evV94UJibEYac3ZwFtGdJVeUfjRBLXZl
4AND6xzKkSOoFsfhuDiXiotCarPLnyQ/Ron7PrETomN7urNBSZ971/6A6M8Buormbn+tzqoTW4x2
gRxg80DlvhRpvdg2iVkHjNgMOoTmYjXT6iPTwyngRT6fYVXn9oBc971Dd8vmVSLD8hWy/kz2E1MO
1qDA/05ZdAuZH+2dhprfEA1nHN/NTrDLdWOOzTWmxbHHfeyz1GGXF11aIpXeRLAKDr6ljWa++2/Y
BQVGRb/FvM7sVbZ8kuhDIywjK1PaNqwV/VnqVQQqxr2oJo0xBdtmLhtms1/VCz9+07WOgGORq+9e
6PI85Mb6KVsU0+FGT/zt83XCHMBNFRFmnD4CacjRpqO4PKlKQ7Dc9HfDAHikUZErD9uVlzf+s2Nd
3GPruukYLWwzalGhht8jVij6zFjz0KdZykeVjPglGujmFAuau+Az7GuCrYOBqOrenmtLQISk6U1E
AkYNog40Ff7vVmKcYGEpDhBjj86n2zbZ+qpYJuMd7HqKHrJ3dalKhOA/oBIxn6gX8yOtm7ZBCuAw
MCpH892TPEs9LBqSJiS9h0xOSSVI32UijeyPnIWNhaGeJjyryTIXrLcSOL647pY7phbnByh++FeW
vvF9syw1NZ65Ep+uB9DlVfoLRm86z6VhMeq+BpAONR2SiXc5yitVcp5TlAffxj5G/Dww6nLwG4qU
xwXV1KGee6ZGN2Wi+ahBTlt6+EG/W1rRYHI2okiBWHjFSa0HzHKKhS5o492NPguQwaBZ8cKYh1xq
8iG6cxcDbu0Qo29SEZfb6/DF5FMsC+84jwn4ghj4RfTmlu6ZGljhAq19wNWosKsDN9SyqnKQOKKB
+nQKexXfQMyhK92UqmX5J4uPnbhMdhGx+iPDFtQ5kJlxkfmDHqVqKHTxNI98SBY5tQj90jtQN23e
sYKVr25F8AzmdHU/0PAZP1refhXLuOLULu4PMOQARnr7gMnIgBfGv9hPe21yRBmQCkdINhMMcGTa
hNAPUNCnWAqZscRk+jn9uIPpj4K/VX6t9ggfhRXJpqsc5FV9hXfuNmjevPeyzNf0O2ejGoaESH/9
KKK4scYQbW0x6B8U24OyhFZ3TdWizVClOUllItmWH8/XzI9tSjZpBeZBD1Ewm0nfiR4ObcjZ1TKx
G5Pol9ZRUKB3UOLpsIe/xu00SXLdjbCk0vs6mHOp9FuGHfQR39QxItQ88W5tma6NFitn6OKSyhBk
cMZONbmmZ2Z/Q//2ZBg/U7U+WXFz4w/r/wp4c0+oLFqfawg+sziAoigkNtMr4lc+Ihk+M81ah457
q7dJ1ft/a8W7ov7yxnmxrYtqg4k9/t6bxeKARZbsytGUKWhxMWcol9ry+kwStrxSM3lTTwcXNe8a
hVJ+tF84o3wSQeG8IQZQboj5WOhAt/lQT7xcrvA+MxBOnHN8O/2ZRnX+uQHMhOWx73HqpU6yGQyH
EUbiMimnMBIvOOR3UjKriG+H5lESg6dhg9+lh7oaTCfS9LYf8i7DVShu+jWvpSr7u+6DbXVLe80A
B8P45lAePxYmhU4zfNB9uXRU1o06LgHrLeE8obHH8wNwXi9nc3ZlT8qFs/xX35tZT9cv73vs1iTN
PjcHH+0RkvwlZYlwTFNM4tcG8RBgEJjjzlf5Fq/fZQB7TuhHEbWoGmK3ydDDjIdkNhDsNPoDafQd
XwvIZHqi35iQU1tvziwkn5JxVADl9qkn9+okplajeWYJElpVHtsEtxc0I9KQ608MBIOWmGyTQiA1
vE5CGuNqeGWc5a0l/8b0UdtGYVF5cJF8kea0PBVcCT1H5O9EaPq8TV0Hc5nxqTX1if4/87bo29OA
HHdvO+RF5JxW1lEeebI/9cwpP5wi+jpbJwu3Wdhh2yvAuh51EsOJV3tAo1ih0k9yQ8G42hayGtYD
yjbVYwkJm8qXIiOjQYsKHa7ELP+BSUR+54k87kQftHuGIwgCX988vhfkfMysB2+Ssjhhwn9dz0Rq
ktrSaONXDvwLKG2uzPxrpSennHyFDuDX9JKgvIYrEBYaGfjGGX8JYyZ0/pONC7GlDyMKqLo7Ihqa
qTnUKzKul22SeGqgAAIgAv4Oazrc0S2NTbSSA5y4/uxsrl3MJ64F1F7diHxn9tB2L+F/JgpFLWvS
mpiFBja+jZ3DHdlHS2q3vA9cHlh1upvB49akIXTc6vfTjcMvHckscVvkO7uI6HF0UHstSCSI0Ab2
BMjtDULM0GRd6OBLmYl2eAs1XSI6wICBl7W845GksEgs16msKf10fKggLtb6oTyFA9wC8DNZ/5ZV
GKP435kGcKGcpcXgL0NriP44i8N7bVNQq/gvoiqKNtmv0nCwvJYvLIf3WWRXp6HbPpthwFkedxLi
KnmI0Wnm00cWJSMw4M+j3OC71BCa3vYLSEZxdks/r4jXLw0rb4A2RnTZmUqe1kJfmous6tnylRx/
yHQ1KtUZiQfg9Ix8COJ2X+MRqaYzRU9c6ERwryojvBaqDfLNo3OzfAeHOXy2wG6X8VftPGfcHTFJ
xxcMMx9ybNLVXO1T3JAXrNlQFbbYXI8sHo/KmSXFI2HlUccCwKMS8v7WvHP17v5inGB1X9tWCICf
q4eX0voKmal2aaBYt26+L7upfg+npNGUpMYq6PegYVgMVlcbzSK6eWe2FKeHwbohU6PmhLIS6zSe
wf+mQ6tkuFUcEzzOqtFg5zNH4R56H/pjjbchMV1+A+9RUpYDA0XYPFfEk7c8ZYA5M5iJl59xvyUE
TT1wOUP2ZkMWcIYlPbp/BF1XoG4Le0u9m6f411jaGvCUDGQmLdZKwOTKmswFVxBDvEkycgpXbUmy
x+YHR0dLSGeJwXWuSujVTr7PFfR92R3CTtrGIqDbiENPQJvY/bByY/OWoA29oa08vArciGBFjy5H
hA9QUwBObeq2DPSulkyWYQGn4Mk6qOqU3L4e7ZLmu6cx+xf52W2otp7k5GnWoLAc18Xjf6wK27bH
AeVMlK6UYmIMcn6lnKOTn1Repmfp+0l642qSMEsvVMSvNoe0kxTdJep/bepC/a/AwWEPZKBIj3H7
YkCMxLRmUIh5QX1JmtkqcoyoLgcxNt2NP67LBYVV+LWMVCBog319YHUzEx72tNJaxddUeythKaJU
MxIUHEJiyWpmwwybgd81sFB8p3w87quq8Zf1H344GjOwAaTpxpO96pRl16j7A71i8iAFlqb4mBxQ
sc/iJdQyDTPXjnFvEbhj0n41Bw9U6a+gDw7tjbT94HEYkpRwIE8vRhxs+2jNmDK/0Oyz/IrXZkZe
okTKSSGpBrT36lq/P0H4d9IzNkKfV7WKdCplnAQ+1Jv7AnzA7OAJbrSw6xaqhLw7G5yPUMHyPHAc
26aj3fwMNIAeMSbuMlusbUcj06pvzPCMtnVue9Nn9FyZtAAT7lZDRWWltmv/C/dqb69vE6X9LG1N
LqqmEFN8zAFRtrXYoMP4BeI+imFjmQ35Kz07zfLhy5a6WKZugnnt686cLujSvjtXqihvbrL1fgTF
VLPAV74m3buu8k6kp15LlVCzSJGQRFInJPDDep3tk60WSm2afF8HSHBUQkzKTFc8iYU6+lsJOHnR
eDO1LHbAf/ui2VuchdTuc7rBl+6DCGE/S48WdquYGL4QnLTjnSDxUH0qN3KiwSbL/RMOybuYa834
xVlwqtoz4GheV7ap1jFy9VvVQl6pRL8kyQRIDvyGc5meBry6qJTP38YF6hrxcvCk5PBPm5xwPNCE
4jXP9X/6WdHxO0LnOG9tVYNtnT2OKPLZbRbROA6R+Nt2+pn/WTnZLq8WzTwsw9GrgpuFXPi6vjPc
FzHwtK40mlXy0W3dFNTHpRnYrT/+VbqcOiu0zwi+6gUPyAKEhiKFTh8lQuElWs1Rp7hgN8FQbjrm
868LIvkHMNs5iSt/Rtl40+T+G9FDWoiNkO+WAkFxAeA0JCG29xpU+yW9Fxy045EeJ4xnrDbEaiXE
rjfhKTwtDMtW8fgBw/Pogf1I9nbVQoHmtDXcqGVjHOQ2SSQTFLgNbem9nYmK1FduPirbsZ6i9Xvc
Ylklb2o+8fc+RVob27rulwN+4B0UjR2drACpuJAVIqEwtjwBOt3lAmVjc7HKAUiX+BfiwnbJH/sE
e6MWE6nij1c/7DDaIfF4AqL3JMa4J76kG1v0Ou7wEzHtKePnjYoa0ObGYXf3UwYZNXDu5YrYzgc7
TO6cbt/l9sMzM43VcmM5NWoChp3Kmi3FX5bacgsiJq2kL2sUE1Pb/VWskNMvSDWRwTNA1Wcp/IR8
Q5yuIsphyjCHZQxq0d6RvNYld4uUqVWyD2rOsZrzlIr7DeVteiMjnSGwGoyPnihGpyBceY9HbYBw
SEEjW9Wir2CA1iPA1zBvGp6Hy7te9AQasjHHKK2VfaNF0CvspDdrQwadeed1n+Iq1DaiuuCvNBJU
Iy1/MgcHsUepSk4wK/LkxtA6G4xkzfxb1pwvbU37OH8Hmvb49uXCISoFJxyKZgQn+/Rr/xQR+8f/
6mqRC5KOL87zcL6jwJsh8QT8gGCoBf87dmga2SYgg0wQEqlEQuStRy1PNmqT6or012UVYRYYXhCe
xaPw7jONO4NAfjOo2JpkIFClKpZk6B5XsKEeWdyI3cMhQBoP2rygMZPeF62xnZzqjMRUlegEegL4
ZCcHITYH7NSjJJPQf065btLpmb4IY8kB2akl+h5XA7Jrj/LAaYxzgXSEo7CVNDLrUu5A0am+n6f3
Z0qo4hrNy8fwMrNutKORBCszROotTOgQ+2/EaABMciuowNnHD//XL/WH4AhhBWe829BxicCVc3dH
1667BhmcTBrnHjY/Q2KNhTAAlDb8lceqhZMOOesjZJzFzwr2MDqnlTETXYZhAatlDn9BYrHzV+WN
tij4G4rbCEjqQ+SgTN8B3FhmI0Nr8WOTKMBHczICvotK2Uh1quQve4SSZT4RK78GrFhFdSQNcyLD
R0ba+Z6oIK/R2Oa5t7ofVRFzpEr2NFVwBSJiVFSV4Mugy/NQzTPjNUSENkz7QDNQv51buOKfSn4b
Fh5NgZ0AjVi6hF+G4TiLgAeo/FOo6dkY1giNBHOghHLZsQx4sDq7AxOplgUbda9bnKZh9nKq6TfJ
cO85t2OkMzdSjAEVohpGaEjXnMtaTfjYzFIjUonmwUXdmGTw1VvPx7oZbS4G3kuV1UMqWfopZTHD
HDjyt4P9NArAGYhgoMTNwN7MbkQPHLEkwTolC6XEfeYeMfE4/uXj1Q5ojyQ8FZzYbpEDejBTHk/f
LicIMa4NxAXPWxv5EEYi4UVIkTMPR+O17OHQCvneXSfVuMf2aXS4TF4e2abQbCqVwXaNoHYZ3CQN
jM7J0GxS/7HC8gR01XMmKGJ1POxxk7vAQlaUGEs0np3LgCD0zMn+GlBaR4yasTa8rfUW1eC39Sdn
/486xk3Kg6winz7sUwcF0Ls7jm7l3kkprb3uvABCHduNviQNVtljb/7mwtMb/1q7BdO1YQUHI/09
ur/qCsOh6zZaulFP7ZPAeQ8JNZysslAUkcaiV+Q0SyyP1vL70wn/YsL+/+myWnjsAyh+FpWOZqAb
hcwJZts20USAl9tZKrkW6YWZwyGmZG1R+eRWgI8jPoErba6aDObv/Q9yt7Z+HjaEf4QIC/82OZRQ
TyojmdQKzuJDiWSIUJ/HRNpHqSzXAle8lUGKVD+r8nm4w1wBNNGTJCRRE0KomZTWwTsfM711+WDj
8uKlZVMhmZWcpkqyg/jbr6hbLe61HpdXts0wFB+/+RIrp2C8UDCsy9JZdkCd7r8RQsZf4H6i5RT6
bomB7ckcml+Qi5lFsSGX7JDPOiTAt5F1YidxviUfR3DjVGSwRpZmHeNRAPvV5V00PZsDrMbSLNsM
hHdKj4sXvkS+TKTS6DXWCvrHYLpxBakBxhPbUyPTzZGR5mJUDidaHNIlWQgHbiw2eBkOsIR1mEF4
SAPuBUQgAmwr69yGtGdnSGPGtTwiRfte/6LoC3sq+5XZIdix01c3kxe/lK8DatnD7degz7S2Xl4d
KqEmkCRkQrooaXJrZjs8MGUKP8WQYgtl4onnYt3jPxP2qiteay64DGQ9naPK/e4Ra6y2A0NGhP/a
q1f3IWaTne/ldFUHrJHM17OCz1XB2EjtrI99eBkzsVPnWs5w//TBJ23v+FZQa9/JV87ImlO4kIQW
EKJ3lFg5Odhl4o62vaZwmPyr1fR/cpGI+4j42r/JQr7e1O6g1mm7XDWjtGIX6ilb5grnMA02T2q8
I+Nhgpb1FrMkpOhiimIeJog/JJEGxaCiuqvj5Wd8yigziAvk8PJgqOiXAUUK+aRgHFen+s7PKwWz
x+e577Dv2IyHXGhpNZUIvdrdeyZGzzd7+pP7F3rQWx72VuIxwu43r4cvfDMAcs0vrVPFZRNuFBUd
CoS/I70MdVURFAeyPN1Xwks7jm09SHNEhh4uE128VEBSMBvFuZZ5xFBfITBjakReWyVpP6zCeme1
XrS5FEDfVlJR3yw07dvYJ0sdsvsEWTtOEm9BZh3/p0M82SouHe2dZBoNJpYX8iNZW8fcUPHauzxt
06xtfo5IBj1lLe25juzsbA5gmqLhM0v/sZTr3zjt3nRu3GiHU70njytl1fseNhSdpwndpKNRsfmU
L2eeZMnfHwKxWBTZspta9frslTBBPEY7ZQau6lDTXPn5fIORyIYhA18HXXHuyeNE/4DbZxsjVIWe
fM91N4DC0+ajo2ciYp9YXJGY7ucdOJvDEw1Ib8UNWnVE3+8SKQHKP3ddtuufr69ut9AtGQyW6nTb
IJV3zkrhnUVgNayJ0OV93kESbsJm0uImXLhZ7Urb5Ovsp7hyjQ5rzPkS8CInMLfMCgl5g6Pml/Az
unoWaSqCE3E2jn6Sx1uib7bab3xNyrJE6eRNkJZyzHhqSZyRkwjlkbTYot1bmfJO30exTTdxFwiH
qmzwLvpo1LkGJ+OZ6x2e8obsUC0TQ2QXr0oVVeDXavvwvkarKSx132ZhJxNX/b6XyuBTutaIVPie
CoIbxj0xv3j79axLSk7KGMy/W3g6BusFJH+b9Oe0Mu2UgRiY0jIqQYegfXBd9SSS2UPoJPlvM551
TvW/1aythUmqez+y/lZxwfxJ3ODKW0ZoktTwQcDjuKmpFzhHL9MJROcW1BUknTtTvMejhXrEqvnz
FN6oS+aQuytPE1+n8v82KPhJrP8l4wbsEbu4Ve5eeiIVYrrYnmUEjE2vnygFpMrX1bc6TEOEAvfQ
2q8mS07JIpz02/NMJeJ1kyYrH6LSfStyZ0UQC9+oP/R9OJjoIod8uysLqMswXbTMK45/NomGESh7
FTb9CE11li4Z1puHMlDm7ENkB9jDixUcRfYZNfMxY3c+6m2Wh9mwUwPYHjI1wraVKIGDuEG3yMFL
JYF7DMD4UzvUnYJEjjpWbhYQ3QNbeOnN/4F0jptRiLKKU46DA2lorDPWHv+/WqsxDRGvx3vGLgxe
45zx7cv+xDbbHUhvhHkcLSJVIjYkKBIJkXlo2bwdt1ycPM43nfStUoOxOhHQnUPzIxg1ygOHHPok
ZqJ4SlunEwMwW8ngaytQhzx8YM6HdJHwU9Scc23kTkVtPQ7X3uo0h4CKtfc/yCQmLuHXVgqXvf1U
cYJJPA3lChesbmQDMsI4N/8snC4QLprFGkvmGdXxzGvkXmivuohwC3g8zEWQlbK7Vpqbq9hiDd+V
uAAE2nUQIrbvthld5cTTNWzj1Up1kk7xKQ7/AunZ//PL/uB+kGkGteLa3ewm+1ZWFhG+BNbAFh/z
wQvvsT4DdbcR5q/5i7LCQ4vhGqeLPncpDjpR/sW6XKgJFrEMD5Tu39QuU6jS9QTBNTcceZ3ENhcx
G0dWIFHF6pQrpL5o1+TNQVN32rhoX9pMbtzyltuRP2+b+MXHzdIIxyNR5RZaStoaIbgX38/f76b8
Cmit1Vhb3p0rmR2YYuLbcN1nQyWuIwOUXezdrO3XN/BA6JreGc87kCXLnLhcjfQ2nVxcKg9kr+Ox
hp/nELk4MvY2mPswZq2xrjwBmsumEttLRQjwdmJHoKLBiRpw8KSEWXvIx8YJrsCO9BNumZsBl4dj
g/vKZ6s9vUuEJO2/nclb5ZLCD/dPBusgE0Hv1+vj4QPNSAn1w7F1VohU7EAAQek2YiEQHSB2v4uB
Ehd8KWZ3GZFwKcuJ0NFfF0T44OmaCG0dNW31+OEYmNMlw+dM7GQ8PfyfvvTjd1Un+qdUs1qoNaGP
z+i53THPq14Nh3iHm47F5IrD+2ZNUeH4lrt+wBUDvVitg1kgC//EOyV/k3x/JHlq/VHgXxNYOE/u
G39BeUyiWlQEXrh460h778Klb/T0W3+RalTOQi9B+riOZP0+Q9vnbhkCLtfc+4Fjbhi/Lw58sTLe
7Yj3mM88q8eIVe2VjGxGR8HmUGeG3DRygtXR1Q+cRe/4mqMShplqW0WyYddA96+R40dupElc7XMe
zLsa6zP5mUO5Rfk6yyP8xbWWDo3si34aFeylHN80jNToZaTthRJuMAN9N1i+0ALTLAL2LWXOgyak
CjVmKqMMI4LBoMiKdlytJtcvpt0W9oZ1tTJ82umXdLpe2CvTXa78Fs+npX/5Bc7iRIQtJCxFS/WK
uX/48/2mypSL5BlSW7ck7rUxI70Gy6ipVGwe6/D0u9FWpUWMm71mYqKbFXQegOmgiGSZQtgJw0mH
o7ZACFEGXAtYHNte7K1rbWvF9Z9yv2BBXT8hE3pqGO7Sh4Bv95cA7+FTJS748s+G3V//eJ9JXLhT
GGku1J8YEsYEZZbj+3Jn/uAYkbs7S76qqIM6vFvXpns3oBk+IgZ40/egM3/Wwg294fqvStKFR0Bw
FfF/9vxwxFrVWewsh6jP9fBckYEOE9Fyqkf51OzZ201PUgrzKipi5ABEKZz20FKz54yUb5cSX7oE
NzTC7dEb+eYQTau7rlFwnauX74FQp6pJAv711EDa0fhmyaQ5ZQNv0J59W5IU5Wc0ZR6mJDbuWvQ7
k8UeIERc4Gia+Eqb5W6HErH5j6iBB8uOeuJQmngwyijoUCQjj71pM0pa8st8DYNlv6SD5mnHNSp2
ZKGu8tmUUIHh1fSKgvu7khclXZr+7l77x9wSo3MWXzP/HMRpEsxKEnNzuG19Gjrx9aHIKbarhc24
gmSBPQsFbyw4sw5Rwprte6+Xy5Bx9Dh36F/ttY89sRTZGcEE96XWEvd2F1xWf2xva0u5cXlzG8Vb
OMGJR092Mt24XwJ0fz3DdX7mVijZYdak6kyocSMLgEXJrSEMZqDfkJx/MgictfJou4uSbTx4ZppA
YrHLLwIDebwo/unxnibAlIZy4A4kDIY0rpRV0DhjDvkZoRaFP2CEqaADYHcNRmL0bXKDiNXISrYc
FjEm9+DioSfdBY8m1a8Fof5ssV6976od9GwYqtoI5xZJGS4ylsyj2XGzYYbCg2D5BIAj0GMtEXUJ
4uf/nyIqtNtaMVUrw6Nejk7GZkvbLyBbnsmfKjd5dpD3vTdN0qQFIrmebgKZnitMbay7ppG2BL1u
474A9iA+mXSIYCDu0LS3LlsDpvX0Zy9nWtI1xGm2K5QweJEdUXT6sPKrnmVMakvcXTcMPHddxwmW
/ABYpgmw9pOPZG4pmtZfqmz89gReh4Fp1olg1vGAJpoPF/GgZ2zTus46pKpSjvZFwr6M1HDZOZHX
99/WMOgUD7YInQZtVoaj+PBTVQl+NcretuOtjfbbpdVZFhzAz80EKxW8ATgctXgjRa/N9IqzNk5W
rqTGCfxa4S/MVNkSWhMPg4tKmDRziZ/U24TLrx7Lo2NeupWdiTY5mDs/+vLDq7QswoJk4SEoKU87
0YfdUDXr8w6dUlgPTxPo1A+G1lhJHjgXDQScTAJyXaCLVscXNeQRksaoUJW59+TIAd+0lMRDQAOs
zcP3qkXVJwn9Q+FtURO1Fd6OnkfLqhBnK9xyqZ9AiJfVB8tu2ayq8sn1VslZ5uWM6bM7sBcYs8hd
NXyMiaLYtI6/2IaoITnmq5pti8Iq0Jzhnrh5SOJoyM53gvKSqkwl/9FjOmgD4vRQET8rO8xpdXZd
TcXV5gIIzm5pjuVbf0XhnSUQ7EUR3AN9dxNCBps5+wj2MQuYMYt3NgC+BJw2Qi5rbzoIXPOeK7wG
4oMv9PcIWGZhaj8oA5CKjS+3fF+yOYg01Pxz7wzqcZWRutIn2ASLs3XXiC9u69pi8o7K14dRQsaW
EbdNoy3dduu2fsZDQ00BlawVz6LLO0l4ITm4t9GMw3/W/BEKn0Ecmgs+kew7ctbXT/LFdRs06T9j
HWm9b5VPlRtyQMPMNzPIfyjbSCWy2RGYGamThHtec96AzYEmN/pkiT44NiK9yZffwCZTXjJU0c1Q
8IBBDkWUA7YW12x1qle3s9QvJxgwsn4aA/UrFbicVBrUBiJwCI+/PEbRj0uY74HAObvTsOgYBaui
D6DGQXata5go/KtKmnJkzV/h7bOBc08qqSjlFWT4tWrSDfowqty0n9pW9JGqyXciQjAtl+1n3o6h
OVD/boQcggSb9XdThE+3ZGs5dJubLvo7DhJtFZXrfxb2NErIgyG8WzCFH2Evk/0wau68p2oB3TN3
hXe44WObfnakeabcyHY6X+qlHwcR/MObTRVRnYeq+i6p5fd1UeBzAh1WdTpIc9IuD8wSm+IJPLY7
vEuiFjSXIoCdGQ1JT3ZpHTuKlJ0Jz8/fwa4Zx0p6lQiLyK744yejREWG8sY38cH1YpgSCHuANfex
KnlsEtlsCgNtMIUBDinONDCqZqT9kfzjexVI4KKm5smTH5iX4n7C5LKzLVdUwWZ6al97QC9zvapL
8cySmWy2Dyk6n9oU1OZ4eF6uHUzqgzn8pxZ0G63QOAIVllXqy6jm13MPCO0btv0sDNx/pmxMJepg
ZU75D7c2+/whkhxYGSKEFY39M9Ntwumx2HIIb7OqBin88jm8X/aemUYG6qbR/f/82+VY2u8seMy0
P+ecORd9bo2b4tdVTetYXBGn2zYOPyRN5zM/tBSSW/7T9JoY+gXf2BZqTwPi83Zd+DaTUjoCRIzE
qAgDxiXLrM/Jl88ZQVSZP9tENtKZ+r7r37UFYMFfpOee1b1IqNIT0HPrX1HPpsXKc9TBzeLqCHMS
BPniengdWm+6AoLAmb9rmHG5aUgL+QUMaUAje9k2G1CSJ/k+skf9hwZ4avenmMCer3t2LPTrZas5
EzSeGswDtChdEMNN5P5zuScaaMWo4uEWjHSCi6Enm0wF6/Ag/wlqftLFimoaWGfi6S1VQpiN7a7q
E70sfAYj+sVm3SsIJ4YumyAuryFAnMs77AVfZj4QvBRvtyxt/xSNg9l3XZ2lZKy0D9vcZAo6z6yy
AeYhnGmotwFdVmCqjEswheon+x816VaOFtK2s8L4gw45/Gn0nEgsDzkHQGYI2+tFq3rj91JRdMg6
ebmVBZTHecT3SxbiOhbgKLTkj2fIRsCFHQj95S5vtMhct3uDTFldl0wurklskLFEApW1IG5CMAS0
wt3ZR9nvaCGB61hABEwbS/rF7E8mi3XXyT60o/02Ynz7YYV+SRWe/8SQ8NXVdWaBCyb7ozQ8HnbF
l2dahb3exATh39REuFHkcJ+kpwYBkT7+Sbva72I1tyDAHXlCyBHzgf9IU+SwvIyCnuJub3X8FdB9
C6g0O29/PsxzVjDhdxu6Tm5FP6l+Qw8x5dtytOhvuxNWG1F0zBZN2NDRLGI65S/n8QTjxyx+OQbi
bLTtSB8n6ofGP1zQaYHrp9uUr4bBRTNf2OPqc7CkVxOFOc8rfpd3a612SoQNBXmDTHMHhX8eLNv7
ZbOMkWfyBa0CC+6AhXUA7RtYH6vFDpt74FWSKthInhoyoed0SrhEiUQQ/syDqE32+uusu497Vj9f
lQRTGtSZ8r3jFgjcTdQKMAcsQH1kj2I+36CC+P0kVi0KQX33eazgC0rJWQo3OnLLsP++pJvEyQuH
oU2AtrInmXFfov9pDY7Md4ifNj1AQoUYtMfObY76ViQmC+IKW48VQxE0C9TVB6ucqHrqlwyQEm9W
Tsfh7W8WcV6MGtQetzHmRPkyodDNmCNh6ljQr7gC4IYczS7dAzLyOVOf2so5A2+N0a2vdKG1Ttu3
NPuRpIUgxA8Exosi0SGNS02Nfrtfm2/YlTM5tOATZP84C7iwu3B8VUknohMgaVZ+k6GM3EzuESuL
OFHZL77J16WffCxmOdZTrrj2W0rYfVrNNH/uLROPefjsE1CWJmLvvhqek8TPeozE/VtVgCB3ywuW
x/pUwtDJUCQCM8/5xK9WGzDHl0JfGPwMmFT0wOhuFhQyR2Q4NWAgKlhe5eH4PyHbe2en+4supnqq
vCW1EQ5TwskjugwZN2IBZ333W2MQgMqnu8KBOrjWl2FPCiWCb4oc7DBwsd50/uAkVrCCI8cOWQZj
4I5+tIxOdRczkn5mcIdV/B2AbDS1nwQVXPPqlk7tPdsN+DB5aajkyd8YmKkfZJbnjJG6NZzPymXa
gAGrRSkjyOVg/kLS+jYNQEI03IzGS8yJupgXa1Ozv+3pfDM4P7is9T/k/M4vU8iFMJyeUu9BJhIW
g4HfdDSCJEiN3dcIAxwjLbEO0n81B/Zf16eBJ+v6ehtufuTL54ST7WMe2VFR4GJu/KZSYxNmnAfZ
ERRqWKthNhy0uhpvRompIzOTnUTfp1BXtx4S7Y2ncaeAsc5+8vJVpjBX3yNlIveY+tKHUJ5Dy//w
f6/8a1V1KDAgRu9ooYuQpHsDu+Ot184wU6zeL2z7PYieNa4EcaB081Tg70gpDL+nlrOJdvo2WmKd
OgcLkynlHe0r0+DrIxx2wGZPfbVbJ8RKzFg2Sk5f+i3gDN892wJWl+qTxD+nnOYh3stWT42moRo9
hMhVZMTt/5E/Yb8AT/33zVN3KhR3AXriKCIl4flaqWEn6fHaO91JHwVUI+5M83Z2CthRx5vfH7zX
86Vi2lPk8Tw8RrzEvmOBgv0MDRplWHNL///qbbMg7DWCQRbUAbk5hJy0veV+0FT2digsKsjmhyEg
H8T+36RZJiVnDgqdZk66UzcC/QCVy+6e1vAycLJ26c+/aNN4mQ/LwZEeO7F4+SezenlwZ99AGsrB
B9c6UXScBlylcluvzW3rv4e4aMMgpGH0/H3/7+E97G0eP5byRvKr3AUWuyiflE3VfvY+OO7wFr0i
+EJdHvEtfyzqS+tHhDlrqPe8aGaAjBxqSgoxE+kI0t8ifeskAgmbWsw1Dz2n6M0fvkJuhctb30Dy
1YTZKodb6O+zgFRYs4v1adssTviI8Etdp0aQBZVvYP2Zg87jyrCY9AvUfx8tWOzYJCs5mEbDdePC
+iakNkBWACp8GMnyhHPXl+tW0a0qGJCS8ULy/isof/kYISuP1q9roIK/OFNe8hnpT/T4cnSRHNR8
C/ucgXqbVNLq2SuM415xFEECsGaElmpdaeFcKShDgZrEg8sWdL7s/CdxDicbRz+wsZKLdnSERufH
k7WHCyAk+/4EnaB43IH+Fs7zUmgvDvEAHwXc7NyylYH1wcMZgnjKnWHmuhaoCtaYCTvZvRqNkMkx
jmPog5e+8K0Zg3ua8AAm5Ic//Q7NW5HoeTcm8+PBaBJKlx06nhgQG4gRfMlbtrDGyjRxFuPha02Z
BKcZDgsaepJxy/twTT/PvuY8zKdl8FunjYLg8lQq7GltM3vj9Uj81yrhRQVi4gGl1gzm9MVXys/H
UgMfKLrhyapGISqaSxlT3HetNuee2rDtV00LbdUSwPCZY90VoNUvsp4+W4dR2M8SdPeTMfZCto0v
6dB93TRJO7B9ULDX8I0o2dgASHlOuLIfPJlxrdI7xgO4e3Da7fXNg90XU1rf3cfTIA/JDUlQkUyM
gy0cZ+G8TDUeD8yf/KHea+irPLUK3vLZAvoXMe3NccHa8hT6hQbmKz4ZM3skyupb/Yil++i+tJRG
JjPaiR808pQiD398EAk7Ko/x472ZCZmoezMhXBnPJdxVXUpHDZ0haPpSF4+V9UnusBp9gqkQVbYl
DjQ2aLFOhx08eoK7GsD+r9peYfQcVR0ZymrXx66Vb+Nc/mLyscrsATX41Qu5mWkzsV/XLgTOPQUb
PR6d+QvisGD4GyxVHN8tCQBecYvpWpy1ID2xNQQyqApXOnhrWJISTREMtLZ7kmf7db4vze8O1eUh
5yeYhI/8VczM+hmZ5QnDgCqm/qnJWQjKRek+UVr3FaL+M6garM9+LlF2ZLOKv0gDGS/K4+9fYr5J
DPyHki3TpetY5sXhPTK7nFmwFgKvE5BoQ7yoic+YPL2Wp1hmdNlylkjjlg+2NYqUEiSWLSaTKV5L
v9iLzqr6cc/PCWRPLyEfDBSdRO9+VazugmzSWRfP+0Ifhgo0ExxZDY9Kx6jWU7KgmPPN9cs0XmIM
NFofxEsWwRCvK3WolhlMI74PEwBbBytx0tHMrWecMwEs4AkTXynmlU2R+vWBT9cAxGusAaQy+JOe
JhwDc8Z8mxsmcc+I58o8/FkF292v8WEan6ZQQ/k1pskrCoH5Xl4K9gNHU0VMebzm3kWsxdwYEFRr
UGdFtqKNwoG0DmZtmNGILjRaTpAOsLoFMFpG/NRhc+gG1AH6CBWU/LoV/n4iGLC1/nJreNqg32aE
20GPYhHjixyrM+lFuxANadf+FKirDoL1mAnEU/Cq9NxpsVHNouMZYepufQ1D9kIeDIpxHzltckSa
nIfER8jR1u2GTCnN/TrpoILIMN25lS4avALyTuz3X7a9RZ5P2GCbHax5OaCmvO5WyNXIAwNFWsNN
xULzryx/klMhKoVaXoZCo24Tu+6tXMagUB+lkF2xkyTDO/KZFtSE/Um7tP273MZfA38frilbKxVN
fnbpbEP4hdCyR+LkZOE6LoTNOG3VbFt932XchaPJYJKf/x83D/WCfUTeNjREiHwaCu8idnZ/Lkf3
GdhcXP4e5j8DLYp7rRP5ZgpQ936hK1gtwbIyqhHOOK6DQTgZtk6qGd87ZhijLy7deYKs6yeJxP+0
rBC56vxIhgF8B/5G2PPqHy+Qjpe9woDfnZaYJtS2QEhbB7Rx+VEsAkVOip8WkiOUpvsxBSiTSRdI
GpK90wFmW7PCRPSMVMkQ78I7l11gvLTcek0UucBFwEIu34Dgz4DgnR08pVd3DipUxfftQOdz/yXd
0P3/r4rVwEHoIzCYsFysEcAXGh8lplIapbZ9ahydxuCvag0ZItijunrIkDEbOE/BWkE+p63MmfHo
8YISMrI++EIsx8O3TZ49+A3zgMJMWqCLOZewaEzFWjjbyWsmFC0pfp3GCOmPc11+FAdHtzeDLpoB
qAYtcFfq3uhPIekK8HAyx6m2KGQtRnUsXdmnmw6OMM9yxk6YfEahfk/E+H71PGdrxJUob/GzIz4Y
FK6wVyn4T3F+G/qrEkyWmohsun8DfvIxrC1ApswhvdFYxL/97RAtzr75YrQlm3t43A5aeb2liNEu
NJ+JexfgO9jomYY626Oo07cPvSwFpy4hys2vH0l3ANG7GMxOw8B9spmV9FJA43x8TxVeIjX0gUjw
9aPKvdGbCLhG6VElobtqudjXFtg+yhZrzsSKUVqWPvM6UEBRA9s/IwiVjj7cf/CKg0grwGVefH0Z
teFixK7xMjCY5UPuhYm24U/lK2+5sWHo5SLynmewz2OxALZ7PFYcNqdTmleMNizkRLOqy7OqSxVn
jwNvSaaP+c1E/HU29tS272EZAlJEhzOJzzZYuI+PZvP5kG+WeayS4Ha9UwUTlX+AJNEBeTH9qH5E
DHVdolYOeLzVNmIaEEjbkTgqIycA46Mh80XTziBYdYNX1+22FMw3ES71xxkgP9p6ZBLXqEY4/5lQ
pXanmVBJG34ZBBuVgP4TBt+zESp3OWykh5WN4mGmZdiDrwLLo+o4R13DmWPcR/4PzhBl/qICdp82
PCPabD3EdSycgLgPq9OSWd+/CEDPqRZen4q5rdkeLh7Df8tOvU5bKzwx/blPiGdFLPw4zNWtdnNc
+cXNqhk5uGZePMYRSgImlxMTtPdpZi4Uckk836ahOZnQPNDyDA8/yhlQVol3zjVzvb7rC2JPQUEH
nggm1qCqxbyNeeP2/hJvGBzjwERaV9ArjZpol+RbB7AGD5UdRZBmqCgtt7Pmy+rmP4jrlOnPqSAA
UGDkUvFpfYJbTceIbD39HDqzESW6XEZYO8AHnVPKnEqzDaNRwtEzDvDD6aqTrnFhnQhuRHvBtyOl
JBe8na6Fvx/a13zzt9OGmxGYgl1jRLG2WYBGzPIoJY6iR5yFWpKj0Pdak5e8BQEmsn8/1d0MTTOS
dQH8uPbLhJC015dtNBCFpkBzQ4sr0On9ddzJ2VSNsJAJVO7Y8SkfKUl0RITYhYJmCjcxqi6mvKJq
UDpyzht6ElbfFsdOGbNS2MvdBzDKGwgSlVzlagnwV6AlIH+5VfDuCXmKrwKyOfWbGoFjneaIx7Cm
zXY4sbe97y9xxhYTtkKoQg3ruGQVt8iXLrMT6te1n+O71jbyvj7oBRkSK5E31F9GOZ2VpvGy83ss
DgPtuCVvvkmPJFOmbZXOULMQe5O6ydwFyk8cdfxzUtvnJd9CB16v+QPxecSSXKGpZWLTKpa3rZFt
ldgSuDrAWj1QNTUASzUT2fySX/hdwLioJ4HPigMjlD5dB1EScEgYvUi61a7zI74Zp7SMwDEVICeS
c+qp1DBYyh8nwLiYNWzdxta0fwDnyC65yFsqx0opz/68kE/SvTFuDVpliKEANi4NH+19KBs/cr+S
h50qoJlfF6fXzJljumXCcfh13ghpV+LL6uRxnjbE26l7Ds6S9HwvZanj9/BS/CEr9/On6FyxjFEV
yqihx6xR8018FmIBfEed58ql55Q63aw7vt1n9xk6DudL6c9zasX243jQvidgGnPSwUc7PTrh/wgh
5Hty6umEyHZADiaCKbX9XU7idUBX8bqDVdxZCInWNrkr1D1hcqrvbmJzAYNjwwgJcxg5UWYhGUps
qDi4SiRyme4LP8N52wvMcN/qti3gKd3YlksmcbE7kzvaHx9ovBDNeLlT/RdseTovmE0P1UyUeayN
eLIt9BBbN9fAuLwXKM3+SLvDalFlDDJQkLAmRIUNXVfUAiPS/YNOO4y+Be1E6BQ/SR2TfV5t9+aa
mhJMH0fPdWuPU4L7GuWczGo2pO0AROPWesRnMnOppqUG+gToT+7oi3ksIQZhPPzbnLF1uYIG2ehC
jqCwbecDTFPaBA4JWhzLiEuJecUSPcguWXg6A5oMJ7c2m+KmqHzBVIMtSeaeMnCB2MJ+ibuB2c9q
RjXJ8+6pMvxr0jBV6pDaVir+eFGH0MPV+fKvDlUN9O24im53gr1GJqJL/Ul9vksuS8mqrbNrlmWB
2K3TkRCEuD2y3dqu5n2g/0hs9/QhAcNlmWAD+B63ZxmY3E9L0ho8fvyeRLAXkyGUUVSp90rpN6zl
2sh1+TwiLe6tRqbDflpYfEdseJ9SIAZ6EVRnXdxZpDHxRJOajLZZD+ZzymzoTQ8JpUa9s7uyqX37
vZTGxGgY+2enb1fSkkTy/D3n0Gw8Zrvgz7h0na+0TfPKMGLgelgTwKksXrR9jWznf8Y+utD/C6Ip
pfUpan6ImNFrioKlIuUaLoAYPh/u9jWqBb4zVM50GHL5mA69MepuSIqCeoLJ1y/xen6mXmbOUl0o
/bxyWuAnKyOIGZS0ZP1REozOfamjSew8dkg5NzPO66rdK3gTUWvjAR0VrcA0HRKfb3nzJYhOgpvf
kzvDXlbczA8Y/T9l58c2XyJafH4zqiLkqQHOTCnL79OFlpZdy0jj6BQ28CrW18ngCyjl1XxqWfXM
Lisj0Ryo3+U95NFgknmyQ9Znb+KGcjqi3aarrbgh6xykQOF5sTvrqlutdnXWbbc4C/7c2CludOJG
NmktuoBi2gp5cxY0T2welf2yRCKH10sCtdsem+RbFhb8kWBFHpJIXnRDP4wQ1NOcg81TLLn++iy9
tEdjMLWlSJsPkC+7Mxs5wenmqnpAGNdfyZccqL75l2o4GsXICF6cUi+wP2nUjx0mEyOWgOc9wnkd
WLVczccCVnXG+Uac6TbDkD4MA/wg2Pe9pMTopiCqY+KCwMAO2pNPCcOVVEfquQFfQ25fDenpU+6D
uFxxPdZa+NFUpn+kKxY/sJk7mcejp+02AyB/Ha+GKn8mFhxSuhLkFuM57FRWY3fRkuRC/z75tVGA
SR0Hr23NHJPDgh5RTXjLOg4TA1UJHepQbOKtItkzRwGiXHGpblxnWt9i7ZESCG7OJwP52wHi9498
tKqhvg72MEpAsCD9mWkTApRPOKLgUb+RQVTva2VLzQmMPGEYQaqTJ5D5X7kDFTWafP0gXf6sifp1
06ro8P2qyD42HWt8aOcIaZzeVOwlh7PYt34E6PxtdDfDTEqkxmfyxVoOAbaogdK46KAcY0eArThZ
ZBp2rHI4lnZTrWFdsXVDgCzO1w2IcLi+1Nk3IeQQPJA9hR6wWy+AMqfuSR+b+KUloLEn2/tVHomm
IW7Cuh7oB7hbMBz2b5WPQ+43Q02w966BDaN5//64bUv8HWGIwxgElWPHea2qFijGHNZ5sSEHClJ9
gaPvcu22XexHaFfvT5ZiLvqgy5XBA6MoQqlqTpR5AK6ixnvqFX1/q+fOvPJbio5GZtC4ew90A8Qg
Eaocke6sWERh14Rsg5sXotXjDrG63OjPzAqV2kuBiMe9AEsNCG2fd40Nyifw+0wDanLnaqIrkvgM
8zXlSgj07R2kxgwGhxscwRYFNum2zFyjM2XgGwOKCkuRWQnMh/LtmQ5WwwlUN9rgGZdsRFa9M2fc
oqgT1i3En1NJ8uNMGnoOzxDs10ytr+0DCiOWCW3gLLctHo+nevwBmiWzNemxCaaqutWYCqGAvbl6
0topAV04iagPMK1TRVQY58bLB0Tr61m6KzmxMz9ZN2FLH/ZgftjGNZC8c+19Za15DJ9gFsyVMFHv
pxB8rX0Ku4olh3Mq1uAlAcXTY1zPftrO/M8Nit28dH7By1s6EDhTqXM2Q+H9b6CW0oQyspOJ9GRm
4Ei8zd9GHGJjkCst6I3cHNuOAWyYKiSCH5V05HTLyRL9TVYRJjdTb6NabUC3rvJI7We8R8A/qagM
/Js10sL+xTJkQSpvModn2ydJClcp+IwmN8qd9ytlLhuoss/bRTqhBr1cs2H0ZbKH35aprB/rLn0F
whLokxIUgs4P/P+voZNT+hilh2TTZ5JEc2tAD5GrQIRbP7HQD2VGAWeNNdFMZlxpChPRQFK4Wxvb
ukeTXOhoobWTdjdgiyC5PYtgNMMqcVP0tw34b6rz4S4gImG2D9PTV67ku6904RmcgZP2oNsboqi7
8tM2XEY9XuQqvw00VvKsYbnF3fH9Rnr2XADYPFgSe1pFGOjKNB3l/KlQiDO6CCRLiKyufd95V5Lu
WTjlh38r8E92M4DETFbV6WdGZzGdSsVQo/dAiuMCCL4HNKKOgDidJPKvIWiekusTq4d1SnDA26K6
3hkCpO4fLmJYminiFuWe1bP7WtSO8N61FthTxmBpAehrLY+p7xHv3v4zwZ5tQO/VkDIKLwrKPAjS
MJe9qjCknD4bUgMNGBx9WYAdErWY/Hb2ic7N7gdlHHR4tYTTc1Csrl3brr6AQWHiOxSnph1qZo3o
FEeCbTc7x1B+ti1dJhfhWhBEukrw/Pvh1Dk5k11PHXMSVjR/7GdXWMqeNJEMCPJHQX3+B/3A3Aib
Jqi//GgEeDuUci617an54CK+1hU/lFvTtmEKBQNdMeFhs+khVSjkKZJcj8QHCej0yZvgFgO3i0Xk
82I9zjY+NkkqAYlq7h4Uf4OrYTc0di4I+iRZB6m6L1KR6DPxBtbGDPFhsYkF8SL5RCxdlav/LoFe
YdSu9P6x5gbb1HgHiwRfkoidcrA+kVic8WS8ePZl+xEvYbcxG3B2Zau7MBqq/2CbGE20/cv0cGzZ
mLWR0Z7+gmt1WuAZVp5OSAJmAxWF9c0O9COfsl3kOaxHnnm7hrdJVqZoL6U/s7Qb5mVCxx4yT5Zx
En+FyTRAlDy0HtccT8+mcJW1giGaxwG4anTzwcCKlKeLY+1j5/g7NadYpA2JDPaM1HrpjHVfdW9I
NPEfm6HUG2c/4zlld25ZEd5y8d6Hnb1TUNSjn8FUVc92IbDF3KCvMS97gyXP31YPQ9/f3Y1u6qGH
ZubVJn/MjzeAD7I2OwOeZi7edTOjCHwWNgwRfa+hYXAKajTkTrNDGbttP77nETdrWKEG/1tn5Lf4
b8XWJFB6E+6wbKqkS4G0U7W0jr5caNaY+njZIxIglPkzuqtYM2lcBOH+ePpGvRRfPhLTMjJg1JrC
VGVseHe11RouvzY6Ee4JhodAvZj65BQM89dHZaAPkBPf2rgpLPqaqvhCTRPW9THBJLjYihBRZaWC
IO/cNgyg8HtkAfaANDY1UiRT72aYqEXekLzjVuSxqChlO43o0F1208HBrtTNl/a8zeUpvC5P/T7G
64zCYDDz+KNweVOg16U7vIGbApVWERDgDxqEnUMAI1TNSHyPRJ1HcgOMB6LU3PqXnAtlrpUZ9pLR
ds979cuDqRUdj0DQC+5mMNOJ0uiVTb5ukqHZQMQzTtio/Zny3uL+6Ad5stW2vNWSPMs98WYBSB6M
F3KiuBML6zaLzXXp79Zw8qT6Qeb1FnpmSm/+DVA9YFfPpecSXNmj1AafzpFhfj7VqxV7wMdvtX4x
QT3AIIHdivvaNMpzOugIVWRHkoIXN9SogcPzo/L7vmlCpouT00h/H4Z6ivd/FX3xszoZ2StUPf6H
qtrowpbWQwqRu+/Lt7hiqN+NfddIhs6M8r6hnNFo1gNIa40cN1e3EWtA/4Fr5K7cFRNaoSw+0bw5
wIWrVttBvbuODfn6pMRToHFC50SlkOeuPczYRbbOzPm7P7cRhgd+ZPozE24U5DW5jAym+PGkhz3q
YWmugSD9ahMPgNe6Nbzdh8R4coTbsJbUpH9cItQoe21v0TTm5GuTX21wBLn8HJPdz8dfL++oNcb2
270Zwg0MDUFJ6o+h/g1TY13aEySfDJL44P3EFveGN0hHZYknJKGqkC7+jgL3zX3Feqt/RacvZVm/
CY+Yoo+4ghtmuZL4eHWmEz/usxk4yEaVgLTSgfGcihrkC6xxugUW3BGnTEJrv0P/B2RbtpuL1THj
pzlN87fkyhFEmrqsjdfpXFW3cM3W961hBcTHAVcoioog+1tktO349eKM9JyiYm4gchCG/UlETsc1
9qz+XTQ8ykcLHgkcpaa6ku7C5C63Cy/Mc521zgDiNJk4NnrKmt7HZybxHbMutgKPachl5zjQQlMV
x/Hx3OJCbJciGqsGv3egPpmVQADNPP5LaNMVbSsarHmAaRbpPPTPdJfW+/YCNycsjG+bPqt1s8fI
TeQY50IZ1YvF7hJ8Q7OVRxQvCEakw0XwUoZBHmuef5nISZ4UISmuG6jJiDmCwW2PW55DOubrF1e/
GujTxi8N+7QQ0AZTIZ60iINwMQEkR9WegrRmvZ4/RoIgvc3lew/fl+DFAbcuFaDO7nZYk+s7YqbM
FY+B0J/tG3TH3wmz4lyzHXHCHXS7mU/7AwV2JhndBY9e2siiTHS+pEUR/uui5VcJkPoMSjmROydi
ynK6MQn50GDopNzjh9yYWALkytscLn+pVkAiMyyQcfzEa0/au8HxogmMw+EYDz6HZ7nFJxUjL96c
k8nTSt0L0dB+9NFOU/tjC9eCGGGtv612pDruzGrNAxPmckN+8ePrHVFw9nhWa3fNVbJ/9aE247Xn
CoxtgHvzIwyBcV2Xk1IfpjDI8fok/gAAEniUY9nOwMtvKZr3vLEOHli53TpJrDMW7Qpj39/WmSbF
pWur0KVQV1IkGMpu4sOuezBqadZ8CpbQHziXqOg73ADhgR8mCZIptb6rjQx23hMKLPDr8S8Xn3Db
rzHVhj1jWyB2RW5XoTuhl2H+LgZ2mw+P2W+z5kP7qqNg0S08E7POpWn61SLIbGrpc8Nth6Tr+rpJ
7zfOA7LF9d52sVXWRgdHrJnkqcKkVI6pn71HNrwvs2SLIIPAJCTgWoa/X8un3g5CIPrUxxnBGPt7
XtHMFLsWD2ziH8EiU8lpQb4tAXOJkIFEaaoTK+/uVLKM2mawpC7ixVyh8srwRi3BMDZbgOlmRN2b
rhVqXqR3+NKjg3P7SwBKTML9q94LGXgKjhzFBF+SweDWJZzzkCvv3gAflSMDf58bKGPmbyQrXtc4
eB5xfm2Jn1zchFyO1m5vBhexKt8ov1lUBsK+DpXCKJWPrd2e/l8/43Ybjl7Wz12x1+/5Rcl7m6IC
IMKKDwXqLYIK5Lj1lFgkdwIW9XYTk3Po7RG5y7DrFMIZx0iodNB039FfBpxQKVeo0OpWQbXxbweF
5omIkKcnviGMAmoHThx6P9raJojQoeZOLMwW9hQ2LaRon0ny+PMmDAdNP/Uh8EusEVmMgd+SpasD
mTy+F1be8cAwthT/N+n9BV+2/Zi/wY6RcRfrpA+f/0UuXhp4ylAd/UZT2uwwWf9txx+UDucL0bqa
ahCKQCMWKTaQrFjUxTr/Pl3guzE/kbTITVM6Ur3oO1w1U2hDiaaA/XQ/wbqE4hpebQPNRAUFkySF
8i97re9GPEv/doErTlSD4gLg4k3KnHEesul7qug28U1cHMdf7bT4tvJk4NmXTQRJjNbx7/01e/UY
V5jD4BWK5nxPY2THOroHOzY4qN/mMnh+K1Vd0aKT35xEpZp1gj9ElPmnNipBm2Mh+cQ9MIIFhv70
fkihwfVfueA5w5mqHGXmNgIFuu0mTqsfxhHJIKekpL9xTw/1zXPk2CEACxAzWbLSgoUT1kmH2/9o
WIZhah3D2vrHzlpY/q+Lz65/ysxUD4+evG65xyBy+WA8o5rq8dF4ZIB/7v2TPBbQTtM4d1nunk37
N3FrgkbHFU03m9ty6PRPcEF2uOZ6vywcfvhbg+ULi5iLL7xTGgPUK+lQ91GEcHd3AKYiGql85I4a
CkshZkutIqhPRndSOPGXdOt+AqMpQ1Sz/zWPEfMXoHBUGoIqUzwjyQHmprXcAlp6vZBfRNCwRKBw
nda/3g76cFln0vez9Tt5uktCVHrxAp0LEdNi8htgcCnXStsizRnZL7VXjUE/wB6CBe8CmkYrXYTH
l0h5qzi3CyXMhLxi0cPy28vMm6pPmAxP3l9LkHGLLiD9HZd49hF5xiQZqMoZVHonU023PCQCZkLL
odQg3WOMZxpjONEGoZhCegFhZQptgfJu+zS2JPdCwutHuJsHd8f92USgkTYqkr7bAR256WuWDp6p
ppCmJvDt5edAfkJGZ0oXS0gPj+5GlchYltiJSIomT7Mx6mToU8AoY3IPRK1IMzHZjr1uE90mm7lD
l+6ysG8D8TkvTkCZ4ELEib05YtQlAPjhyE0ZIVHGF3GP1lsgGfB3kXpT67vWQXfUn3tgaFFLtfPs
1lW2VDldRSVMlFt4VC+B1XJ9XSkZYfT/oEgLZc0MTbeV+oqCfEc4NVUwKQM6y9wa+Z7I1zQMqyV2
0Ninz15oyzGNNY/0ECpcIs4P7mHvIH4/hQ+Hwtts8XH0r6nXeov+9OH01LGpsFITGKKWSIqk37Q+
n0yDGqjuHHiih65gMtj6+4vP64MbKjNSI6jN99graNNtEGgksZxMMh6I+BB03aAJTv+dLQAMsqZX
EEyxwhSpNnJcJtSApdJ3w90YDF1UgZ2T7Rx1PKHjX3OE5kkvWL6NALzLQJISrQhrpvee/wcZX/ep
+teucxMbl6e8i/AGnQEbHr8gSszFKmGlWZoPNQPf/aUJq/gjNn+s3wfmyqStq3DnNsMJsuU2Cgkt
RrQrPdyNDW9m8gKE0onSDEAzy/hn8WFk8WSV4r0xN1ArvrzkgCEdBUu4iYDIsT3McecPDT63XJpS
YqRK4kmNQuUQIpGOdvDgrAOG+yVeF+5o/c03PlVTw0XVPoWeZHZZKzi5oXlumFBId3yNfnxTQdGv
zdNVP5WFSiv51/MhmqadaXgVkgmQkOzYlAHFdrlUdiLHEh2ilZlL6PCAbtleKpa/CziGeaLT6d8K
D8u6e77BoTZwaEPYj6tXqdKMA5C4qsuz7szGtZs/6xqqmck6wNFWhZ/0ImbZmOMG+j8E6/LD2enQ
ipYeBpYYGuieYaoCnt0JvQ9ffyDYr3JL4lv5AbOa3DDIyuY8YGFfLXsEGK1rywY371EibGH7dsgY
Sfg8/ic4JLYYjiNJVCoq/ytjnJckBZn6bB73+dp/Vr9T2GPdh0MBMSRg40ywrbVCIyKledZSsPEK
etV1zE843e36gmHgDZ9JHsf2WC5rLm+jVXTpIKmoGUO6PNeV9XJIbgaaA39bBbfV9qwvo/uU3DBe
2I4JOrcS74VGkGpsUa3FJB4X82759XUUL6fSV2+W4LxaHYkMQlUZLs83hfkKYkBnegOhsSpIX2hZ
0BKDDcfMlUUu0oxSFsMPgZqQmLPH4AKK6mf5JfMaR7CLM8q0lhaDz4DVYNX2FvqAhJU0fV7JWk9K
IRHJNip7d9yXhXl9CDBhv3PKplAMrbEwprQZbmAp+pk33dzQ5/r5Vjka2BzAfH8yFoKRVNYHPK+M
5rM+zIJey0SuWeVpwy1iL3NdeqEg8mEZAS/7FyNV/o7AxAx4vGW1ye2r/3UflPcB6R2uH6RfBfPl
1Tu1vXiAe7t2LctwotX/54ibDDWTkYMV/iv9LPt9erzMcphwgaK4JEXbuJNPVR5fOencW/5RmmgE
hJksLa6sHrmG9H8WjrQ6eApJHRScj987S2lGdCHnlj9xklP1XkULz+ix+iKSZVTthcJriM86h6Yk
j07phHpP/1LCbfBKcizgsw2bvgdJYu+quVoWnhB3udWZ293TKZLOYo9Ch7ia41fF7M6eWgDZ5hjZ
R/opSvmrXRXUtBqm1yB6BdchdaXyYJGrF+MpCUb+dMVDlt9v5W2Rh/pyCGzVpkljo6gZ07IwY1MB
gUp6B21yG3ZSuf2YzipYbMhoH4bIcWXvORE7hYHSzu9YFKfteAjL6Hiq80M4uQOud9I7LhwEKMrF
IKUIIAYY0OyjP79JnCxV0HMRzYTjyGKwRyJdwplRFq/qpaUPKMZ2Ace6XlfTvTs9vQE3GA7Xhiu0
e7OZFAI8L9LR8eB2IbyeF9qm5qydP5/vbm/832oMijw5qekoabQaq2701jMT4NWutd0W5t5L1dBL
fb+vPennkC84wHV26SMivDeAvdtpENKke13ek2xkIuYuqmLFlRuVOUCbGD6Q8JHrB94y3wHCCfB6
6CN1NNCTrgmUDLC5PfwW9HFyL1Ud9ud4n4xxo4goEtzUEukTCVCr4M9wgg4LQXwRIF1HnJWofGgO
rwEHN7CaDK5IZLJtVxNAcnl9q/hKBlbmo8NPVpHo/nczEE8lhm4+o4GSBzzk/Jbj14sBnMsb8aiF
bnUdRYQdwAHAqiTUbURhINxflf9tMqjnvo1TtcqZW5KMnYKIaBO4+hEg3wbHfnCGEqrpNfFE1tpD
2pSfRgWDrGWT1/FYSMYwX17yYLm3Kzu6PEKNOLWG67jnJcnMDqZHK0UQUyX0zPz0GQihrHZVd2l1
Aw9P2m+yzwmKdTVJItyqmy0fl2oMG7EazXsBy3jMzIU8AFabUm+kYpIz0ir08jWzQOS7VSXTKrmq
r1HXDbyDEAhy8Q2JPIj6RkHgBW8GKjE7Tn4SIj2zXBcgkd7/MRbpDi/RsCZpwW1mSCRZ0/I0ciu3
amUnN0VnWH54mMn/jXgml5LmK2uXC45RubMcI3ABdMmJFoblVG8B6BjkJ1D8QHfudWzpcqjiLhEO
RvFc+mfYay8WLCROecoNjlB3s6TCym/G0ywSyZ+x5/Bdw/fxGMEtjwArblfv6eLM6yAmo2nJ9Tip
y2U2IJKPM06vsCLFwR+o0wwzWkae/09/rT3aFvwVIcsWvbB20gVUodrBMwc2rbGnaw7EGqehdIkr
LHGWGJemyWm513qajb/r6/6QAl8NEzOTDJa4l85mVNEPQ+jNyb3BmHoRcgg3eo7mf7zG/bwCkOYc
Glz8Lr0scHtXYbYXKx96QxVDNnfNMB3IFTd8AQnxjpqO1qArJpYwk65toKcAic+OEye8sNzFNfMB
87inNWtlbQfnr9OYY6JpxEBnkExqJGr3JRuOHiszCd+fdyeLbsMNye2Nm5QEN2q7DPqd9mX09SFn
YUAxzrIuOWjkT5Bv0GAzhxvgjNmfmMO/1SAhsBoecIXaYwTxqg5hqMquEgEkeK8mypLh6CIERfoF
gWiHgGP0WXq/Lgw4E8kMXeUabP6CKaXuoj5z15HDRg0z0OURBgLs+AfOwK2xcV3g1QiirK3tnA/r
Rn+AnzyiVt9Yu3uyY/udU16/lWQqyFLUySMTW+KWGn/0d9QcSyEQ8HpTs0/eD+7Xh8e8i8JtxraP
y201fxfyg9DBTh3WeWVTBcskaqGTNodp+xQUapKDJyoymdKnFs4pgReCwreMtTfk7fJ1hXJzhvN6
a1r32g1fkTiRdREXYoosCRaYhzXkQrncP615jG5CkbGivEmZVrw1uKOfTegxtqft0qY5/qdIJi/S
mo2Srm6HFffKjeER/FrdApe9sada5VzLP5IcUTQURgl2Pg0dj2tpVdGcX3IWQwKXnE38gfh0zO9o
af5bZEidelXaHuQ0U2DYgtICdN4dR7AUZ0cVZByThjOs3DgcrugqdbB2jwR8vwh/k4mNJ+++fJBQ
UyewAT+R0hc0cPBQpqcRIrjIhc17qIZFc4eaImd4c9IJVmU1IWfRP/SvZhCkhQo7aamPLYMStGhA
8BHEYI5AHApOMf50MGv/JJ3eyx8bwqtYuTivIwsyI5VznFyJlqhH9178ARLqDQx+bPMz82MUSmG5
A+XWwABW6ejIvfkCck6l4UpD1UYIhmPt5kDg9xfbTTxZWeGHDKqvLlTTvCZqTo8u3ZbzxvGESSaf
daPvwBv2dfmxNERrMDKaBX2d/3Lzus9RmkZ75P7PlcCULUbsDggGqEd45QnHpAMxg86D1/2GnB8Q
oIjIPB5brZzc3J/iKN3kRqabEuN+ibVzyfj9nakYPk0i/G6kVCKwFxNB8kYft7hvmcWi3eBaN2+j
SF9ZsxRIM5TTv7/EH6iRmyhG0TnhwLsBE0fkmwxI5OS56IuEZFgBPcIAolaeAVjKVBGvaEmUF5Rj
oPHnzp1qTCoUSdmwEIqmN6KAlcUUkyECsfqhWede4uWqw2lwtSF6fu+T2RFp81u+ViXnN8uMugy/
pAHlQiDwWywo18P3Xvp/FiMvDDhXcKOPtOitUwVzzJDDx/2Pa69QoBP9Y3DUuB7MJ5evqp8DXyAL
0oUCM3ezzYgxHZ8O2JcsZI0LTvf0yKK10AiDZf2lNGb9fWRka4pRtLCnh23H/2hd7PoXVBO00lmN
rNSJvQ9CpwqzjjPnUxwLuzW20G9QLmdUy29CqSd5ajJzNDkvtNi+9TwFNL9pb8iCAqGVcHEW55dQ
QRIwV430SgeCIA/tSTgQAEiSUdGTEudQwAy4fPBMeGczye2cXZAEVWzhV7WwL5TcWB9bxMVGMEg9
F5SB0L4FUt/nvrMSZEwZsZWlTD9DY+g+P5/yRxU69D3ETSENZMUz4RWdKqukD09ZSr1M80EUef6i
hJv2d9vAWzaoWN32ie50T6sLsYWfBk30PcYglNiDVkY88ckJV3EdDSu7G+5mzgEOdGM9mvnrlT+D
mdfVDQL1wA1KO/PDEF3KuKMXIx2B9ttuld8pL32eS4mj7Kvu5lCZvLvxnpPZ6ebUQ+leEpHcWqtb
3c9Twzip5foZZlEYJYsUTXHl8fghWbI3dnuCBotpAVUgE71d/2THYXlJ0gu2gvga4TjhJfN/thC1
Q7yTJLiDwNZI+RhtyDsbCt+zQaWFc864rV5JPTAO7eYNc7u8lbkjgxwfC6z4w2pl73d3hYZyOsNE
zDskuKyRWVI7pMQPKiMSyi0716CTW4BN/18lTDeUfI5skIhACJOc76Xt8KjWEussHN+Fxzz8bCsB
8juTkcHwHhy7oG1Me2ZUrrOTmATiOwbBG2UKWt42UmNrnQc4h1KFNEkZ6cfgXKPAlpice4Zm5YOS
BQS26fvZycHPj3H0kdd5M/6Ac0J34me/tGblhmh7GPi5MHvFEa4vCo24054kSLPDRE+yLojlkiKq
2P4F3g/uSejhGJdYjxOPJUSsI4WEDs2oSYOTH58Y+dhOhw9lmCnrLzqK4a49GdIqoiRogGwEgZLo
AruK9bjxfMEy4Hx2GrF6APpe9npm3Smk0k4gy9VvCB51AvlKX8w9SgMEXCOd+1mBfLL4t87/m4f2
T3opGIlM9kGWq2t62Ys0TmB2cH4zSM0zXwTUc9uZVTrFY8vyb1/xrk1msyu2ovSofmMa7ei/xFij
yOZWSE7476Cgt6l290edWsuj+VbQDfZEVRfzBUCACJdoXpyAGKR0F4UUUsRC3a7Dw51hh89wPZ4v
PCt+PegA3knLvA1mkx1mhb1O8xrkDeu5Im4xKTFTt9Qdu5fLPVz/TPYOsm8usp5OUASLnVBodrl+
3AMKYVRQH/MTjhJIWaKbeMIGbo/PKAdXTasxKHy2w++6373f//pXVgxATXstiay65m25vl9e036f
2eKLSBQLXkJRGSPkPYTWTNAOPQVIIRV2ecgShcFzw4n2QfiBnxHRMbHdZji8aNpSHOOdXLU9po38
dEqEWpWWwkr2w8FAT3+iruHEzTqsQaG3+15/OdKXNRoTdnK0zYAJ4RH3vy78xdvxyzwRpfbZQZYJ
UX09tlEVcfu5fxuVRVVCogJ/byfldfFGjpTJaz1+5x5xafvHHIPBKY8j7xIH4QMIz9oTM51iXUrk
z3VAt3fsB2mWQ2M9wSGoLVnaXvTQD474KkE9ZHtrlqAOQyYhHEQg5lYG962qnGpfy3ydUQToUkRy
y2qZgSXq2yQjLSCvnbdM2Vp+e3ANuP62x7ZrT+SWGCWzJYU/HUVdiMm8b7y/a7swNJeGINP5Rw5a
qfWEhnQ6aeFAjbUCCCoseR7wNARlkCB9efvp/ZMGrzlH/V8S1+Zq8w2l/OWzHbeNEW1hyWGBNsZN
FOEcGJzZOnIhSbO1PGRxIjeUpMSslu82B+2Of+2fsSbFNG0HTPNNGDa72HUF1cmEOE9xmAc2Izto
mEndeGVcd+pmmwdK4eiRTjqyA8tvuYbSrIksYWOa+5n1IAkYJGw2iVNfrVEqRqM5flgxC+YWprUk
qRAuhAV6frKmBgzlLN68jEIEWWyhAyUhE4CdZc83b37EDWSRu7bTKgy6L9/kjhcu1CnvFIszynqD
oGQ32+Xt2qKMwei6qRX9UW1nd9D9+dPmQt4ne0RyJGs1Afzr9ZIhYlJI8FuolghxHaeHbaxddFD/
yyHq4V6bFe/478nTFujDrDtHHb6U5jrq/1Jxucilr5u7eQOs+hbhEcxppQPQ0uzEUZvzlPDLT2ez
wFV8VQz5kToCGr+fEztrg1JWp8bgw+YuIcmGuwxvLweqDcLC7S3Y3jhIY2Q091FvesrmOAPdoZEI
nDghJov8hBbC7ol7pBZkBimuGqxdUYpxy0H7KGCTC84EPUZT9eItcMWZpbetUcRguJHmiWSy4Akp
j+JjdXpHr+5Twle0UjoFzrmNNmQB0kteUEVA1HSrW7MrDYo6A/dMmGNP6zGLU6JrOJE1vksb5HZL
0U7UVowcQ0a03UVjfMCVNbzPIe8Am+8Tt/dyEnvxETZfUVaTTbD+h6CpWIOrZHLQChkhxQdrl2vf
xfQlX56FbjxP5f5pAr2ADlg3pDicxGGyaN/9d/92O1SQepDZxhSo+jFZViUNyQPsutwqZvzlcMOY
mYnIUsKVFP1Wp42iYQ3xTreZB/8y/wTqNXPp3RmEGpcQrcC61WuBVTFQtB4WSmBuSWMyLe8ldOIU
NuDwc8QE5IDTfJHmn1Nd0WJXGlnputkhF8TRguyaB6e3JItFscZoXZ5tUDcAgmLgZxSCOuDyx9W3
Ss+iiIyOnZqGU/9+rJUtd7m9vFuylaiugH9g8GzafrwdyFW7Sh7sS1+XErsxp1ZwqFCTDrFCWOdJ
8i4xuKy/+kUB+NeXDlLEaLm1+usFdVg+KnYBQGPBFTs88ParbfE4ykQc5P1Zk+rztCLg0www1I97
8C66ixEtT2ZQ+20DVe1W821dcasxEpCK07yCuVBUSjrA9kiaUQ58iLpidNU3OrmuzilKV/BcqWgh
by0s6cMzKLJ2xrPR2oN6y621UPkdS7uE6WPCHrB/tpeyWqBHfaFScAgosjlvdlEj6YHIglXEy682
NI8OKnwHezlmcObLVfL/R/xcSWctXCXWv63lIoAG58RaPPF+Iz4K6PV8A4QOXr0Gi+1X5SqUpUAQ
hxuEOzQBcqZvjZhctD6V9nV6Bw6Y3DmMuDQqJfKJJoIxOHzKxQaYmsu0C1RuNwEQtp5wCWJrSRRA
KazC6cKRt1ZDqoNGRpFC1qH4IhLrSx/Dfimq452E1FhnoOcQUhiusK3bOEfbeBAgrgXlNQRQPliI
q1V/kn6KEP2gTaU8YWrzNHTxPL+eGk+VsHgm23sVZtFx+PkQbSrua3DNweFvFwfqd3C3TD0KHzbi
W0026dRcSm3kZiNDj6tdEx/74+5XG7W7LtpZlT8dENM/0cBLi5NfrpKYJg9FZCOAJ+FXQ6zUOZ8M
kLs7fH+ImpQF+uuX1LiNDKPJ26agfzDuO75WaYjzT6nFZfPifBSkxwO6IYQs174rn3yrmWdSSw7K
gAerTfG6SqZxCjmSlJonwSrzaO2MZXfJREBFMcopIXKGgk75SmxaV1kNbxM7DN3pmg6YI/gNRUxw
gwOM9A4QY9qUlyvIIVvianOxuDRhF/5ydFZdKi2KlDW34X1vhL9xGU3JWWq4ahDMlmeR0i3bWWDz
F8AENG/BlxSAc8BAuOelvuVagVjgH6cvUDk4uhciqmMg8l+yc70QNfJj2q4E/k922CcXTnLMRP/k
WJsGm8jujfoxRgY+qYan7tyJZL4drqENYYL00QMXmo2mOmqPzhmHDbEy0831F2unjCklyh/xzmiy
1v0teCmd0qH+NvlZUrDMB9l0v7cwSr5UkgS6/jksBRKsqMP62RpfmrUQwZ9NMy5K56ycV73atqqZ
TkBlM9ilXbP/Zb8mZ89ZgS+4ZfWcmr461fyD8ZMc5KGwVQsk+rtB1WrSoKi/xaCUWNAmbaAr2qoE
6BoeIkCvfv+9T8E2HnqZdz6NYklyrZZQr+ZzYls1wqVOa55XVKl+OiJKbFjp3GojTY5NP9EI38n2
h8FWXf05NtlaRO7JdFbjjsx6u/wqUAnqlBavCxNIkruxm7fbm7/iP+iKCdBc5W5LPi3Rg9a2KO0w
XckKyrbfXV1IESYGAKyv1ryNbFn1X7x0sxRO0Ig7IV4UcT2nufZe094xR3NFs7b2fSdheCG7MUqU
TAefuOu+9HIWRXDRHbBvtwQctt2xAxxKOS2Mw9UjD2NJVOnaJIPFfYCRyGq/+bC0ug1tdu4m3jnT
YQkfAVE5lD8K9l70QVlE6fSgfeiE9coCJi2fl02ghwR9SPbLEuca2aifa+GgyxuLIpp58h3OTnzR
taWMn1QzwGptYLDF0btDIRW/cUJB4Uqjgr/Om+e6uUNIrU0fiwoTVoUc9QkRtdUAunJxN0xLxJH4
1SU1PoFWjZpKxy3dyu/i06dD6u+DTHRIRrNur5rRXmpalVTX+tAd0dRLpvrDr0HyfSNZ9LJc8lta
h7EQqf6mbemCHzCzFaVYBAaZxZDPIAk1V7YO6AEJ4rJHjeM3pIB31hPXpTk5Q/gpcxCtGf5eWzHH
+a4A9GXMkXXEIVImQEeyLm19ScxoXZD8cPcBWq/kb1G5wKSvoRDyf6YLdEQQxiaPu8LM63GzkLe0
J7fwNDk+TX8cgjnMuOQlL9PWipbwIGpE5VuQ5A6hZ31XKp/5NMp0oFze/32q8e2bo5ykBorVS6GV
f8LsExe6H3fDB8UIDx+90w7Q0LJ2OwLRM+vrwtTBcaHfkzBZ40UxJsnUb2kH/U8ItRCnn/jLAmuJ
kR5dzrc0RstDOIEFTtcsfQCxl1tKUBXBSHcEgS5MrkBJ5dlEq36TSy8Lh35hPW9XlqsJhx7Kv9j2
0SZzmacAE6gKdvPAiP+qdcqaVKJZrcWJdZOvqL6wlJM5MrzuIHwKIyf//GzbO3B314Z6CSKqyqLv
2Rwh0dkERZvKtEB1Zo9zl04lkZqZfFHiWn2o+09VN7foQA/XdBN67MwxjIBDMb8+uFPiuiHRfmac
Y2zYUR6cluc2rE6ffzt1W8WiYEl/fLD0etH+GwaVBCVSHYw0Whss5kBvZ1NVR/fSnbGdGvbRTUM3
8JcGYPMaszm1kbXuytm/vQipOsAz0zmoXnm3BMiR9W8NnXrznyaahJ8MGzSD1UqDJHqtPi5xVW9a
ssVVDlN3PHVhwxgzukdxpZDkqyrtvBOrX8Q9PAO4Qdvp0tOaGKq4xRa63EZAa+QHLRLqJXeAkQIn
cVLpkAdtalo5HYTsXzeA1bmsJrcGlHg7K2tTCqzN1GfwwrLiecdDUcAZDyHs9a7a58qY+Lnd+WZN
Hl4/5L+rzJb5jcZTgF/yBnS7H6tCRhvKaXM4mfycRP+I6CNPl23ysiiLZva3i9Bm48L8hOtWUehl
xbkavRbgfisQoX2rI+ImoI4Seb3VN7jA+BxsdOnCvH/XI6+jRXyPgm1dReiDDxcIGKixhQtSpa0Z
UBFQ2uB2l5eC3CMMXfjDURfYrKxmxwn6CEew4ajdbAitjqlW8tym7kdNu83Kz+cHq2Xlt8tZu0IB
hS0IH+4BYDQ0jR2/CDtPKh+cXRpD+D5ks1zwkh4eTHQi2+DpClmkpmUCa//iylkmK6i0Q+O6bfCb
bUkDX6bI2+Gxv4asZDfi0AD7EqZP2cx4Ph3eqO4/QZ4qPQiNebtmuMqPbec9t1doD30iKNCsU+dH
2BbfXHiNZTea7ukomuBI1+1ry0uN/XPPEY0gupliIpT4nXS5C5Ufu4e1c1nhLMdE2H9ltW/WXnbq
Fs2u++zEeH56nveQinXlF0vdO8dSraOlgMMjpamXH2TUiwqxquO747W7/MuG1mWYtw7693A6b3kQ
4jHyyCVzG1MzRUAPmE3pK+b4q17OTYLkRnxETVsj/ZqYtgTBwAbFchPQJDqVUuP9x+6WrMz4GeLo
u/68ku291/xdLt6yWOFjZPi2Cs1sfNAKo8Yy9fQsR2vDu7b8qpQNwnqHU9F1RD+XQKR6Xfdl1JaG
cUhtVYeQu9WW63Szmm61TRzMwkGzlkCgCminCBZLn9W1Wvci8S6cCzaOoLztwIsT+kKVa77z8Tlr
7Lns7fx3Ko34qrleJzeMSKpSAxeIRQeQ/mvGixCfA2fRakINupsoZB4p3XM0XuY2gGNzZdhlrzD4
uaEV1HNhJHzAqcQydaKM8O1HvrBW6oYnsGC3cTmbpBi+0r39jd2E5Wf5bfUjB44wTLR1qkUt8ci+
4+lYSzB7v1mdHMi8J/WyTGySUGsyDMasoLBZy3IFT7rSg3EX0RpZb2IB05jYumACvjp0eP5ll0Oy
osLmktxLh6WfeiFBbUVbYRUp+FWvqAHpEvHxzENPqPo5YiGBaOpkL4xOQWL4xXiyA4lOJB+bhXLt
V8o8xYoiIc+Ax3PozlwkTZlBlZ9wFOqur95V2aO8C0LLsp9NBOzwexRmmF3Cmb7OwUtLO1UMhivG
Xb7fyb2ZJt2nPR537K5SDy7pHVB/+EHrzaJb0sLE5keuMi+EUKOT7OHxnBWFDwq6x+zR8Tz+nflZ
2sg7kYGnNRP2J44+r1rIZ3DjcOK4NVFv1Xtoxlww3XUd6mx6qvsTBuvyrELxVPWScDYxtctHSxxq
jUBdAAmkowAENZQJ5Thhk0dZ/AMgn4cYu9TMn0KuBYd+UBOHglhGInN8iF/v+VTjhrSnmfZc3hnf
vIa1EoeighpDm2jLtN6/vwszhdVrtlTNB2Z7LL3V9MePYR+qv8Wsc2TPuThnoV7QgYE/4pgCIoPm
UZgTELzg41JNRJ7Bp+V+pGXGt0IBW4auQ/mYdzkRzu9Nd9ssXfSTNvO26YJw+MX8D4sBXmRgJYnJ
I7q/LgCd6FuksiPPlT5a9qAxdG3Bk0BBh5L/xDsRU1uvv91UM6A2nBWh9Swnt3AxU/4LEYZJo3eW
nre/g6Ucy0K6y3fD/skm/DSwQlbJuUB2TkhxJUh+8YJ56RtnQgrQW83y5QsARC4i0bE+7NGDYig3
DVEB1jgT0Y9PR/Ck+qV0R3Hit0KhlsxmcbBF+54EeslbB8olTUcDCbcDC1saATKcsWb/Igfe1qGG
fp+D5PPtQsBaFnMe/1hGZXgGDMUeNxf0sv5fTqvie4pZwbvKK/yyUzLYz8SfH3lEwPo2ZAlYA9r3
2p7hEjREH0F4JObGVPdZBdkMgo63BzEiV1LkPFfHbxN7E54fPUs1oZQMqRlvY+sAoEIl6t2+Fpj9
K6ZbDd1mRdP+jLXhSpdb8+hEKweG2f6sZsPNmFmU5m5GCDwyyJOlCUX3dM0mODvyZpc2IzDmhaEY
0ZnaWVMmKWjuzaP74iNEJ7pKn0o/E5EYm6uulI/VmtEwrOECvi5Tv+QXYGnKR+vO24TXC/ql62dV
uVb9waMeyrULaglPlWOw8OlMKR0nFizjpNKevZyCh0ymfgSKbOQ6Hum4c55I9kw5Y4Fy3GaMcYCQ
Pqi3VlWlrC+nB93+gEunT2UaKWMx3njl8pBq16SsbiuJvO3IDlRRTbjyYQu21BNUPBsnXzy3O8TE
VA/YoiDvmcMca1HnzhjR92Z2VwdpzN7lzEH2XLVT6o26Czzeh7noIbfCa43jBlYEgIbvkEPCkioL
HGBD3w72UrN/7IOSb7Mg9zefWAaSeIeVU7T6I9G2+d+uvhhjCZdQjgL8jqvA4DeqIm4lrZ4yQKkm
2qPIQhRMb6UEtaN+kl0ncoVYilDtjscqYxLzL4A7/9blORzOsvIHn6mKuYEnAsyZwAcQhw6SkRTF
IX4VeEX14ZuwthjvW3g448DJwwQSE9If5qhi4+16RA5yJk6LMumRbJmXlYc73OOBG2XkIJtRdAjZ
4Ori5aOBr0Yan+eLxgCTO2dEZ51tiF5T+u58zRyuo8BLD/dv58NlTdQLlw6Nh/Gju+vU0k+SO8Qq
me9f7daqvAzjTYyrBaQrHvTHy/kBs2JSq37oWSqBrcPF3Tp59z1EG9X5hU/qaCuEZhvGJvicmHOk
jzpwQEg/rk1LFdQF2XaXtam58VGDlwOcG2uFk+I2yIHF6SOrYcxFcRKDdwY9u8ZxcCSrE2fCS7Lj
dStQseMt7Evfya9Jo/7/s/ACAlg4YELDoU2wLJx42D2MGUxNKG6DQJYrzTzS2y491pQgh7JVVsAm
2F3W1G+/OyhX4KAmuA8C4DoTaPKaCU5vr1gSgNaNwcPXlBfe2ECMUVvF/GZ0V+nxp8M3GHLPFoxt
KxRTmwTdUL299Ov0zd2XWWpLx1Gs6gyU/24xCbfUk7VDInJSsubrX5Vg6iRijaSAE8aypj+CsG5u
XskR0QQxgNlqXn7N2krY1dIonEDu5bav0Bsr/Yy8f6mUbI0k6Nwvxc82/qisWWnni9fHMDzcXKyL
8MpHxEaOuOh4YDu93+X2Ncg0XE63v4Pj1derJGF9hG9zuK6EitHYqc5Ms+uFQllyB21brKSKilLP
MXS3RsVu6EkoLsesZtbPBzOkr1db9ci4nppalEBYI8evT2Bu+WiZgZTC7822HmZOJD6T3PyWdDVu
KkJEwgZ62nRoWlditcqUGKdsH7lSUPEsJpiaRftE+AnwXvxJmaRGYXzGJ3ukDf+Nl6uC4XHdzjgB
kNNZGw4bbY12l030/6WhmGQGdNOxOb589KUfg6goXynjO8Co/6PXuP3mqa1G0zJbm2rX7jTdxtcI
Ir2SPBo5stFLOnx7tZOOvLFFM6Pkv+VToarfvCiAkTef2XwUJUyDIKemDJqUYGKvicD5uapvfl6K
i1L90QkYmb42aCtNA+UUo6qH6dVDwi7KESc2rhrHvPFwsbTjlgIqhbN+6Zz4kuJQXcMoXSQ9/ocW
U7yAZPznSvNLuqdaWv+q8MKLnWIzg+NPseewhaueFpbPaLx350u45wowwsUX+J2rUv4UwJ65Z5rS
ACOBr66MoBLbbNg3O6m2a96nKuvdp+GhMWJu4omhcIyuNIfuPOZxRN0iqGY6r72D2oBr5zUIgodQ
W7Or+t2UGCYMCHr6a65NjtOxgwWUQ/m03d/qq/LT9/HgvLcJB3KsWP2tqQXjtCSVRDJxKpPD/K3l
Uxq0WKBjU5c1Kk7JOmdm7/i6nmXmvHph/EvxbFjghIIhymmmSWRJDAMnNC16yNs7fzzRSvUwrmKj
EWb7H5Z2nSXr3paZ0wigGdcEjEvDDExav7bETQpHq0Riw5KNAXhdbqTSTgLd9dMTm323O1sV/q8X
DEMPfsvLDBTigF61L/PiCFzyoZPOS6t3cCpA/Ax/RriNHyDkXuex1iW8ZUvhhbUCNMe8mLVj2glE
GDOcem/QZMIVZuNXN3MsOHiQdJss+n5JP+DbqOiUCeaGOXgxd3NseDK4mOidVOK12LlxnZikMFCJ
TwSdPJKFra+/svdJb3MgxhwZtam9rMOHQFG9udo6Ms+mvkAYQsjlqjhq7iI3eJIGdD6Qn7yFq8se
nmC8vdmhP3ZTJwYk+V9ZMkjGoFzLSvcep54w0qkT+JgQB+dlta4Yo74rONx3MjD6iDxXPijmUeDS
LsQs4IvpbPtmQzB1EVktthY3jTs9gmQrawd1s2J/0EKj/77I3Zsth3eP5v+9tZVPXK9sQclC+aW8
/+NvvVclzXiWtpsgK8juU7BT1NM50jRQkjoJM3PE1w2cJEUYHJE4VRMRm9S9v5HS7jTGW2lsE8oS
frwXrrO3vgUOsIsGvmBpTRJ62TQeUz1zwo/ANLit9c5IUjxHi9zW5gbLYPbcOX35tAffVC1VS1i/
wQt9ZBJ0g0qOEL1zn5/oKGwTnbTVyDNta+F6mvVFnfPhAlm5OfnqzkjP9i9r9iiizwhEr81AEJlf
G79nfLZVSPu5jduqjTmOKrpsfRFmbfNqpmoxjdUrkX+ueTCeBrHK9KCHwYUbCq2sFahpur2HkwpI
UwSGRvRNJhUwknakNoSRTTFZ1bDtcWSOy79vYXZ59yq5tABQmraWX8fc43JUB+/Vb3urjM016GTe
pqNbOkqwiTKA5wNdNsgPbvEsCCvji1I/S3p9/lldkQ9IitrJnNxCstVikoZ4t4z5Cdcm35v2sHeq
0lJoc72jH5iBV+O+2TJde7vORVdRFUwVJAALKVgiIDKE+4QDvcZS66X1oKhHrvUa8aVpdeH4s80V
Dzj+pDWtkdt31AbE152jS3HCoJqvzq+zQDfxA2PrDA9cz+mV3popNXO5jtNS/NaH/pimMiW28RFx
owZG4kdzI4/TW0T+GKUqKxdstnuENB31vSPBwfIkyafpTB3ZncpRUtAeaewmdtntPecQAuxCXcsM
LEEw/NF/7AWMzPMdTsU9SfdNF21DGu5k97ViqYvACQByKO5EjlDQTHMkzxqyJO4Hyisv2iHKbxOY
u6IvOw+7wFD5md64etA0+p6RPO55Ds7rMsWPl1kuHvdSNK7Z86nOPRMtftOE7PgXuiGeBjsROR4s
4+W1mNE6jmkrUFtY3T/TqqmF3F3NKZXKtnazqmUEVWm3RUJJUu8LW0pkHd+1ce78umeIJxZVGT7i
aq4id1AUBDNl3aBOs/W0fomzpBszTr1x4VGId4prdfAgUGotO76qQu5Q4bnzoirQPQJ/7tBvE3Ga
8hqzB3XN8wettEBg1R/7Jcrb/jBKyD5Z9XeKgpNZbvePQU+KWInek7w/taHIVBmG2CRsmqWCW21y
9qGL47FqT8cqNqqN86xtCsglsUTYk2h2kr8cV6p8U6RnuCjQ1c100I8XScL7rx+SAOzATL95aDj0
WEbX9X4EJgVdc9eJkOUAd9jrYFk9NxpyofQ9hdx6P1lJ99FjvtwYcz2EMYMBDGJV0Yuzfdaa854R
0YkuuQt/QtPSTilNlSyRh5SeAXGHoW1T+Cfs6A369L53B+vLskqTcwx1HcgrWCelVkPrZp+h0+5H
iLQzLcxAfdvgVeoZJitA+JRsqsoZfnjoHJd3s1rY3QVCrH9PuwlZoxqG5QBi4pML9G7vahvyw7Mu
VQmwdin3Bqw9dl8cR4+c/3c0weuA7vDxKEC/HtNKyJRPwkq/QgDKtNU8owLoFUNQ/f8B7iI0HCZT
ef0SasUbyD6q3gNu/0bagafob/5BOFpUS5PHdp0we7WI+YN5x3f+Sblb8LTIPSI48JBmizsAg4sV
hPfFpS8T2XoewSb+z0qXWH0XA0s9S749AWjfl5OOqLwFcsnlqgSUobjbuHiZZNiq4yBx2dXau0wC
voPI681SmwV+8xb9xaYZ61SjZg+GW2D3RKOB6ohSQ0aNNhs3Yt7W0zXWTg5ZvM5G5fUflDMqcKpF
zDjeFbZOqo1Bw2QCbTgVDsXmpvDF5VFv+0YZlLQMzJkN/qhgHrp7yRw3NT7LROkIOF5vDNd6TT6g
GtDAhrkf8s7vYcwgtT292TQodW5dr2mewMXIG4SFhyxZpexcoHDMgsj1MEvviAjj72A6KErx/8GO
bwHqLcrDffrHvUA+pzB0ebVxbiKtAv0JkUSCCPy8CoN1VZmFhm99bABT7w82JiWp6kSpIDHT0oJo
RJ+EO28kCTJDlTWmzKiM4w+/OT8shO9IkIE9Q8AfgmQdbcEXhtKlsHww5XkQB8IA+GY10A7ey2qt
5E2sco/8ahzAu7l+Z2i6Fr76DBoS98lpGcbAv6locyUq2ftTiS8flwLhkvQKEZIb1Ij2SVz/qdQq
1fqh2hXM8L+PYYSihEG12d2pgxw1QmObmfdZ56o5MlKcZR4i5D10/HMNLsMUXXgMUwpwgxwajl9k
UlJOB7Pyezb3NO0+S3jen9qAeRQZReALU2x7o2cmGkKdyoxa9UVy458Zf88RTqtW6ayDbcS9Xn6J
HXjiRbIyi+OR+3VlrapyfjJsCe00OqsBYxVtqHgSDdNVIbAHfUgyPhT5y+GEu+SvdiN2vb93VYdT
Nb5HrOhbp0Kf3YvczWgP1vLGylrw75cdi60ERc/avD1aHQ+QjCYhDNgupFcFovw382U900pgISU0
RcES7A6oxJgDJQhFVIH+2N3ZxrTAKlcsu/y9MYco3/DyoCdRXsGD9lAIA0qU19ugwhzybTGBwx+x
muI+a71DWIRBzKaaDOkwrDbxsXGFVvQjVRxxYerAgLKldFQmu9uuQ1AOywHzymZDgbt6h8gBj5uR
rJ5GSJAwVLCb/8AJtSI80pnOrexk8oI/0IJYuEgm9ZPUD+A0/xn3Z6290SmWKZrkwFDc6zNTdRhF
zgZpNdpo+kyCS2Ktcd7bv9MT+JX0R84i7OGhCkpoGvvhih+4pZ6dXuHLbaLsRMaDw5s+ydlK/bP8
R91HQXW3HhVK+Oa8gbePK0XajpcCHw6GM77GkB14HT2vdencIPaYM+xn9gWPAKlCzryIFmc90gUn
hBaqSM6a+HdNvhrRlvBj+NRUN74FrEkDjpkcA4n0ut75Bp6Gii1GDWjUPYM1A3fJU0szEPOK8z7/
2vLVic4bi6H0pEPGYot/ZvaFHEPU4h9aRO1MuL2vS2yTvCCOzVCajV61uPRn6uzpnsaVXUbZcGZ3
ZXXmOtWnYUdoVH5CUr6VBiYoi/KvIHVJxsS0l3I8Vy9fzAWtHK9gH5NtkCa2VPeqcDo5IJw83yHa
nYng2qKm4tn0J9igRF3Xw3dOP0gIMPptAnkNROIcrDhxJHeMNlfWLqUw00kUXrGwyQxgndQZYaaF
a9rFzHAY/MosblqunhA+mLplofSHaFY8ciVnq0SQUj5ycHE/9pFpORRv/2d6XckRYyLeByq4cdgU
HZ4rfv9f2wxfvq8kmr3QNEqe75MDyzl+Q3lqWiOFRImVL1e5vV3J3Fnul9OJEbqLu0eNDK2BeMun
PFLUzITvSVm8t8AnHl/IsfMkVbNfNbKtp3fl0WH/JT+tQAgBLfjMNRex9+hio3N4r13XVUZ1nBPl
0ZpCObI7BHgaQZwte4jOvpBJSylG31DhJVTCmu4NrU85TBReTVAGkRU1IcX+XI+bH69x+wcP6TB0
6lyNPoJTzb3VE2KIKU7/RdsErYitlHU+n2Pm4o840mZvbeff8SLJwj7tlJNuRjeRZG/pu0kiIu/f
O4Pi/EVdQo9Kx8lTYfgDXxTn7ot1QebUWitOic9pctgm7U6i/pIDfZugRtcrroRoW1cotKpnrybS
5cYaU9G5omLadXValp9k5/05cPrqTQs02Utk+OtDAkoMH2DJ1hVjTwO8gzAKPErrV5TGmI5JsH6i
SskZTqQL8RzGWGAZkrHjZivz/TF518QBpS3dEeKz0RrvfNhqKCBEg52dlOOx0mF6CoFsw1m4yl0S
c2OS0j9YhPRo9IroB+0Qe3Dw1t38+K9kErL3tUhik1dCszxRAUcsnOqo3LeUlbupOxaFqxOd0hoj
Hb6igQnk2dpFbWcnaimpFkqK0ZbFTwIIxs9sBx6bwd2ctEAMDRBs4qSJly+Y5kh/JrRdcbNptZSZ
xuzXgWBAgHW4BMOq3yktB41OJ3QY+2i/VNqbrKA5bVivN2SmaJqZUplvXI7xBvwFcmWS3oBhODUP
11RcQdJQPwESe0axSiXqzJqaJzxmuk61xI7ls0FhER1XDs7TuG3IzrvMX9XTTbRhX0FxhrZp2fw2
AttAzm347Hi4xuNIprdVBnJW92CNvWCpVsNRt/JyodEe0+FPSTbH3WU3qHbKPpOJbD8cwkvcVz4l
V195WKkUxiPlWZwwxXbaAAQWNo+B53IcDZ/kyYLRAWO08KzrHEjhm6MNSZo8PuoqpdZnOnvVbU3o
Z4zRdWnwdpngLRrhgIKVzU4MdMHIdm8P7stOqEW4pLThCZFTVm/bjjW+5OzorsWZ9j45mDCLMwUl
y+it8WyRYRxqO3x19c8noRakQypMBZriSvAMlCSv2MhgihMnqBsCGhK/QZWJSzmkZ8EmPojsi3Am
VdBobYZWjeU7BX7sWCq6C3b3LZ8Oqk4iraVtib/llgqFKbdJLt+Gkg0FIEABHD5KMEibtREMPDtl
1ZmF6JjNUJGCl9vv2UWhsa29JkLodd/PWZbGwolCa3t+LNlvwc1OocLZq/VXvpjaztzuSYESORPY
LwcVdGVXLy78tUGto5A+DfO+yrUA4wY4CLYyGH843HU9o3s8i9K3f7HXpGSu0lKPaOkVWeRlXdwZ
CvfJjLeLdiEWbwTW/AO0uwQYS99RSTzOw7ZUpAiGToLNFB1n0ZRt1OCTulKsC23ypYS60oKNYaqO
r5FvC4zTeNE+tWs3HWE4H7fb6QkvQxa4W1scKw8wEahw9F0kcC+Zu/OEALP6GA6Hm5pMpWh36I3G
0PnleWvHwNqPIGkarLlLA+4eKRq6qEPGQs6wqJgJloAcjOTiK96RbUEe0l6sq1LiqulUf88XjWPd
nI3C6LIc5gtE43qYkIMcmhVA4bgroFhHfAM/2FOEOQPVvfbH6uqv6SjxMPYYfBZYdlyLIp5WR18S
6jQFL0t4tqqRlkyszARQGCOuh2ZiF3Btq01cBO7n1q7GcYxwhCsULsMUIBUqA3VEPolE1slLiOa4
uKTZOtOtzR1GFS+88svKdPckeK0OpMS7HPumFxGQQe1m2YBy4lUfUKoF0DVo/EKllXgM4YcBkjjz
K6MUokLNBXUa5kh8RAtj/4/FDtlKZYdR+hT7QKNzMy3SUpnV3INRITXolyFHCzesVI+67V5+lb3d
E+flhGyoRpCeCHqCPFT99SJ2LO1Py/ya0PMv4caNmFFLqnqJf2zaCh1gwzR5tFiwuWn3VfTqKzkw
obquQzBchWAUWdqX/Vtxy09dZadZnxWfLp4hYLuG/9vknohZYA4AL3aXZM3K5QeEEQZFGyOOiAro
wS1x3n5FDSNJSNiJOE03kZ46P1ZQ9XcfKKAF3ak8gzgpOvvDEKtpQiAFGRioIJpfusBgqRYr4NAT
OoLysSPGFo2HUGcv8ZOdl+cN+8NUtdfyVWzbhutdwwjNUMDjJOelqQdxON7tLHN4LjDFfjtba8W6
pLJOANiDBSE3sbfCOxFwS/VVcZWqFAvpMWGafKyuptLCdBPU7Ssaea/42NakFQDIuC+Gp4LwGdDi
gfq68PGTEFVSwfIO0Xcws3NEZ6OocJysD4eS5T7r3JWef1vTG+oIV7UDlBj7xqUNOfmV8OfKP9zQ
xARcFAdmCnhB+gUrcaO6JagNZAKr1+7AcGUvwTNZ+VgSjwoFnvgfnl1JCS10j4O6p0p9EEjliL8E
Tt8+qG+6WqTtbSoYkU/lIerNAY00E08N/TQgDH3xSv67S8NKDU30JvcSDeZpX9JmwJ6S4zkfqxfm
mC9+acAEEqwAI+NTTvvD9TP95XUPK7+Dv+jqLYnMD19VUIubio/z5oxlMbofR9kiyf2eW/q/IHXE
yhB8ERaI6+xm+HhRKtp2IAZzRhzba3KO93ga1N+mq9JDWqsEO9ElcPIL3QSb+H6J9SONbQUt8Jx/
7+Gtzj310qtBXmhTgNFky9spx7bp6gU9JsBzG31oAyyA17oiyej72lCj11dt4MrVzO7Luk8PMVT5
/UtE46uu/HCvtDTgIk2eVumsSamzZcnMKocNvjHabHJtQ5ik5teXf4Z0VxIBs6OlPWaMolLwOV+P
z3iODVcenyMGs2Dq33Wb4295wmxlTrEgSh6gevcNHZfPT71gZbtYF/Bc6dxzxaiIq0hrJOXOOERX
ZTJIWYPCCkNh8igWqiwON5xpZ0MM2bWbH5gxbaGzVWj9ypiiRZ6S0Hc9NtfCucPWQqWaFuT9kYjL
wJHoUpp05zdKo3ztGm6JDRlbJbo6Q9ye4WYveC+SLlQq9ydxdHyvkHu5jy+eEe2AhvKQZTBqNz//
+b/6n38pM0uAWRQFuWMYGEBaw82TtXzH5OrCYGHthti0lRf2rNT28+fjwqGzrD9vhnaZbRG1KHDX
NCCmmjG4p8wQ2dCbDL0BbPgiRWWVluubPLBnN4BrrEI2YQmo2+Nrvi7plEjtJV9kMd2XZO+rujYW
w8b13cpt6GUTKlcxdKgDVFsct9p6TLq6KYCIs9puSbFaRDbLDQX6syBjjmv4QP2SNv+fhxpHYatI
O07UaPY7WI8lQoTjRlU9gOZVoH8BbqKu9xFxN59m04OHdiBkYhB+ocdDH+diTxGjRZjR6U7Bn29U
NsqcSVEM1Hle5dRCSTQl3OEJAqj7QylWwC0DSLBoZOGjlG/ZfZjol5cn78MHuOzTZhTb3wdyE4q6
HNGW8iciJkmvbUPNVDLTu5HCSGCc5KFD87JbyGAbFZMpRZmtcU844oIYx64dj68A+wGVVRY/zcSf
x/JrsfOTvOrLIfgg6CMC5SyxUWo4woyPpQmsFj4Fui4eIKksOl0hEDC/awhBlmRh+wcuRRASoG7B
0Xlea5fRycc+fL0yiX56T0Mdo5uVfhwV4DdTpA4+CD8ZjzjOem9ZI8dTsnoPCRL25iNVgZm7nCj6
a/4VpVNmWcplLM6Dm6bM3gK4TcUlcBfow8PgeGJ/k6i9H568sROcCnAFndSYzxcLrG4OIxtyh40K
hC5pIVvi3Ip/4PdKut3UMiHZd/AH+4OUTv/6FNIG/sYK0BhgZhirfxTRbf6AeUpUIRGVRBUjQOpC
fX0i1S6XdxqnFxWBn6kqgilBiPdYa/RY/CXh1TlUUwHcqHIzXPTN9TQvd1q1l38L7nGbjZFOMRdK
GmAKsCzkgU1SZGsrfMLtroNclYEV1iI559VSuYvxitmv6InnHu4WTIAy3ao6FxuVynVHNj4RAMC6
hcAuxrlt3HyBVI7ta++9HAZNkT2CwYRiZ/6WhY20IOtBOzR5YeyK5iRMnANS8PxpxzOFKrQARv6O
jRiP+Ug+XZf1GIPwcT4YVmoauiJOXLGTD4zjMKm8e6cUahSjtZ982M6Nx2yb4+l0HviugnNQrxg5
EKw5KfAzSMHp/tdbarO/HjH1nXlKsfJlYK/yO7rYIz5x6Fiyq9u9iMV8AEjOGjwOTQIyn1OYebLw
RJBCDLPDLrtUKYoBkt1o96pGKIFn3dBU9s+4eOrZf3MLUAEIuLKR/T+cONVWrxYiJewJWLsHt2sx
g/NKIPgFEL18fQr0HkJPhDeiNH+S7uF5PZKctBdgGXwBvO4PfTUXa9peCEv4qtUwgkYyvb0blo4S
C9W2awfWTOPYyfF3PuMRpbAAbSiiCgOXzV38La9sXpyjXVaem9LD55FK7ovi9g+9d0ae4UWAyIMA
Ve961VBhMbS35WJXWFMy7utz/VmNWLABpDlEyLQI0yKM3LTLfOPypHIat+hNYbVZBhmT0DbiKBzh
/R6ddAlZDuK3NoFYjCqj/WoFLQdhdTXoAd/lVGlUqDHAdWdROAITNEuNb1i+986HECAX2gPanKSk
ijrnIuHZyUgTQEfaUJt9RzDyVV1yAzCgcAsJlWAQWrujgHDx/ROGJZoLEINuXCiidHGJ2Rq62vES
hTQzN0LVAVueTFEqsSLrvtP9i1Exi2VCD3p17QIgC4ZWLBf5d3rHLekC36vrvKjnCB6soCE38IlH
9tAQYrRCHZR1rblx1DBIjUIKSX47BKKBTPRnzwyb4MQHxf03gwLOn+403LhBLExxMO0bryLPCQnf
E/e7rksTrgshcNTyjaEuG7v1wwKWy46BlXLqV8t1ELBzWc1MsGNJ+kqTLQ2hKFem02wJXm3h8qdY
8dDq3ZcoyqYw/uqjv8V1iVFmPdoGU/dMPkUwxNZDn96i5aHCrfBD/DiuZ4pc69KtJBMJ6s6+UZ26
Vr1TdeODJmENHzKKoMGITpgg075YZU1yR5/kljW3XAi4okRxYOYKnQgUYx3X3MWjMHl++vVujtkm
k9evut5/cy7KutbQd4XCib5MtQdlJbuSINtjzk4gwvcUlvHZf33UnrjG7cJ43yLmPuiiO2X/rvJl
0e9d8yOLTmInmtXz71hIAgBnp8E58koaxYe/3X0zbxDajp754jDefQarYXhNR6wmaH9g1Ge3+Tji
H8LxlUNc2+oOLkTqOPWZvUc+tE5s9VLbk7KQDTdz3JhvzsaJxf2v85MpQXNGI/mhw2Z/KVGeat20
JstcceoZQYNih7PxgQUEfjzDG+fK2zqIqAQgCjizQbi3gdSALrN1ku1alEo2sJX+woi2GE2+Qfcb
mYgw8Ltu35S36Kvsrdrlu/e/cOIZepfV2AJAG6Fv1nbD0j3KkD9fUZb2f5bf6NvPB4lffKoqLziL
6Sn7mIpN/1NzoG7l1Vzuxp4EQ9QGIDlqnNXFSLK2YG7njmWvBtXb3uMKI22ID1pS6qrs4rIG7wPl
Tj6pddo0BX2IHOs6KQ19HEEs7eh59N0vzmxO/d7sJfFruim6VVj12Yev4RKdtDwMU3peunEESLEG
m898eLyt6FDghfaPW+cOu+tA4Ss5JInhc5cnR1Ubxp3Mg/SkcmOUBZxXrNIuY4LZsDQnZVfbGde6
gnxVw+j0ap+ZKGGGQ4JAVm7mo6eN9FkU4bOlNAPazz9FIZu4JCv3xGoDrOTQv8fxKLLmSimV7V/o
I/JHscvYTf41YA2JOToN2V9ALSUdFBIsPi3DsXS854/tQi14iUMSqNyqe7omI9X6JJewJf5gQT4X
HocBrnI/212ByLlvg3XlqoOjr2wmXAhOJZipg+Xb9BpAflbTBJlr5jq+fkQV4KLEO3YzAQAOUgLm
ELN0mJVvhqKo84RGbzKPT/IpDkjxibGzAZd1T6HJm7b5n5764hIs/nphumrB4/ZIh/TIAQU12GJw
u7ddU7I4EDPBPrqUVVa7Y3xrNwU9UlT0OVzu4XJgzmUOaiOK/SKumTBdF09rQkA9kqNcexOaHJhR
SWcvFFzTtpM0I5Nb+oCk3isQOLzkONOMJjghnGGjDSmMm2ogtOSYrnjT6RIPY3AWgM5M70m7jeXm
PDKzQIKyOg7Gv7fsMtoq4lOMgMb40n3tj/SNLo4cuVM85ZwJ8fl/vm4lfEvqeMISbMuJSA4+ATGL
+eeUJaOs9njfR+c9IFUjYKCvVQgo99RLh3eUXkLZ9nDdWdpBSlBBJdifqPYzwtq4Y8SOgUijFbp9
6DoQDmvtnDK4ZQKRX2tihC6L3D5noAAP0HPk1/4AqKkp91ZpC4y6Kg0Gv8qkEmdYz6MH5MaGdDD4
zWWoTCF77s9UF7ypy6CkYrwXiBlNX+lAUGMqhqD1mneNhLV/o1Y4fY9qoTYWYc39T0Bbkai/vuQI
l4nFxsxvS+dGp5WJvJv9yXPX+1uf+HKz/xuSvIFzdCTqyvYnfcS+aX2ZyUvqYKjt9N84kOG8kS5y
Wt1e7IASo56hK+6w6vYHUo9f60zZ+Mk9Un49CqUTqy7lMz0mUZAZDo3NGCnuvIh+ytxkAtQw9UBp
sHTKcWkACQiT7yKuL5PfSFNehfxTzD71WfBSLzfcb0eOaa4hyPuA0FSouBgFHuku55YO6aKM+mI3
fmiRN9gBYVcLNhjlfod3dZhH+DaCteuAnfU8fwbw48zxvNRZE99OX419oF60CHzBfOOTcOtMcBXa
1KEqsjOrACkOjSL0mVt1FPyUQUkMX/oAXEzwUKXNRfjg93mD9mA6ENNxPFYmteMRdnVR7fI6ZIE+
sXHIcQ9Y4izUosjizztzcwhcJ9vVW/Quczcn2F6/voI4dxQTuGFZj+j32WT2OTlGKPqYt7Atz0on
T/9Xj6MvUmQxnBYjZ42FjWJoLkKz/Mo4EDWwGdD52Hp3SPYpWI/mkj/agAGryNWer+pU5592ZgKL
5Ey+npsKmlm0F8HKLBFtoqPv6mubJ84oL4X3yR3WDi1cdCfJMyogSgQjM/SjmWOBdsvLv2Ekid+f
Yg8Z2ehmcmR9PIVcpQdMERLe/+KZJQB/RGCUmdqK0Vglc7IxHM+7zkK+RdL0vwvDCamNWqwXNl3q
+EGSglkcIhi9Lzm13lnRBJyop8/nctE076MlO5vlwn9r/0GL2VD6BEiCfdDINGJsr+MHF/Kejq/L
thi1GzbZ8qWbDoeUSCXy7CXUd0S3U0JoQk6Ffy/ZlT0wUPvw8OVvpVoqjce9mh09xeHbyYBJXp28
im97Sll12MiVcp9pNZM0C8VvXF3j2RfbM1BRCv8EgBLGIgz3thzfFvCrt50UjUYadHsB38vN62DJ
1kH8SOv002wCpDCDI/vRTehV95cEqpPkJRL+wVP/zZvQrKg0fuHg80+XVl/WfPdkOsxdkzTdaRPI
XwNy28qXMrVjGXunQMask1bjWZHt54G96SBa5idDItOEKPw+DpLCDnNhLu2ng2x1aepN+RK08CX6
BJaqPv7XZpZk/Iwai932H0VmHMkSNnmFH9/ovaXqeP1vbVBjBlMakWAQ00xs3G6n/itUWpTdCkLO
D9IYIWnvnEQEgx9YETaY0UqoUECMT0keQ95zX9yk8MaEqC4BOJ5c1/dDCkf5WZCKjw7qoSvdKSGX
zGL0R5lKXjuMAi/ke+TgqP7DTg7OAGTbmm7iU9M7tOuFgO8zjpidjkh/A6wfchqSUH9dD+tSgVWM
dkXB6K9Sm5OH0xw7sbyJaqs5A5b3poxpAID0cboxZZ6PE/Lfjy6AAqM3G7TXEB/op7NqqjmU+pwU
02lbUYGIkaYkf/lFQaR8eGUEr/GP/0wxC1UaKsgAE8YDcFUMHXCRSqJJ19/afdZQxmlUABQLZ4oo
YY70/6mizwFLQMaPI8+8Vi516MRhws1H5FX4wbebqy7GQsqQeYOpjFPA0Q+V41/t3nRKrCpqmzNt
mKMvxB7Uzmo/awvTDVR7O4v7uVRzzidpQStAeb8ebLrBMdYkNVvrYarvlk/JlOj+cd5Bwq0qnnX2
xK+GYCTVSxn/D+uBTuag24HKi8k4u9vNw1anPgJWLAoaMyVi0Sxdo+og2Nvte2NFHl/DelrBBCRM
2U2pQg+ThHy/xJQHoEaWwGOrRmoQ/Olj8VIYEnOJKeHgnKiKj1OZvDzijvDJ/15CTQHEy8aqYfiL
eSpnOAdq0R02+6qS/SdIbRV+liwzo3VqzJYBVS7TVo5hMVwlJ4HoCb8Y9rbYB3Bc7Bin7yeOWZxP
e2Z37Lh9gUpKcB0tuVWGREKpzEaHdMpz3/gUFx+ONDyQCzx3LwsdBLohAtfB0yXj446UhDXuY60a
6wnMVjCyZZMACoMr83Mbcvmb7ZEc4NTL8hfszlU0mCsEhj7fqDcijyUT7g6FrIeNoqdl+XHFWJKf
ZdM5Vk3wj9r2tTnatwk5KTPvcgmzW3b7pYiDoZ2lmOkyPXIsIFNQFcuF4bmDxx4ZQ+4FiJhxXLd0
+ngUEkWwE3AYCTl/r5iRL9UCblslatyfKexYqUyuH9KWNYAyQc2aTMm0MqE/pvcHXu9wkglzqWQo
G9d9NHBOdYiiTIlDswSnwmeUVBIxtN3gOvt+7u/2hMV0J7/qvVn8equfoK67TT+uluYuJzv5ivkm
6k7MzxkeXTPSN4XkG0zk+Q+NQTznLRFTDXHhAa9rmcKrVpS38srEuY/SFPI3t+XmM4n9cMMB2xPA
sOQoE86ufyu0KwDcuBlxDvMsTyt7shTNhcCVYpajVvzUGw38ospCeGD5cIr/88nhuI/Gv85OpaEv
QkWABUOh81v2gp2eWjaEs/qzBwH8NlLADFtN1jRVfcFGo37it7tw3bb6WK+QsAcTYjww81TxhDDN
/vZ+ghx7apprvAFl7Ire/N5ZhQDgooesrGgAVGfgQFK++BWgjQqLM8X7UJxos4beV9xaOSufvE4N
vQrTkb+3g7BFz3Vj1DwQPfmjeTLtnVtod9Tf/mjey0s2Kuog1Y5vexAoqomnmE9YoTTYA5Av+0/7
efGzcR3jBh0+r1L4LOGRLrhlEQoH1rkalbTloeTAjvppzGFdQAXW+9I+SrcCsf66SL05e4G9Rx5D
3TeeCpuliLed8VICbkYWzfmGFCj7YbfTkPBzI44vCDaHgRVMjHE6bUZOsZkrCWaU31FZcPOd2/CU
SuYUN8kg47X85Il/41Waiv8HeX/cPsAguZmJ9hvWWymaqcbSh9ChesBdy4Xv/z+PsMhHmW743LtF
+Jzv6TqyuRXFJQUJ+HW7xGMC7jUAWm+3cMi0UGw65Vbu0iL+1jdt/xKJ5soUMO0ZuzdRMOmAQOCo
Lm1qOFcubrzjXuTo4ghqxNjwsId+6tS7XaAqepvbqmEFYCJW4x1Byu5tRQ5m3nK68HI3exaaLPxv
hOexqz96ZAhf+htqlpc4t7Se0lqxYQX9nVqqFoQ/tzsTZZeBtYiwG+KgSmptpIG24yGIj9+PtBTB
IE63Q9Vb1pvYdEVzwJaa/FZUeH0iLzlNtuNr1Vob4eb6apywGXFB4nOTNUZdsnwjZmhQARsQBxJ5
TaJg2MNwX3CbpkebktuZ6Oqcm0r8y+J6FsJeFFRJBMWl+Gz5S2vuW0PbaAGD3x/wziBruM3OpBpB
b38T9JEj0GIYuq8hr6MwbwWPMNYuuh/XKMzk1y0OBmokhebLspA74GIPPgBhdtHfMcudVAmi2Cuc
cNewFDkPHk1umC6JQ4Ur1X1GIXllCctlIPCyvHVY//eKOmziVMqRoj3V5Z+Mvh823ygE2wGJrtQE
ydB0ChLDX8wa11lm3MoKowkPUvz1rzWcu87551jlGvJ+utWH3E11SWDIx7n2tQzo+3Q+Kbj1qq0f
DrAtaRPibgsMqJagErvRkFifpe5oVl1TSeEd0WX4gtP5dLvN1ump5b3nv71TnkQ+xzCTLorhGKlq
OY1CVazhQJU1gRcpghJh4zDWXqF/MU6C/h7D3Ni1PJMTmcsLXsc2K2nEE/9ubaMX29Lm57dCGkDx
WUFw+8/ghISKXmx+rFNbtnyrjZB4O7vUse1jr3DO6rbeMGf/L7biiHT3paqAAX/jvwrR41MILUGk
MHnKq2k8xi8S1bmKsnqCci07yBkVfQZUIK894ezyJPDQfeW1DWkOj7VXP0u0W/4Yh1GHQKZBSjHZ
D5AJrYxlI93bZFIMR5QzmY7PkDvZwwxqy0Xi+/d4qjKaxVHiz15tG7TH8ecXHoSRa7NMTFkFfrTL
hw7cD8B+duPbBd5TZlFWMFhMDy1+u3PqnVg2K0hbJx8Y8wTqzx4Qnm9Kwr0fkPWwU398fePlqosS
gmkCzNvHO3BCSOBnmO3PvVowIyPdhET2sHk22S1nq3a8YxwQZESCdy37YIotNsN/uCFvV6b92dyF
xqfyf3Tlxp6xtTJcvnduUHukyKk6Uubl2K29z0ydm8jZSPSdI3rXckwkf7vFINqYbwAF6EZm12Nj
BrrVEAQKw169BVuPvhArKj9QhsWg1l1FiGMYbhtx9pwlVu8+MWNKTZM0vjAEaysHjlkyVbrvSYFJ
TnUxcAJJ4BGD5BmGcG/3jvcJCcW92uo0q42+DLRsRk8bZ9LXPhmzGLmoe5UgriWphj4bscoKnvYg
0j8063R4D1IJ05Zr+Q7KqtfNBkm8DQvKV9r3ai3D8rWOYW9UUTa0jhHcEDAVaeAGKVeOeZOv3eT/
io73KXPqHW8t/kXFfQF3C6YCbp+rwCOBwGa1Y4Jh86cdZEksY4DfuvsnT4fh3YJgS1VO6BFv3iNk
oy5nGQTXHfMqlOZjbf6U16By3VxRRqmcJFk0UxxH1Ch71hrOR7568FMosbvELyOeA1KRivZxOfSM
91efRIA2s38Gsj8TTe5ZEeI7zRWleImpPnMVTiDHfNnLapwujBJLYOTq0m/YvWrL2Aab9FpoW2yo
x62g/8fKDRhJ/OB73xjzPvjWD12PP5kgL2lylAQUu/Z2+JDus1Awrapf3MGyN+bbpipUh42m/jU+
GxcXNzikMQ1s6SGSAqQX6nq+jUMiXUvruEWKuwSv5Wxz3HhHz/8NX+s8ayAl+v/1vfnlmJ6kl7TW
8lohJNfLSOGtZ0Sm3OmJUNBlrrg5dtx6YkHovAe7zJLxQNMdiqJK9qNYBJDzKqGve1zxUuK4GMqt
cxy4zS1lBqHFdgvTaZ8tiGtzSNGGHj1ChbWpV2T3pdhiwvgTCZlRLldKqo8Vhntsci6/sXRWsCTm
Zjlxw9PARhpqnSihaPye0McLicxwipzu0LnVRyBy9kS27oAGcFnFlzeXk/y+ZG+/Ib6L1xfiof8L
EEXHbLMQXj1MKVzb0UxdDWWpsWfOOyn5PL5+rCRZNdd579M/5pjoB3tWhEblEbgCbHX8u/Od5CFq
yqpvWsfwQ0DWkI77YZalpdBEwpfs0ij+g9BOrn4k/flY8+zVE4iReSiPhdG8mqr72q8MIAjo3SC/
O/anC6UNqlblBC8zI+HniiVc3hBFQoB1ELKRB3xXBJcO1d7mjjzDi72FhAOfAI1f5c7OuMofk0SX
dKo265fVJToQCWfM739bevLZgkzzyq6dwz40PdeU9xMpHtbm7NeEoF+VelWXei+0hHRjutChf7Qn
ISo3NAXrfO5sXADUT+XsdKJIQqgvzE9+S5huBht7vkkRmfTr8g0jS1/XccQ0tqkUSym7wCl9hP28
xBddymAhApjnkJ5lb2uXR41UWTyTU2J2ZRC+pIOLsYTXvxFzLsw52UpVnFPzabGgau1sd/DDSSEr
43UyjeTa7XEzIE5IkT6rcwsejUL871hIcNxr+9dSH9//CmU+dBKeQhIOkYFzVeyt94HgiXZrr6s3
xF3S8KBU/bCUZ7w70UItTZwzikdJeJu5L/EIXth9i4OtJVKPhtHhWS0bSJ/Tkcx0SIdjrM1njLYh
2FYC2m59w9fEUt+crPj2SMwJmKlKU5AD3JhG172hYs/cRUKUYYO22EAxMtISI+naPh1fYPLjSj3r
pZBljU81jRhUAEDD7g0q1JhBkXzHsrJ6He0iCRJURcTF2jYnDtYadO8oHhNZS5Z2pmqIrl+vDv0q
2+4TS4Kpkp/VKUtVFffWn0UVCvkmixL/NbLjie4JbYRI871GG8nSOvrZ5quhbv0QLAwPF4Wz0PZO
95vG8OQIK+GaCR1gTyfmagdOTEz6ECmO9qZslWVJqA74gYrd3U7M+dV/8P5pom08X+XniUJR/vsX
Iy2D1A1rpM+u52zIGWCNLHssqEQxCE4pcQMhwl1oVxSvb+bbVo5nNgs4+XFV7ywwf1xDVfdfNGVO
a7ziDVZ9VM3pKeRFd13AAoeX/7ZWBICMjUzWLf7KsfSnhoNNFOT+cBoZZYDHZQm96uoVlfWIbwJB
IGJQ4+OibFVz6YawMiriTW0ovn9Wr92n3zRrSXaQ+02N3bavZaW0LUM2tnlOSLCZEgQaS93nCXwW
xb+nO4eFz57LyLzZt+t7j2TTCz9CsmdnG6lcv7oynNJEsZVvVd1gMDTomonmOylPsdG9proBcXPg
pASkwyICdWIwBdhTNE+Dldks7AJyrR1Q6vX4tsHZ4n3Wq7J5OxeEch4CIPk9+5+f4tAB3WJibsv9
fbxcl85Kkdnsz9ViX3n5UlUiAnpJBd//v+ocxuvqzftuxEPsyt6C8wyeqjcHXWUGPF8/5dV2L79I
ndyaBq9e0J8vWNArZabJN58J96sGH2f1AvkT1vW5dwY1kLla4OsFadOyd9K6hZd/7f5w1HXBoAp8
SA5NhUdhEFpKjDMkm4ZE+XaD7xLTQ/Euh4wVhd8rMIDe7J5ucaa//vXZRRRp9A8zYi0rn5mxvo0J
HP5ftzZhXYM04VEm7KPglRwPVjsUtIr7MnHI5CH7SbNAAnr6ylpcRKdIRERkUGRXoDAmHGq0gFY3
yU8WE3HqwOV8RoOHo8FAdQMfqwA9XtwZlcwVyd1PhdXkmforPSFbeX9wpQQQ63K+bjNFP3Q/amod
DYb7yWG0/OI64IVaXQPLKdzqFRf+rC9//d0RV1KfVQbNHZRvpIk2udsIhiaqXSfUmQcE0wMelJhr
NpLHD/l9qgZrqAwwN5FmDoWOFX4qLHC06V5oCQK82EX2R37X13GBPP8VIwNVegF5Pf29Lmz2N5+O
VPNxn9b1Yp0aaNWPNeK9hhi4//TaHS26LDr2wJNdgR6dCIHBHwmus7wcSUUEn2hI/GiLXKVrVJLR
1ayd8HmVDzNYesjl97U834vDOgsIdsBFRI30Hwa9H4wdYqgecql+VbLZrDez6b0PGsTnEKx1AqJM
TIwZCeY3uGfEZKUC+bFtJ9FoIyYjzmwE9KEpX94qIiGpXo6BaWb70tdrFWWU5+lciqQsiD+VGezk
NZicSbBTiEbCVZkUrVT3ufB+W7QRQvKb5cV5uj6KNeKe9Q07m3+q2oOZq5qZA4XMQ8hpASqCQ7GU
Np1SNDnhWyJRgrPBvxf0b6RLwKX4mKVgiXT9DPVM67lB6Jw2IOsUu3t4WWed7TKh4oICTSeBQnhH
+dwuWphSFdUznknciD0kE3eddPifD6vedW3Phgur2xyM3FdsLVNm2RW5+bS0qoAKhhGf4gAtdSch
lHNAbIz3hw7BrNvSyiQKXiWcPeaeO2sYpbo8GT90wI4hSN/bDzOwqDPaZ98G9WSBnKj61SB8SwYU
TbWkKIMXeY/KL1WtDM8xUdasODqczTM93BOPf3DNmkuQgD9NCh1ZRus0g1ku19PDxEsLIs5o6OsK
8pNGQE3guoXXnNv4qxcfZuEP/tAnDQDlxM+GqOzwyPc2jPiI6XrhgFxQvTQIulo2sJFuXz8LcjXr
YailCDiPuOQWC8YvoTz2JszqdmEftUt+J6oC7G3n9n59HgiOGY8Io5BMMFBcH0XVRC5gBL/hp2ze
wGhn/xNYf0rTAJxA0JQkLcVjqh2UY/636o8xfJFEnsV4bFn5RvufbRK+5iIEc2e9oUNYnJhVDML6
hvTAdeZlpud5kOqq8KOE3T6BWeMBX2JHMEXW3LUUGvE0xLfxXSacd+Dld6RhhIHqhn+/pJkXCUed
UjybwXJEZCImApSBcT1siMXvmai2+f3mwMm2/ADXt+zx98kgKq2tNELjxauBHr7dhbHU9BceICTO
ARyFBqPBXh37SELL+oxYPdMIRJLU797DCJm0VdyW357VztwLFbYE7vVn99yabUrxufL/QIHpMezA
b/K3hCm46VnqDV3GfxjcCcfR8EN3AaWNby62pQM+PRcsNwCARn6/S4HJ1QGhDfJblV2C10NHAQ72
QbyjxxWuM2U8f5RQVNsyxiai7fAm8Wrfz3988Hu1JQbTrYV/eH3KOrTkYcfiuF7YsP0UF2Qg9rkx
E7gcfWgHGl4kLWC2skOKEm4IO9NuJhEKAO4VWBskm/OISOqST952oJRHrCdzV6guUae3DxR44IKY
jebYtM1gwz+MsDtsAJGFqUpu9C84hOp1h88Mn5X3B3WMVM5z+zfUGLyFC/vG9hjkwLtsa39WiSnb
z0jp7yNX32FlQD1TlASU+0lW+gkHzADKjLRdjcR0ct82FphCielXaHENtbZiPMMkxFusjQXQnFdh
Z9OZoJKk72aAoi6HZVBUo76yutKDpQZNgksg0NbyPe6yczhQJDjNB8jevYl6cofJdFee9ehxkFJ+
ZvMRX99IxFts3yoqkP0F+6rgTxNnY1OFaXTNujAu+gViKgxRWp4toP7qhnojVMRo6vWHinXcjtfa
CTmw9zbC6HaS8+sgPV+LIKlVOQflfUOZHFMtKJV27oIM3bzh5l/0IQuqkjxlysDGdB51ryU9IMkR
RAOn42HhK65Bjw3tKdhlJNEeh/4riwHHg9IQX7sA+fnhH9sG4y1VDQ2lgtshkFwg/B2r+u1hFbc0
AvEHcu/imBUeXcLaR49G/dp5YmU/n7gjpBYb1SxohMCP3aJ34JS1taWkKEs2hYVWlqmP6dWZ9t+8
6IJ7cZsSa54PZjNWcslnvFs4D8LnGBN8AEZ2FYKVlkiYoqL4i29gqb1e4jqu+N1HAMfi/Ygj6BLj
CpbNChIICQ1ZmyE48Q3lApUsOo61xluju/Q/wnN+CNdfS4nCFmBKqpfzc5V4Qh0HI3eFO5BU2mKP
5t7/WgYhDLS79MfaO3sQDjlLerTK/mcK8PtHjg2+EnyFr0Wppku+jQia7uQVWjwuFloJ+F5d8qaI
s3jVsmyGLsD70ahrJtPx+NXdJ/ohIIHgdvwyt6Jest8nv7keQ4RIphHosHGR1vE25HJ/9SIMbq30
sBxLY+Vm/A1MT1fKpTso094pCzH1+hCLaZ/k3El17ghvFCF/lgOmALWTZ71jHDb7mlhAPUmoKy/V
HzUdeQ/7Ww/dCTHw0hQJKq6KBSJlnzuOQJEOBD8evoNU3VB6gJzucjtjVV0JUCxQFHAp7MS0Lg1Z
ERV/WbfTskrGZgOEiIkS/4FobfHuo25kpeDahekpj9wTWF2jmbMdQpNjDxdqRZRX3M0H0zsyBlIa
oL6v6NwbIZKgAji5VTM5Oa8cA6BCkisLI9PztVA8seC1BsIQGZZBAI4Mn+KXOtT1EMlrBZlbecO5
GHFs7LUyOzyrjKpPIIKu8inkKT2YnZrkZ0hNFFCde72TyZzUvLcD0+Wg++Z34INA0w6o1RVV9je1
LhMFfRx43TzaSVfNUZuhG/JoAILiJa9dz9WmTY9xMLCZb9eBWs4XXTN1HoL5VY1dqRqqOJ/p5E0b
QXSoNf7A7FH4oMIz6ImZlp7/7bkF/1aTnnjqhUeYUekMFl3ap1xJN4wrYW+7cc5uLDtEo8O/myX7
IDD8XkIE+rRhNTrTw9L2FPpiwevvxLvW766ZftBnOEdvCbaX817bVM4k37j8WMjNBXe8XIyp/Qmt
9Faa4rJ3VwOhgVBZhnNwEhmN/gUG0oGpxbN0bnnLerE4hFfunI0FH/VFJAiHZ83xCxeOyBKiRTul
GO7S6QKZ4wvRAFcJnz+ouWPYHr8nWJCDLM7Ljja8HOUexVpzx8gJ8lg1MlD6m0FvH4qXbyjZppLz
NGhHAfRUne7ZoHMUwLtT4oEzyodfHaWMHMzmyRCUTHntzAIPrKMHWZR9CD3Ro586uvkSNOe29UzB
FtxeRu+jjzUacj/ExmgUW9wO94Ws105rscgixINlq998kMlXAC2IqYHjmIvQRpR/758Wny0yUn8H
LJPLmuPQXN5w6TZXikJTCuRrgjb9wwf9H+WZr5wgL1mpUobg/Qp8BAxJlDqP9QJRhczdt6L7rg7P
I8tOhKEYBvsNkO+WqC1VMfknsOBzi0JSDqOANCFSML8ogOlqZFltg0P5GKYDw5a0cUiJiJ/wUaFG
r3LL1DlrZ0Le9c58nxxO8TJPKWnLwGpBqQ0Du2TNMqC4hrp1rPxU+aSkPVjzyeg0+p1AQ2j14I6u
/RNfuZ0pgo13vH0FInkYggd11OgGQC3SscVIIIL7QmxRUNwb46sSwUjpAyNolg0NrYalF0z2YhF2
sTJH6bLwJbrb9CgicY07nMMSd8EwWLujwx63AqMOGbuIwVgKtubRXb3QzbIfqaAMbB0YuhCGd3V9
ZPXl4Dclt4FN9mg9kIao2twtZHxHvtCmies+GVvuOoWaftTzgR2KWnxjfpBQhNGc39GL1LBeJNFi
62YmAgotPMdw/vAimB70vqz191qh/CzKKTAdDzrxehyQ+MPEKLuTv7Riw/52f0WsQdSh5DVDW/As
XHftcd+vXRxsH5sgZ95LQTORfFmrm0fXkv98eDcflfe4iZJhRQW4KQ0W+wfaPCimp8NmjKjkL3tC
6sdgnBRnHPKWzvB35pIWEj6RfV3PD31aLR1qtXtLVpiWR8DyCJULTddrgRHB/hvh3Daf9Cvij2qL
QX3q0c9JxNisAV2SGnPpontgH/5zHi9Y8DDuKDv/+KQSla1MkY1UGUTdjvytlwKUWMIPkP8oE9qy
aa8YDN4OLgvxuOEW0FmYnJrKj5uJsjH2dyzvseKjCUGCzI0l+B8BIWE06ktGU8q9V98yU+2jV3Xc
ExBgp9GkoW1W9WZqGPTnGW/4GN85ktEaQ5kihyCHuhMuHeIzkHQaOOvujsX1zIOr3O8h+09vvm7i
gT4d3HdI31VKn59KAifKiZqczq8iEkDwOx9WBIUPMxZiOyRv4dLWQPB54c3OnHf3A7caON26zkYJ
rBykB54UzE2up1XU1fqmb0icaKOHbv9gICd7ubzrBl6IH/MV73AE6AR11ihYcWFKPkPWupdxCSXu
YKZLuKKfjGJEjdqZk6hJL2EmgYNUw+X56MiLjnYjRzd/CuIfmtCVLiBgwDiOhLa2qwkcAcarUkNP
FOCv4mAGikyDKt6/H09NlnqFb7lEXL5J/2OWXTJw6dCYUIecyTmoyr8zqG2dLwvRyGpitxLOuQgY
zYTiXkRFyQk825ktDUdiCup1OspJB84YmvVpcq7nLXnzqBRbzO2SPeCy0YSnt/Zej8YBBeBsvM3o
moh4xrE1Ln9/GrDTTY/Od2CMXIH0wGGYMf7EZJBJ6FcBiRADhFghDxYJuDVceSA7dKmBpGUkqNN6
6D9ybjOjV4AREp2Djbu72gqXUT0EYZeWtG6UHRYLdWNhoPNOVALarEvTKQiDFGtuqUqj7J8zb5/K
yBHl8pxUm+nWbBwRh1Tqw0BFS9MSQI9PVUmLlrS/Cx01r3zJf5xHQeBoISGWSTHDbxvtAGGbUSLx
E+7niMrUYL3j5TCI8gwZsSG/I1O8A3JbPI6shIswCSc9t1S2PjjkJW7atkYf3K/EmvNcSSNMX0Td
QGwe/zTWj6TwFBP4gLcpI+7zWZiNyf6BxQ4Mqkvv01eJewj2LB0MrvgU89csfxiiAE6PIqoe1zzN
EHU6btZCIaNTfqHykzp3F8BeENRbF4l/pO/4dyKz5kmyxSrEYwgXLAkk9zEdEp4BJcSgVr6wvPbA
fbvtaEzoBanVygSM3B7uJovDw5ZXCfgFskSG5za8FYr+24drBvdKdbgzgXKH14yLpGX2nXz52BA1
XB2b+XAB9ZsqQP6UgwYGcer1FlGqZZlYekHquwoaokjdC40nVsZOlROeWComnDAEvlu3Dsjrf5fE
3xYP/sgGia0dOSUp5z6qhoky/rIP5DJVPzN8mNIPJbKaG/h10CuWCYRJyODR8bT/I34MQZuZN6Ca
5MKQN/gYPudjiDl17s1mNNWQaGEyaffQRxdVMw5Enkps6cn+qKi8NVK9+CSyagxrAGjxTGOaUDPE
GWiEUdoj3HWCvl/0skaSNIJCyLC9IaZ9xxQKmsI8Ezz6JnWsYLZY1m/jdhbPKXbT2Wz5VALlaL9r
vJErCkOfLtyEbSrEKdIIUmIV4u9yHQT2coaIlVBth5EJU2zi3wZLZaV7anyljInBkS0g2v+kjioE
EvXtizZDe16moAamKnoX8ADRrIgf9UT19zgp5hz1IlQe7itOd26i9DDmc45xtJwnEg4UP7Kx1lyn
ED9OUMmpu/oZ3jbd7pHpO1Y6dcvbJWKdKJpEZCllBrOk2IuUYGkbYYDB/5Vf+vm8z8sgnv9W6qBZ
0blneRGZY/1uXhtX/KYGvsa9ZHSKPeGcHER7tBJtGKt/YIdSHGsnW1eW93BlKdByksCl/ZwuvX88
VvL+ElwKoaPejEfd/totZhrDYZpfNnWir6HGKBO/HZqNu2Q4Ms/9k1GGAGdkvjpZETChMlDv+6Ec
ggEj/Xpn8iSr+57AmzzCeTSOyFuMKzn1ERcg09keJdYk3bkj4BtVn/JC9cG7aQbglM9aHVhzn0Wr
S+ChmBFHj/VvjVAEg2nIguyF5Z+nu8/9IaV6QzgbA1HKWP3YJ4PSu7SlLT4nddgQ5KA/09oWoF7C
Z4h3vyFikhvm2TpvdMvWjs9RkfWXsadRhyvy6vnTftG2xOe2Ep2hxrzJF4pP3mkrRM9/VIfvUQ5x
5yKjiqpLDpGf/0TO1XiVj9WLGqu3DHcjxR0vFVttgVXhS4btw2r32iraCaUwPQINB3/1hhnZYWge
C7qOghWDDylPB6/jNQxjIIHebDTAEc+AC5wFkNWgJ4GvhVVROqOF3X6YNn2FXStE3StsaTEJR978
3nmwbMrJ150Jvc+syr9D4Th4nW3WD4WA9RcCW5/bZxnf9A1tcDpGZ4yGVUSGY06ATEdH2wrPSG/i
s7e9X7bKLhHtLO/gGT0d6jG0umF9NEwgyhVu9Gau3gWfLodUg/T/Yq/0MRf+/qoVtqX2wuvtJReh
UgSfB7sUI/XpFbhhSC8Mq1ec7YjpChTNwKGVyWS0lz+UGJs8hM7GuMnvPQaE026GdU+eL5JJW9Ui
i2ci7aT/j5mHK/10qajCsIOhiaklcoIUVT1EO/kevEuARYjFyMHvzQWp7dLsAcrkyhNFY6FkYD4C
5HWSy8j27gLLXcPu4tGr/FKzFtdLvE+dDtnhj+eY1WevPNu/D8suX4LgCRf2w0jsa1Ovmd8ewwt/
fRYZTFBiRp/IQOcA2nSXl5V5GkCsMAEaUHXe+mEHixT38Z22vZ0Ql5J95ckhd4Zrl86KYuVCpZtX
aUWKKvbLMCspYNEBGMnimZNLQt/nLyVp9+mSMU1ryw9w5YGBKDgxI8zr7KwMRMrEETVu5Ka0fLAr
Spl/ub6A4JIMXd+Yy3PaagpZ2AfQhJcpBoYDu8P3GqMbypWUxl3sJOCuQNPhziIoPbr63mfnka4T
MjQoCN9jQJUPMIE7+yD/9BVw9AlRN+v1IiEisuU4m+k2EZSr6xUaSZOBiSmArOqj/GwUSyImw7jK
dWZDWXTeixlg8RD0LHE7uBBdIf3B5eI4jgniBkLzH/7r/dL9xorjrCKkcZ9PRxRDcsHZUtHJXAb4
tpuRXUC4cba6YZWHNL33vw01D8YHMogW9L0e6UGcPSchkds9UfFkzPCEHgAJDZ0aZN5hFrel3Xec
6YVg/u65P4ckCRk0tRMhMhBCP0W9doO46EUp7N7TcIEfH0auwfdWX0CiQkiEM8Yv8ozwKsilq+fc
RVkWsAMpeFFpr85w1UyOiVk/JuvDaoZesVYfg/D7O3ElPR8ZSjszHksGA33wXmcpan+azRYPAdLW
0/a7jQH61IFgIhn4RHVvVPPSY9XPwKOoaMY9ovrNN+EZ4Dwt6T9rfB6F7lMG8pR5cqwrMiCkhmkJ
+9a24cojY6FdyOU5eEIx4YiKeimqIMsPIVdZgDr8jA0PlMvZyDORkHmKTdEtnjpnsOyyb52LDWap
bXSecpnlvRgFPgIErMOV6wPQ4Nfsh3Ts7QzVtOmtMeeQ6+M+NRp5P2hbFoQtGMtKca8FMMg2HDsd
jgQu0QTu8Me0lLDzOy79vQMOBevSHrFs1qVmrUgU/nJppZJ3IbUiB8sGRuchs0F8dPjOlxpwwTI3
kshb2gOSHH/bZv6tfALmwQfQzDKIRwS3l05xPdCBcRpsLwMGf5AFzjS2VKOt/jCVT5qkR/ugSHNh
k4xQJW0YX2Lq7gUsaK1lhy9Lt5DNBJHbyamDY4eJSjy5ZczZAWewdIPARX3gR9zrqBop9J2xGwKj
Bu+RqRpmxKE+ZsCCemlXOmxFpywlM14DAByoQlxz1PaTwoa2aRYFi9S4J2nysLt6kClMs6n1ojLT
LHv9il9idXXR5K6ZT+b/8TFENIr8HS+7/N4MTUII8mwl8UpqI+u7yTRD4B3wjeWOgW+Q1nLLhxnr
RdaeVvjs0kcOu945P/dnPv36INa94Nx13Y6IDotVhUL3Bj8EXaO7/Jg1Uo0tVsxcgxNRLcxVCrx+
y6MwKdlEsK8i9CSxvjZiO4VUsnahaJ/qFFsK114k/OccCNJ/DIlaH3PTivX9GxCxx0C5b8JNY3eB
mDzGhDDoAdIF0/rviP+NRfIjuZhs9JwZaGpVHrtOcAQkTvLjmaz/xaShyFWc/e6b4w6cqhPy1M/e
xt5owsHOZ0wasZpGdQVIZqWz8P0wabnlx/QzEBSAAW42CXAdsbsMv3LGzSJF1giB+Twxj/K+S1wI
+Uf463ZUTbZWOvX8PJfjxobxjr9pG4OJxNpcaz5nUBaSix2sEgsSB4cciwFL69acbEYUoy1m0wIY
uF11OSQONL823zVrVR+E+ejidTa2g+ITEUAwphzidt4h+qbubLNEmsbdzFpLEiANUSG0/e/g2R3I
GJ5+k2B5WPUFOQh+tQfRuWytOwVKQkKjs1GJabWA61EHRHgablgDwR49JhRvY1xfbGEG0Bd39V9w
x43tAy/rv9ujEn/WGFRPbEmewOYzeSFpQXHqkGskidGsTNIMvnkco4PBbVwumiWpiFuJQJFEt6+m
o5s3fa0cF97nONcYM7nWuF5sdU4Gn5RTM+pKvjX9VLsY8ziWooA0MPo8gyiJ9zq0upJ9x65h3Zx0
Hawmaf4VYgWO3YJz1k99Mo5mezEeYar0Mxk5Fp3iGaEHrk/pkRHVvB05QvOGL7ZI9qmu84IU5uMh
u2biJh1V171woLDqgGgOGpN7nXlXgarPAL6WIM+rBLu/CCY3EysPJ7jIbUTc6yarl+Qr7AmAdCaW
+/dR1WigRDZnPOxZzX1UUSIf8N4cG2JOYn/9ERudWAsgHBUblHWQOsQTvwGVBT/XzQts05o6k89D
cTjjquO36aNWwQS5ITN5KYpGNPIdgkPd7DrQwfJ+1PD7o8yB7pntaiY6u6aZu3rCwnnt7gDPH7ai
ROZF1GlMmfMkrwkSVLKzlISBRvPSr3+/7HAXZrtJuxAYZUPiy9BeUKlQLdv6v/FlwcQ34P7zfU2B
/AT5FITrKnBkqSKREkACzm9Ks8iwNunbAFL0CKwYDIaJtAfWNSwRIvOC4u/7dfpZH3JT5RHDVb9b
qOM9974W1SuK07b1aA/N1mjqCWY2F1Zxm/ULTuj1U0qpRguewnheOKTLtzzcECPDEADVuyuWD7rV
UmwwqUmXWjcu0S5AeN8m2SAGBltcvOwXAD5PqDU5LN5RNSH7ahaz5reh0L6fEAJkJ3d96FgiyGvl
FF1haW+x3r9jH45EozTCuZoSb5djPpOxWKxqt/SRAVWHYBPBXUmqCyYP9XlWHw4YMFh315ISYB7P
U2undt6HKjIDQYLffn+RCPcBmgdxv15Glluq+SsZ21opABPEupjphpOWm2TnyYEvsSjgFx3gvH5d
AnZZnGMxH7JKtCRWXkqHV36e2nt9uI+YNFAhdi5TtBhph8efeGiZpv1kyQCiEkBXepkkuOcP1anO
pAcjMS3oEhbgtV7O+cXHpcECJ8K4TufOSrbtfiOqfdVKE9RjmT0JgcQnUeTUchzN25z9zQPVVR2P
0+ulTD/9pp8nYWLr6asAwqb3l4h3I9ywhjpE+obaC5Sycoj/Z/zt65yXHRw1Vh7bpPgRjcdYd+g9
ptOY57eBa2gd/4V9nIN8bFy3DXcejA1K69IRjjlJLk8pO6fdsu0xj/KfZMi6nMaBCsyNGoaCk2Eg
AuBpajD6n31pOw1sTU/Oy+9nKmqyb+ZGFugAyNQoZivjewh2S0ZXfR6RmgQC9+n1AWsdVGN0dXd5
Nq6FGrZmbcxLxUHb9BJLehyihOKR+L/+tWWDeGNswpcZ005kQJNOAMCoF9FzXlMG2RuHE3pituwo
OrENu/CmwzPBI8MO7gcz01TRyBs2GprItjEuURfx9HHz1AYpiCCXuxmUgnGw3nC75iEewTuzRQ9C
aq5lGd2Mgai/JOm70yDfYa4T450W0r3TyVDsaAMgE77njWLQFA9QLPlsLQfd9Q9SKLnYvDS0r194
VZjLUSzFc1PDLEXEiZx2m6FFKszrf6zMZh2tvnXDFWmDx7FX9sJB6iCAZm+UNlngzpRUDzxbkxhp
8dn9DT3GwZ1r7mregi1vN6s79jWKbdkycp4M4YvOssdRD2FKxOtTj31eEhyn80khtA1trVFAm6yl
E0iCPKoPLFk7pUKdpMS7vvo9Ha/Rgu6i/Ojmz6WLIr7iyUKZIXplZdgkb484x9SWfEU8nrzr9vaS
L/1Xp5vnetQJVV+YK+hH4H7zu5xShQY049hmqGUxOk6oMebxa+UngrxKeGxzlxx6oHXqKnQ0TMR6
528b8FaADSZgjRgz90lm59UEzL1fnph6RoPwV6zJA/2dr1FnFmt8btks1AHK16pct/6pNfQ6EpHv
q1wisoOaKtbJi5B2jnNLoGwkBfVMR5yk2ZRC22uY2yZb7taun8J4/VGWFsJm7g0Y7G2TCVFwloGD
qG25K21mPbIrHl2yXOORBLF2gxJ7hxGyMa3BmoAQjyAHH1lmyIWItrtHV0pUIE/OayRrcW7L6mTU
j5xM2mOSouSLWxtBGwOBpN6Ac7Ou9FjEolezuuVc+RAw5qNVhNJNIWiZuLiqVmIfxgL8dJ5oOD1J
Qz33WW9xV0+DI9HHM/BUHBkJCgwYZlY4AE4Ica1/NwOjqtXiTgQX+jyU48dIHfkRK41XMcmzO/F6
y8nJvkO3HVpstrhvsYHRyz1CFWs+q4SnfSfkiR59jgEeuf/SHoawYOVCTWR2ZgazTt7I0KDLs2E7
7PosGlxGfA1Lgwbrve7Lpt9KHm0t4o1VxMNf2rp1OEqj+OGoz1PpWm6JusYNnLw0iU5HIP4qAso4
UJfMgemfbGTdVMW1GedTRcma2M2Nt9UJHwuUqAG2JNRYcko1D2D89pFkXkoGZXoPgUuSqYr62dcV
rfobgE8mI7OZMsFFuSS3WK+0VDb8FQlxc/7JISgBaOWwAGOJAvdFJYWjv8EvLcCWgq/qGIqxFJJj
0YQThJEyYcvm5x2+MxHBStSRB0Hb+pxRKEjlQY1qwdmw/tbMVJ0IKKIIjCGozqiYsf8xaMShlWsx
LRdQDGU/SsbnZA8ajpl9c22KnY0OmcSzEE7TCxZBovJeFguYm+Romrq++MEGkjNUgkUyOI0j95Qc
hpMJzq6ohh2wgX0IA+p3xHcEND67EGmTiSu50yoMgZ3S7IzQcSmB8anUeYPNZgNvqogYmpvA3/ai
W7ldK1wKXDc2wnovk+REqVmj9vbpkTNQRelr+jF4jGMShV+OEBDytRMNAadiiBEp8pndIcd2APH7
zyzXEMNdlcMPr1gA20LCmusk4QaGP8XL3Fhp7LAuWFsMqjcPQUWBCEf3gVnYXtQX5oqYPMBpjqGz
uToZa1524FJlcoRx7/iMCt5BfCJ8vvbaL5tHmrFS5MKvGkiOPZFLF5kXqq/1udsld474LrPSuCBe
yh2FH+8I8SJ7GfVsYLQuP0AbxOCgo0g3gz6I3hvdKDGC4yUww/PIH0fq/5YPwB13GYXRtETNKG6x
mm3Tq6YaZkr26g0u1BbqMRmrMFWlMUb3H+X2+R47VuXcSTuW5KDBZgZqMLGDVGJdjRmnwcCOi+tF
57C7VBZw6DhRziEBr12kwnnuKPlXW18OsYIo63xLngQU92ohCW2daoJVHJJ5OiXYclzTFQ4zbQNc
YefG1S3hR+11+iTMZjOgqWHdnCWyYVDDtyLvBt+SCzAB0pDcXABtcg2Z/G9MmAQQcwEXlZ9jmITe
mHRnT00XzK63gn9WbzcEHivqrFT05ZDROQ1+dC8UTHIXizogn0gpE97xM5P4jK12ckiS3KsqrijK
1m8OR4KejuJ/ME2QcK/5tCwDTPkz2HKlEJ8bVSjGyhHK4aTg6e0fN4bQUBttlE5wiaiZwPNuEcLr
VtVcaNys9Tl1YC2vM5De0sWhJsNv5apMUNSe0uSgt2C0Q4wKTmH6nGfvTzVg7KecJNAGd+sR3puZ
FRjT9xR4VHi70WWO994wpqzws/Ko8LeLy53MSSF3dHojfldXy9G3i6p5T18jCdzHyivUDhSTWBxH
q+rMemS4aXpJx1FCbi4/aappRFGRrbvhj4WEeszCUIXZqLlHmlw3GdHTlk+FGi/aDvdqPqOLrrvk
mWxYAtoI0FLRhlCdnvZNDJCc3Fmui/0+3W7FfatMneuApEg5jZAyTdnagGe55Zsh6uD/JoLxwJgN
qd/t3tpdO41mdkUDyUEYQVOWfAaxfbUpyaoQIlE0NFHw/HqviXsjR0Id7bssaECKKFLmFslWTHEh
6kabCrMT2MWJSI2zgX1soO5rXH6AX+YgcXj+2UuJPKiitoIc1RenT6W4Odwg9ukaMNSOSTPdpswY
7Ks5NAv8DAvNrfkDlzroY+vGp8+j0TXeYNeZeHDsWEUz4+f0W2yIefnB7ToV9hlp7QFmu7+Ez9WD
wPak6yt+LznXdeKr05hHEAYCWSnP06CgoFeJtu4FPpfmYKjAQQr2DruWb2Sb/WdCweZ2/kGCk/lK
K4opiPMn3xk2DTnr9hL426JT0qJ9yKabDhkl1Za7hbe1aOAS9hHanPhQ0S3pLziu41y97bNjyhXk
wXrrg6FU58RRWIzngGSvmrR/JBtKQbY2jas4+T9FNKiMttwPgUrzS3YzF+oLaoZvezosiZgQP4NR
63Bx8wcRGBYTdyJ2gyl935EUkTOokEtnPvtnbiiGtH/OmDHZUVZQMw8jdV/cYWH7QBGujajjG/iO
nJ6OtVMS2mBn9i3rRuk9gyfg1/fSLW/h7JqQ3L5VC/Uub5xMw2099MlAx9E0EjdmakHJb/AhlQa+
Qss6FHwNUk+HmbwH3Q9V+fFEEZLKfPcnucr1UrtLQ8q2OJmmqo7NWRqxhiuXsO/LaRhW0jUOSjYj
nNz/eDCnOHowcr7PCheGADFVbgHm9KjoKjlUb84e22BRhcXamWCKS6nClEDGT+OvlkO5Y/k7Yu1D
7hW5M+Yn9d/wjZzlliH0/ck2kWiwiIKe3feRdyNVyesaGKNZKWkULp2GEFTLPf/KYRju2ikbMtBy
XNggr0MkoRqxTB0lMoABWCkdIPP+LAzv7WwRw09aRcfMYFXHTzdx+IgzpQEDhdhvuFOaXMp/XpuB
qQHkurGzv9PZoSJpPGJZ7TcezfXHBo7nvKWCfaLIKA13N9+1YY3RWXBakXaAs1zW4H62fJtUN50d
h/30dsnOu3oBJbEu0ED81Pj8F3ZwJyTzQzUpJD6yTzSQzPskykgkWVl+l8kW53TnzjGQ8gntRvs3
gtqBtqVrBPjQb5McfAw1ZkRTDntPHiMHnS7G4aJK7BhoW0otR/yT3NflbmI6k2srWmpo+SHS9SIw
VarVFI8b62I4vqtasDRfZgZGWw6ZzjER3LFCrQ02Hr3jHcFpKoWCMUQ/7Qq2ZDXIAyYa3xuvN1V9
ezyIDvy2ZjwbaxryrwzHlxo7eqO2gMD2cDYzIVlhk4sWIIPGRUBhhjJDn6pyThjf1qqqm30msXlP
LUD7thPz6sXOs7qx9C0OljxvJ+JtoEvO1OqMKRejKJpmMwh88MXsEHVkMlCyaxm24PxbiTVQf63w
43VutrxsOYaO1Enx2BzDeDQDqr4Z/rNsLLTdbO7oTLhJiOm2J/PobR4cEkg+tzGJP0fb6+YAXNJd
NpEkpq/N0EgYajC+5y+8Mbf1tR/JxGINqzUMZWf0BGjp3ri2+csvzY7ZVJdo/r5d3TpHPNWU/Wk3
SQ9Zz8idx6CtAqYxuk+EhlUYypWa/EQHajHMnH8NWT2aSb2/9ve2jdEsIRhTSVKlIY0L87plT/Xk
ygel0yYT6kNsFUeH5NK37FVAyxGfnPXNJNN/fPElwIFcGytodbZHhFJmZxJZw1Lhf581pZPZbOEJ
WtwxeJ8sfrmzdIB9Tow+sTUQzunoF5Bpu8198f5WbN48SNpuhlwsraF9m/vi6lE33paPqVYLmKNc
ZMNwQFHy7TRgBhxuekMb0QSkLhl/FG53i5hcDcRUoyjqKyPPAMlOrBQCCy6ZIGZVVr+J3tns/r+6
HRosb71PkdCuG7ulyj0Dp08DQUWr18UrOChnreJXYWbYpa8XxuiXht2GoX5iAMsY45uAeqYb4ZLA
UQ4qI1jkBZ7y+qSL28EiD0QJoLvrKm98Tzbvf3hKaDT/+qth2KTXiRwBAAA2ogv2vxaWKU7DGpr/
WE6c4qGqgUNlbWHBAu6PrnsAMdCREu7Jli3Z88F/tRXat3jdLj1gb8sefr2wqROROY2yJegovOFf
D/Ai3Py9hvmzb74fuykBpLLUPRvOZoFfyQgS0PTx0foOwzkqeVHHTErr9qYyEjNR1eOnD52k+3+9
+8sWf8Grg7S5spOc6vG2WepFMq/8e6iUV0R1cqGRLbxyso6n/u53WNgSUFGAtRbviA/ewGNFBjnH
Rl5qvO9G3TZ4IB3xQABXMVkIyZxQ4B2vbLcrPcFMsn9ywt0WbPsW2WCIx2RfLpNTA1d+V5wK8my2
2Dgvgo4FJsC9JyPfEIESZluM5X0Dv1ULd8rs1DLThwMYB0ynRN/lvynh8xoBc87kvLQ2c51BQ9uk
rZNtHY8vHVyA+3AC/XaqveRTtu/dHoYzZJQ3WV1DzuzKtGZCqXPVbyKOP9k591nMDa8nQy5yzRj9
32N7chj0KIsfqrLFo5nlAcgY4nL3hzeVU8P9k8q1STST154le0ZKam3o4cOEd2AaFlEZHbKIEwtj
7d3WVn1g41O3eM7U71BF6uIZRM5vDjeayoSQWUat9Dxu3LuChOYRJsC6LGAX41WqIRGFEAhSeWpE
MEtvtClug3/n6UFA9t54GuD4XjE9kEOZta+5egQqTKhpTzY3rzBem/JQa8DYEnTAag0yX9uU1du1
ZEKQ1bFKrW1APDFYQ/RslHI34hVtbnT/txX1x0MW3mL577GpVIjCBnBzHbUtXU0UREMb+2RInSOH
BKyeZ9WhqLPH8IG0WGFliGZRcee/K1kU8TpJX4sw8s55UW2IxIXZxgZICAK1LywRV3+5Xxlz9ES+
1jxHRxViE/wupi/nulBr3yaqAGFNZMuVLh5nPgj5ePOBg8x2t9AUqiuYN6jPof5BlcXWaN36AnD0
Xk7qSACEpeX2oYTFqjKavZOF4G5YEjDftVPtpS8WB2+yLeiWANlZWRqASGvAZobD+Vu3XK9MZ5Mq
t6hSp29Oy82q19IE1VXT6M75Ra8M7x1l3pXxDlqg+cLLYBGnzL5l4nZvquYtFtg9J6Cl02j3+FVw
w2Xb97drg8cfC2VdXjKVAnjMDf9jtC6sOHvbUARaM85sFXAEDsuEcVsulSNzJifX7ImEqw/4Iqcp
vBVF1Kc+5gVlwtaqFCow/OGWlILx44uVDOcI5NDM77bd+D6XjPnB1IMnwsmJnTR3Y3P710B/Ykox
BfT1h134FgsVBNHHa2tZn0hdmXQX2pCAu55jgQXU9Dyqj2rhKtG1KgoDGGVBNwjQhHqe28q87eC0
rPCgGpZ5vIwhoY98VgKpIqYPCvs1KHsXP+HE6Pgj55jXws9WJIfql5l1fDv4maBZrJBRxPr9jThk
TJlquYmFN0Trfknl12oxbhfTkTcXpnE7se1fB79Irdj/R7I0pNUBEniqOqE0gjmEBTA4zBnvaFbp
F+buXcK9hyjZwDC1wceq4II+j1iKNMZWuCfyrUJa9jzpdmaU1wRquO6BVGtiKuRGGEM+5It5Pl4i
jF7jEkrINADc+F9/cK6xe/VaOa4dwEreHwrhwdQOium9abkG8v8dGP1R/noKhZpFhQwr4lpZn63j
4I7tC2HIL1b8ib0fOQXFQY9GYX4qifPlqM/DZP23ZVtus9u0jxfstK6Uyi654fL/3EV7S8c/u9B2
1QQpfwGFTeRP9Lz9fR+qMSryqS8aDJ737n5K6GZQ6gqXsa4trDjBxkuuPJxmQGBisW8BkUnjSNq3
kDN6I1zQ1z/XjZCAgKoRATLwHcoWg7mKLCtuqWH/Fa4CLvOc/gxz1XocH3v92PHjhfJ39btpefmt
GH43GQIInj5lBaj518XlvkSjJ5wM1XZpaRtIZuQ8JNCG/VNfADHDyV8dC/f1sWFELhX1ZBnCiZAP
pyoL+kuFfqMwQ9UcFqIfrGVwCl3PDuuzzFUmcmSYcodLGcpH6J+8GhUTNwDGIjMOVWj2mL+E4eqO
vbhfWb3+V+KrYTPm1rLM31NxqfAjEIMBER1PMYiHl8nFUqdUAY+cc9oRI0TKUx2CDdHKGM4G3G75
6UPvB3ZLfuZO/zIhkQCS3QNA0BNiWfQzAmkXt5cuQMBN8rDZ0KhG26TJr2Org9q6qQgkqRaVaZet
M9qe/aQNg20kfssjOLjInLLaOZ9BHYGN0PvJjWwJY7qYX4lp9ixpdAx2grP/dFmKaJQYtZwel69a
xtT5OalvCYsN6aNMw3WnEN0f/c6AuJ8q6isjkhGJRtJo8miqYQAlLSnMJ6rULNoNT/dYCNt1fDh0
Pe+cxSi7Z5TqOqS/PWZbovO1b6MyL5tj+MpyzFLX6b1ze2zGE2dU4wR4gDyinvW/5PyCIHC0XBBk
NTBh4T1h1L5t9qUZ4LBhrNmHo/gqLbu8S0bbNfgbQj/889LfvVw9Zzry8Zyw/QFvc1xlMkV7Uub2
spYGWGCuhKCSi6K36XtaT1PWGKoPFR0cDMLWRf+8C6Efxc4SCRYKtvERtBiFhxOP1qxLPoYgG9LI
l3xDmZARSK4AuCcwe71A1v8Y9oFXfXu/FJa1g7qITZmYf2q8riI6oRE6mOOS0bBCGoxrk+geDZ14
HjtV45jPxwrxVoTwrQ1vfjFv+ygxM7YjXb/o9fxSDslpYbelDT5+Nv3hykoCwzb3Hvqui5LXOkkw
GvBfAKLbhaDnBFh2drEXxYVRdNoXwnpi4qBYiiNnnuGRGcnVsI3Xg1h7Hh6tYoVgiHCzP3oIiUtS
AmAMIQcFEqS5m7DvzwUHlyLkyc0Vljhz6uuayMOnhr9Pr7ck5QI05IJC9BLv3u7cKoAIsFS9dIkb
KafjNqpQnDWnmVq5vMIiKnn2dZ7/8us05MwT/5ee6ujxHH1QIDcRH9OMmztUcJCcVkf4dPd9EGZT
8RyKl25lczO9jdnE0SaeBwxV8D0Yp3CiMiJC9rQU5nsHcxwHXDPtF7NYI6R/Vr/T+o4kP8+Yv1oN
UJM++mfSomH3MQ0F8Q85wsWJm14ReB0HaaBw0JgQzi6xUIFN5gG4IURDkGI93w/OGys7A8mcZLvg
+NCcDFFEJP3gRhwIYuXg4RkuTq+BTItAsoQNrASDUO0Z773i+zY9hEpcx1ddrdVhryywbaTvnIAT
Vgq4Lm8EOZE5Tg6iIrsUcZeBlzA1rmATC4niuxEKGkXUdsN2OaFzD+mNeumdVT7jm5oPQRD13QQL
oUXLSEuhG3RPbHJh+zwCEgvCLTLO9wExPotqz25NTxY9PoRd+S6BrJ3eYpX2i41K3Mbh18ts2rNp
SR75bKvX2JFHtM/ZXwfuQz9PBAqAyWQDM3vMRAD8KNZ1ZyPGwESORv25igIhF8dsHlLGH8i9t8BL
QkZjy1EnBQbA7RYZxlEhc711nTBo2MPoyrtHjjM7sw2SKp76JTsxLDcrW1T/EiFAeaMOGDaxyeF/
IS+5NN2jumRYBge4nGI/N4gSwpeOlj2S8Hei3N0AKJF2K7DHMw+2vKmqCMNcO+5eLU50CcjM0SUc
vAAQjxN0RGn0305QKPZD3hMiy2ivzj9u+a0S78DvuSzPcE1qiANJ58hPO8jFCPLjU4Q2ix/TRyOk
T3Ck5T+TF86VF6zPE1OtDkwRhys7ncCQQhQF+FHtaEu4iMEZLnoLEY0ABwbZU2TjgBY8K9m0134n
m4PCLoRJBVvhN4rSEQimJ+iCacFv3Oey7XJlBQcZUTCtlYTKLXEGNFxJ1MKk/BdwKXpZfn5ECC3+
MQuFGWN25u91OUHLAoE6FeUIRiZzVuXF0xo3yUfjZq2Pk0HUU42yIdpkvbGBgYHLLC9asXKAUeGe
s1iX+YVzpo+i7zcsZ0994Yz/9GSUpIlqPwBqRvqet/sv9SGimqLVOztxrON9V0qwX/iFlpP6IDdd
NM49pKX3NLcEYTHJ0kOU6AEkGFgbTh081DcIVZSSsbxDdGEh+GBW4eUWOUYlYbNH3Aip9SWLLUM5
iL6wvivvzJCGP+kXktpY8PMMJcR18QD0FnWMwOEsrkwtJ0/wf2xRQlj7cCAvjxGGNTbkSL5Ga7RE
ftEnOw2zOmuK3vlqzREDF6vstChaRVrzuiBN0gmjRuuL/Gi3HxrB5NMCUOzjaVlY5IXyge9MyD0z
F5EChhWKRaXD5oPWqDwC8Pe4j1/kTNZvU6QY5pyxADgwndw8NuzNaMQwdpSb+SAYLuGBF8ERPLrp
rum8kSksNrI0WytVp69MhC65GawyDER7ny+9vb6SOciz8hgTGcsHKV1mBCcnaBnw3HeFZCasWbip
2xYVEP4xegpb1UY8oApXkAyQYwnRY/jqZNU41O6bVkneYHu4W6SSWpOUdqHm9xZQ//Cc8w40p4nu
z3SkH/1lk2UH2XrLEZIz5pV9Yfgxncnu1xCdEBbCF1cV4gPlnknLe3ouk/L5lnoVQIaMua/ktA52
vigadLb3fm3NGTs+v4DyoNSjrS0P1RpsPA2YVJu4NgByq+yy0h4drSqVI4JNVV6MkBcL584ZDTuF
jxd1q+i/vF55sp0drs7YsoMPC52+9otnHWleJ9JwNrJ5j1IoCXOwleVZEoxdsmEurNU1Rh3Z/FIQ
/Tz9eJU4dBlpLWyRniMAyi01ZR8gY4qv6YJV7tq6X4ddPyOwh28Fou0jOGiK5P/9zbO2jjy/nnpa
3CLiCB8ScG7DXlm+imoYFb2v/tL3nRQCwIOn36b1e9eubC3ChkfkRaEXnTKh+gn31Y7IU9vmQSkf
CNIHTgvXpVe/iQYpUZtv6/BXadATk0gZM31BYZr+YKSbFqkPtsGzFNWqM6LbHL0YSn9A1RuR03cC
EOOGVe9evH8zny7IHXDbfT7Elad8wyuxGZQkGtIbiiWnv27XE6pNfAsOtzdPHOhxGjrE/IN4eUCZ
iNH0GsUoJih9oeIyXNKsNP1x1djzjtf1NbOmHp8ux4GcnzGdF3udpaC/QtaXJjCmYeaxhBnPATzp
FnW/nygCXG6mnbUttwhLwjgEivtHZAtQO26cbIl3+m2tfwzh+bFpgOLSi1UM/A2AKJ2+IPGM8xp/
XxDVyWehZhsVqRU/LYOe6s2rEC7RonALz7KcENJnvMok0SKUvRwT9XVJanFLuGnjouHn4BnVy0XD
OH9VtCHyQjgKmT06Sr13pr6TuEjBts0IkyVWkmQNMH81BCGUKED/ATXKfFIhW7HJTAUklgWEP3Cg
2IfJGiOF0j1RyBYCSZJYn9YAT3IYU90kCt71n/9NMaF4eENfaF/JM25/8qWt2xAs718T8RACwHoD
grQvO7lpWuFiDfAQ71U46/fWwZc+2IffaOrfY/21vy3Xcz3xZDQBU+nQEMoE2Fi3mVXJKBAnzRMS
3coa/6zdiYV4K7Lor6kuluCebJDwjxBm73wcooeUQHiPs2zYl2W2PHE9ltmW/FhXOnQsK9VrqJhu
JubAcWcdM9Y/cYqYrmVR3cArFYbJChkZkLuu4b/2TSIXOmobEZsusjmt8DOG5DOGSLWViGvlyNQ0
N4DKorC8qFqbZ6vHyoftOVcJOmGwr7UweBylLDZRA2kcZH7nS/NfaZN2F6Hst/yz0gBJBlUdR/rS
RtGUu8LfJd+rg2rkDT7fMNqKatNDt16G4jfBi2XcXxVus/M2V2AH3uNCHINetxnSIxjP63g1iEW7
vBZntQhhxy/k3Jtl78w7GcWdWZIr++qw0R3ibJxfE+wZVzDK6SdXT/cqUXL/0UDZTwdIYN5PL6JC
wTwbJhmPdf+m8nL7/Zb2HGEf4H3xw8DlfGDKSizWAShs0n1ZYeQzAu2Lj+KvOcnVf136nH7oSdsk
vKwH/4I5AvJgnLH1pReF55wcXA9SEoHIFD65H02WxHBdtDOr6MnaI2YcD9Nry7qfsrAL8Y95RyZE
2HrufXQNe2vupGA2QLOWPcCCt5TWJ8na+Z2LZrDFZM7e4//7Z/NbsOtjCIt86pSeB3N1f+X7+2CS
kN15Ovn5FtI07ouZ7+aCe0M5BQhoVZcnufEqiM04R793cfnVEMlgyXoRbGcbHPx6+BB0I6DdW4ea
P/WMrPMXX39OafqVYTiPkO25BpPXJ2zkNODyF8KEOjkwwDJsjj3S0xA2o3hM/3MYtt+yZ8r7VW6o
78/nQOi8ExNQESjJhIGvXDd7/wuwcw+ySx3OxfiqSrxx7JtjqUVhHg0m09SjYS0xRX7oCy7bv5se
caZFVsXzJE9h5ZzMaa4LGdXSVYy1LL6c1NUmL4NpLbAh5s4i4BNJRAVkgMp3wq5BIA0uPp5gbeA0
jA9bptGFpan0uGeNNworyx3obFjXkOlxEsYSObSV6ReN+KnqBrD1VQgb+wwRCcSpaEsqfT7h/JhS
NVi1hNe6yUWXIfampL/YgOoKGMIErLlcQqsibmEhI9dA9cJeyJECVB2URLEGi8wYLSrE2EekFw8u
4qqZKaIh7fohh29TK2YlbVvfShDFBDDv9xnaKGb592LftUyoXbsUNE0H5Xz1nayx4vd86u3KhoHs
iyP0PtGlnBffRMQTr7w1scUDVGlmAnL6bfDaQw2lVOLmdBNs3PrK3rJtDrycnH8vOiqmVariqAQW
vcdkU0wBOnS50WR1alGs8eGPeUH3mExtXPryZPmlvHTbJPrXHeze8SGpwj4cXZIcCmd6A/EZbVde
UAtXvc42+ThBhhYQtox2hoyfTdxsjX1TvywTC/YLOCsL1NsoYYxDbVMmyd/Ec8I+ybR9V8WPMCRu
n29mEGWEw2N4eEHDtOjld0NLMVJmoArAFp4l3BkS3bx7doSn+juBazCCnfOXlZ33LMFJ+O/WOPme
04MDhgYAEKS+ltAPwccw3QHk3TAjVDx+hx8AczFRDIhsktXAMUWqXIEPR1AuIrrJD7OwZp5sN4KQ
FpD11ftBvO/LRmVLlNBRfMschjPywbdOqYcQ4PPkjrM93CyZ95546Y3qHyZIa1NvgS0lLdA7gT77
PyM4vLKz/Jso0vBlhcBQTU6wZGbp+o0wF9h9VAUJH+K7nlkmjwlekATLfemDFQ4oZV6bymV15U87
jKZCMQA9fBV5IIv+fAQSmFPJP7vkwjlWT5CJDrUP/MNEvSOv1EMKt1zKK7xKz1+0qcom4wNt8Bv0
iJ68PzUIdFlQZ7+XAN7LX1+EwPe27CjdKVXk+RnNsVwBrOrz0+5ZhDQ52NS3wj8r2/M2zT2yA4yp
lT14W0GQk52uoPKjCXt13Ct4zEydSOaUuAwMvLvXdn6ctrQw82EmLX4Eko+3K/SYzg8tXg8NcQPF
BelVofgmWHBJTUjBDUD9TzOwXI7UEIR2yz1Q6G77se4MBZnuU4TN+IkYNiM8Th7vS6pi15V04i2H
r3gSCmmZ0G8GSLRU5lFg1xlQ9S75Xj7JQR/0gxWzMo8SAguRC0K8GlLANb7MDjFsr7iuGTUoWCl7
vCuy5J8ONMe+ichsLsgrGnQXC+xMs800yhG+pwwpfXz1X+QgdTXAoF1LQQ7d5yK1lKe5MA0uy5jG
8Z/B6XRxsyZd70MAqpe00x4X+bKTE1a5ZTX//kEFuuQUKpsdw7ONrlLnkUJipOmSKojNw5P6awBB
kHqozIcnQOAraBl4kpKRA9oCrJtj0Cb89LU1pMLGLvnXAx2st7C9I9pMT9mWq6YjLbu5JRSlAMyV
41Td2Y4DUYxobtc8yYTAXN9DFgnmuvykEaHVlz1b3rDOJET4LuolGtTOpzArVQJb9s2vPyZaTPa+
6AysJVe+21JpZkZBpcy4ysS/5BhTCFjwonbUFwd2RMvoIbfDrOvuFD2bxZvQY6hHph1nBKdKupFE
yPtushYsbz6ekQQU44kOyuBNdfOPXxWDbycZbHn2PfO0ogY1A+suBRwxI2Npv2yyKgIvFipz7GDS
d/lzkUYU53Stb77ap/QFCEX9u0nx5eM9EIhtCah9MRobQLAe3Yb7doP2gd9O4UIrnrkfR7n2vyW6
P6b/3PbXuC93Z0oJZj+KU2Xh1wu+iNlu2ToTccNL3FfIE6T6SbDpnZ2lr35cANaPfdnfTIxOcAng
I5ZgKMvUvDiH+jUbZTIK3w/U3EXrh01b1zASG9Jl9i2cAPXAQFyAX+nAUzMKGc0Wl0UR/DeF8uVR
R5Dh7FcUucny3/xNGklGmmGwKPbnfOJtM0J3VEGiZBG0G4IATPBf98VdISdJ4AfUo4+2OAOXlPT4
n9mpdif7QPvL/NWLenj3S1zBkbnpjeXQrP7bWmdIxVCKHNQb4A2IRhlFFBac0ehKmlUnBvmi9baJ
gr2tvdVeQcib7quUGG/8w9sMJ/UyMH+lZMc0ettivCPVQ86+FKaJwjtBQB/vyyM8G2MGuwpB6D9O
ivv1ef1LG+yqmGUeYKQ9EeXI7n5H1oCXWThKVpPpYvBS/GQCzlTMsskQLCtq/oHSd+DZOu/f8Hab
eXOP9HdQmlW43p5SvZ1/DLOTuIyas3Ih84h/JKM+npuzSx/2Kz9sg9pd8iYmW85PvPoql5NmNICJ
aC6h3eug+STCsFkDncAgeHmO65CBYF+jOTfHAQsoO5y/9zNM6x57ZKobd4LRKRr5AN+b0aW7CEr9
ivGW9Fnc0iEKxdlMKf5F4pwrJ1+Ny9bzt6esG0+klpBJehSlJ/pynXlj6BRlEQ06F59rbpQoH8bq
ZH6XZDpAwzfAgcZ+w3Klp4ijK5qgNrO4lIL/U9Jt8ru0hzSOAJgUXRBkaBz4KOFyDyC/fxHLgCqK
HnzWdK++GfGcsKEK3sw4dvvMK7rV+zKKMLsrnicN7WAi7HzqZC694sFFLgiO4WKIencCapHJEHik
DKIbJ4LtX5nROZEKm1+dZ9AO1k/APyJAHall+q67DIY92bEXI0pWMfLncq3G7SvQ6FJK7ZtyBqtN
q6/Cu3LGU19ZzzN0zs2oJyz76aUXNjx8g4w/6tpddKAhDiF4bV5F0TLhaQmQPDt+atW8nbfu4Vmj
7uxlwLUNKGleFc+FiXWGQLk/UymObEETYPeUhE/FVmgfHUStilyyir/8fWR/6x4ma0VD72XfpkY8
mTCM4OXAuYvIqIYqTyqLUspLAMH6Ekwnl2Xqt2XUTCUGflokr+BP7+YetSn/nbSFs1JmaB9vey9K
qXTn7YBl/99SoHAA2cKX92MHT+JLTJQ0lXPDRuEabDKHQl/m6D/2RrkXFyFcYN/nIYLJAIWUGHt1
CHA82dpLC3/dzbbPwDZgsgcfJ3nv+A1P4TK9xDlkT5xnzgVMUNuKrYdaZJIRGWg9iBcoasV6uHA6
uJeAHYvZokhsqNYr/bB7mhe7cMK26tRXKFVefPr/EF+q8hurtGvcDEPs+Uy/wplkzZLCynpUnfc7
rCf4H6fx6ViMrP6/vn99VhKrdX1lnhCpAG4+AsoRpTBw0JHhkGDdvG9hgW0UOkgDHQZTZqNhqJ8Z
k99E8keaaxilRGI/LOJjYOTgiBaHa335DP9QeyLZ82jQ5LUCjHDfyFPf4SdDKPa/m9K0ule4vH06
QoMwGKYEKFOc13u+FBatzQlDCmQwprcayJ1yuI0SDiiWDIC8ALNKT4+rc9dbKgVUlmo8Wwm/5qQz
rvmjUFKW0FsVB+0RRria9Js9c4NM+WNp3xNhg70beN/4Loxde8UQxdpaW4ni+tQDhoFB3qOOgZwO
EU4c+xAFsHIQz/zuJEVIy1lluh5SSZ79EPhMbD8vVANc0hHPg1f0yJKJi1pHjh3IuQBJIs3QUguO
sOpsuhcvcwKlxqiqcrBoA0WnFyJ827OyzCa/tKcTXW4+20CWZsAtgNzmePl0YyBDmlvRmdYHP3fp
XLr8Yrvb3ejvDE6+tRXL84J8RFHRrekaCrar7YHjRv4IwqQBGYS3MwCQ5oIe/EXoNBAPngEO6A/c
rex6uqlhEpC67wldn6T27D9oKau137wOnu1zruPP+GLZig4YuMOG772Pm3Q0yvSXY1w7qeQ7fJwV
4gWZY7VxkEe41RMRQSoKtXpu1p/GD18ZSH7w2QhU5u5y/cN7gseLQdWJFOdnDY/0N3+KtwtnFaAK
FS9q+gQZp9GlHAe5YOItsbrSk9HTqQJKi+pVjYrlOono+dq6d23Wyutol71+tqVYAab0RUVJTQ7r
PH2TmAiz/tkXUb8U7YypgM8+cgLsWzU8xrG0dsDpDRv1lmFrGnyPuqst9gqTBzREBCUxLzyS3Kuz
tKOsi6ACrQ6HQp35VIDU3fXaSpdFRlQxrA3zv/UTTxCcnZiJE+WFQS6axDvQQBwSYVKklc9exAGp
lGecu7UzMpkVs8g5YJPNFnHCqh4QfCs8MWB47RFL5TPOdzO0WCmsRHqjn3y65Oce5pZe+UvirhM5
x3l7wgHJBNIPMu+DDXDwwlhueR55X/QlOXmkhpNdWxYZ5yLEsGNQNMt/CzOTjNMxhZgN8JxTsoCG
MqR2Uf3dsimNJ1eXHrXDcPhz0M0fRBUhXyzC+ezZMgQGU0FzsWfzCEt3mLshRzTU6UlqENxIHJiY
k1RGl5sKCE2gMXLBzMCg2qtY4ms90QVrH1JPHgv+Fr7+kdQLWHKg/V5411nhYTRuSzenHkP+XSNV
MEapaBPcPSNc717+fxxipF1I2MrwVWVrSdarJba5R4syNExluz+I4VXvgkvEM3jEqzh5ZnhLXwAB
+z/Qr5SbUbILcC64R5jRwyRX5mO1kvc9Wqeukl5wDjVfOwK5LANCtcXMl0svykhpL0MIgxC6zRD9
OFWLwRZhDDZPBDKkDCzK9d9nVudrz3B7a4fHZpG2YquA6FlZirf+DU8/C4LuUy14w4vN0gfULrI0
fXTmvR9KQkdtSalgGvaoGargBSJZYvE35RjVyZqUfH6iWtuaMCz7sZz6slJ+BJqkUfJac84rx1eS
sVkyT48Vec9J23G2jy7m/ezab6In5aAMdfmYbfOSU8pEnrNYg3qHNgDSYZObEKjGUK7ghK+S7Mn9
bvM84d+IDwO0lsV9BIQs75Ic4ck0TPVmKD73xqY91NPmJspodRzlsXjGzUyThH6/JLDH+JGR9lJx
FmyotbnlrWL4KlsjZwzgJugVwaRRY7OQLznzYH7CzkLQ+DzLFYfdpWNxA1LQWZKkvw8zQvzyNaj9
Wd2IZVjXm8qUsQrH6XWfSHhFsUMj6E5zJq40GaE11qBYXN0vkQma5WnQXEBF6SfCDORsjX3htN0L
IGiKnVsrNOfypR0VQg6nWPWViEc+q3A+uuHN8Z3kjhXfLbZYEzGn/H0eQY/hVkmoE8Lag+cqwXda
UNUTy22RlesTstarsYOQ7f6VyVHUvk9qepDd2A7idurC6SXEVpqtjNT0gmuSGtO2/A3jFmXKQHB8
1yOwJhG10bypP5sey7aNroeW8ctrU4igqn4rsNoOBW/BeECOilPHqZb2pbcBNcw3InShgVIY+5mA
Oq74G0Tlzu5zl5xtepU77ShruagckDXKMTJzUkoPMbX0/Q9v3kKE/iR95YsvZazde8S+VB6N98Yh
LSkmuyphcvSo1T6PwJZL0xrsIzBlhvvpOoOm4CPbZukCtBKAR3jfV4LVbgdwvAdgkOkRwqUTzFNq
0KJvnRdvQ/lfNl6V8M4xdj5if8JGTkOmlvfIqNBRVrtTfYwQNvjUcdwZ+fc+UmsVodOdWFvCjGgD
1s/THKsx9YyN0T+kHVvu5mHm2x6SPZTqi4xRkj2nzscv+grF+LPz44IOAoFwWu04asaUiw4JPQOz
5b59PITojgmI2cxJNQqfqwQfEe5IY67dvfSr1y8Di1RSTK3+VgCbgKUtVGNBa6HffnQHMCQYxkgv
p60O/tJ+nKz37Pp7MdhZZ2i2FNzaur3HAXcLU0qYt6WmlUMlxtP4etFEKOt6u6XaCDBnX7TzCLLn
Is1gyi3fY/H/i+f2tRuJkbOclgWtgc5jvXgmQAOL8G3ECboQqWhbWc7abzwrWBHf+kG/hIjitlqB
8+Mfl0Ya3h379nEZK7Gqk9Wu0JmDFBSVfJDZCoixHgjUeoHjwERfhmydwy3deywW98K8BjtU0Ghg
5KWopconI265iJn9asR2853xI2/8oabOyH1RSCrC/KhYywkwRmDGK+8Nq69grvxeo2wXCZ17HOxS
/PzIQWhlCc4P/gGq9chrjWV5jJ6I5Dji56derQP0OuSd9zAEz/23/XFEG385LQjbAcEof5cqSNc4
9Xah4wemX2YY33mWK7CcrSaJ2/D89LSljEgwFVJePLfn5bkblQmCX2xM+ohmbqEn4QcAFE+mGrJi
8OwAuHdLzFkRWVhE01Z11WJYN6qZg17tNmwQLuD9FrN4BkZFZC2Le36P8KmD4XcHs9mSStdAdVWA
7hWdhS8BKl+C9Pk7kn0ciz+wzWv6I15mCS7GIB4P8wnZ/WM1Mkiv/gWDTl2vZSoboAy3XSeMi9+O
pVP+e/672OCHMAMehKRD4DXcV3OH7CmvTiJsrfJLWBwqGxdIZ8UbjMqoaIdkOFUHExF4bPXLsG0i
zoAJFK5wTILaN2y9R+/VSb3IueeMo9yuDYLBMdFjz/LByhTCKWt9VgvC0EssIlRz1xHH5NmMlYcc
vd2XYaP9PQ8FvpeEcpmM+jOXKlOmCyOryIK1vqXpKkvxH7LvMcJTEsFEiorBHBS/DC5ePse+qaw6
Wwz0h4RKEvIM4jrniz3rS2Ncpd5Ws5++U/ta3Hz6Hlkmg6/FFKX7s9pBWXAw2qt2pzmdndrHTBjO
9nt6ldAdIbDNB39EThVL7yJA9T52Owj/6f0SD+Hf1LePvuM3m1fqNqkJVhEHLWRmOh55I46FSwlx
rIjofK7o6+d0p0tK/D5pSFjDF1AcM4CW5nBDbWeDre1ZkmTPm1cgm80S95qwDu+WZJEt9rVaMfkm
HQy7YC8ykiPZ9ID0qMzFSoXcnhY8eYvNas10eH5dinkYMBibfOEU3gSg+OiB7msOxLkDPcnp0IWR
UuVNAwhAgsh8MxB+fabgws0fTPD/EWdHHdMhp8PK8Y4TNTC91Yno9NrXS9dQE1du6LzK7jOyveBz
iD+W1as7pj5+zKC9wX/cr6NHwKnBIT3oTojhVIb7lHjdaWGXlv+ciODp6kTDD26gvyHxcnjSDetO
rvltF1a07Z56QMJC1BWElG6han9kHIZpU5NDLjoyRmeZD2yHnxf49V2f9aTiQDUZdeIdgzrG618x
L7ZvHpmJMiQlMnqKRvDFSdxJ605Pe4RZhfAZ6tujz7XZ0bAfCBKyCP3ULPWjBa80BOiv/eEm2RSj
bYxPmX40VnDQvuT9bYK+tckttwTeTAgif463HkgwbPxb0DhJcPGdqEkR6zm8YQJbEJKObCwbz4dA
PiqgGKXdhHEYjPLdMicNWEoGW7TPoJwQSrb5BbwXI37g3XbW+pxE+P/GC3P3m5bOMa3zEI3cHvr8
gwDSuBhF2ifGzEpHlF2rvsuX7EvERPDfeY67Zr42CWRrCYf702OWvo4pS43GrdK4rVoJ1iRhM08O
M8DldFZC9hPfVxKQIh1IBkz0eA6WmizimT2iWg0ZTNCVNfcTASnihjmVQNE96aSbGnMI1JRrzUzc
pA2nwf9TPp9msSNU/0TbwL5LqU8Bb3N8i1bC4WFhul4MO1/0SMoAdJqIRsN8fqg+w8StohDU6J+b
joT4C0X0BlCo1aDCI9M8K27J1kf9eAQ2dQIqQLWfu3JJpn/nr6w7fMlb1UEg4EmxaOwoFE9HOjfJ
9a1NQdW61eP4SGOyB6SnT5FbqLUANXDaIH5Vz0j4bQHROnLLK9ogFoL3okdX86crgovWg/bYEGn+
AIJ9lr3aEHZf3UAzDXwkiqq+E4FoLJUMRZGegPtPdkH5Pp7T/MtQfLPNceRsROILXjNpwam2Cp66
CsfwW/NbEBB4ATIiTyMQ7nzUqREu1QANA+mwoznqYxsfoV9zKli2Ri8/EdBuKm0NQe+lk1s/qYXV
1+W5GVwG6pQTC5NTgFzLKGb3AU1sUxEL1wane0XmHKXSZcC5vP30GWn9d4L52N3vyUoTrR2Avzhq
f6+NB/c2I5KPKtUHKaEg5DaG+q2EZ5JT0Yz7Dv8QjdcbHqvnc4/Qc+2SWIIFT7SycxWhvdQ/t7dR
x2ULOxQCK7w7u7t+gq4dggev5/aa6HEH6TaJ0abDx+VOlhVvfl89QpXy7vMoc8ZCuNloYuke9VZ+
9WjmQqsGLwGG0Tzd2T2e30AITnl4tKsrFpdsjUAYEN/wbTOgq5M0VtgBfGVrAcQQig5nxwe9isHe
KantEY3LO/f/CfPG1+Fv0C3r9nHa/IQJvtaKB1Kh2wIcyT7+ELwmvSIueX+MLrtC7evAdZGKf+vc
ExR4aAdkKvu482D8xQYza/eJBTbWwosYYUwIPCR59QYxq1KAw9Rm0jjwMMU3R+sLqRA2p/Ll0p+w
z2CRNHlEi0eem9vXcsVs8dkBJazga/4Dx//IkOAfzjW1r0UMdUrPrs0e13DfSYlb8QnI/AkzM3J9
TV5fc5WeDQ/dOqO/E4tkNuCM4wQ2iW8cPbWP9wnLW6iCVljbki3/usNuLm8li/3EiwEKyhDQ/Kpa
zbRwN3ONJPedzpEhxFJkTrBCLEz6nXjztHULM5+/Rv3BJVooSyU8EyWTEqPzu+RixyLRQGDV9GMp
2HFs9oPcpZEqXAdJOP16BmQI6Ez7Jp+EThkMwc7AbTV2Ibv9vNQXVe257majlHwCZMJz3Rbpfo4d
BDwyXDZd3Vg+kw/bvQ4K0GVB5YFBR/hI3+PDHQZYJxgY0vNWEFcbQ0ZiHWA0uNtWsi0JpZXBYU/z
cdSrJ6pJLZ73Gef/jUz7dDQFakHKGA8wVJEXVUm7ktep6wrZIOFkyRce0wsQhlExTepNwq/BMn/9
Uudtwn1fzNC0Nc4jjdmQp2RyNbU9RKT0TBpsVB0fyQ1uadJmMZTkZ8PMIYscHqyAmXhHrGw5d/Ig
y+i5iMUiaQQV9edwN/8tZSiekGKce459bD3T3UXzr0bth+3QmiAJ+/xOaNulHL+urcsPnaFL7s+f
MzZZ4JH050erna0JMcomm0NHBEM02yAvKVxoTKDf/RwpdASeQ+YGYn+Ctfq22JIMehBIhF+BqCED
01Rh98TAWRqIx4tc33kaiNw8cDW5/h8ajYeZxAuwpiuEqOsWifvlGESgE13/vtbsvFhWXxMMamIr
D4pKN1pRSfrxwoln/6l0Hwc2V5/oOgbM/FpNOstL0QLQGtvFPCLPV2J6xH4q58dwAlqRPtOAFqW9
fJc/U9E9Jgc1tyLEr3oETzYUW5tza++bTW8OIHU/0jVg1Ue5tc/ZJGFt19bhr63blFzrwjL4EEag
M7IioXPnq+khatOBqbCK3yOMFwYvnS+FJZIhGrD5IG/+6KsIsMuRndMKLAbA4dRtqz8+146gS03q
1Gctjzkl0ohdvv7++z9H7t0Q2OHrdFLVXwXfyMbRYsFpZpneqmdFOCT0z85OsXVgv7VHU3HkQumN
LO3yjblCmjPDFGcfwKcjVslVPaLBa/SXWAcWQbzz6xmIpcUc7l3tfL5qEhA61j85pCqIC3TiRNmZ
0Y/lA4DkQIQyT35wPT0XT4RZxiAMo6lhjGmawTu/ZEdObDVDPDV9kCXBlOJ1NXqPOx4v+GvsTF9n
vvp6bvm5H35x2EBWV0N3n1ktFPToZou9Tsjch6FjViJrqIz0G1LDgtjnVFk+qZH5ZxaOQbPOu7ra
uT01Cs2w8saAuZFYMoRYIAO8todmg14oaxC4HzZfKAHtwtPUKz7gYDQ+Wy1GjqjdznGIZjVJKTva
aWeGnJjhXxJ852N/oPEVpxi30OSbWDVIGhAn7LaHKe4fg8fbJmgT7PzjoCrAHQtjuZpuLUiDVChr
4eZa+xrVJamDe34eJ5sh0py1z/9sihZZpagBKH8hrcD1KuyCrpqZo+Lqlc7FZh5qUdPKQEQ19oxr
k/n4kF/JefDarmUVDGACw4d5t/cQakrFKLHVYjKqQvLL4YcWrvxpwkxb5RSdCxGrUl/nfP5ip9jq
kaFgSNsX6iakB9Gu2jEkT4k82mcMutWOLNBmjZgna+qetlhc4uBWj64G/Gn8EsA7+dFHMIilMXY6
HO2L66lQUMXE3vxmfaXL1P0kbgKIQ4tK7reWjmVHvcFdX4CImros8ai0WUPmiZMniPrVeykvR9tc
VW9Vkw2hY3gn9XwNoF1Z1NxDqfqIOZI+dakiWu67kyTlFY/6DppucPbgV8fP/6jXZQ/gswFGHqDn
uIWx58+JWXLJUqtmUIwL4pD0Srn86XudJxzHicfVa2tAc/38y4FENbbyb/Ert8WXDgXgrnDc07Ky
9DcGvOBwnMX2hgFDBq7qBAuCYhJNf1JzFwJn4FPRQtPCK9SYDac/pT/4aUTV8CTGdRXdvETr1nt3
qq33lJ6mJHPZWbm3hZP8Y/NAyDFOltPBB5mM/AC8ASxu3UJJGifdTI1rAmCjeyaJH31ZS7LsTpg9
AboI+B5NYWF2RrdFB1I/KSbjXtQfb4DzukZ5LCkY4ZkJOx5kkwWX90jO+WxNqbiwK7bI0vEfzYoH
QXSoSOZw00lpn2TecTchrVBvpKMqdXW0m2s7vxsOddRtTvAvarUi9pRnMNnApUTexp+NZh1WvPHi
f+jeMKbwUcTsBhq0qv1G36EwlrM8FKPCrJohQLaXgbHUJO7Z8S24X5YGc8gyJfqlKKxjZqsMBuDg
KL0GXkODZj/cI9wPy1mo7TQ+U/ixfaEYkPufrQeQzyq8QY79kudAuw6bnhIAfZ1Jx+dqUINSROKs
KAUiE6X8Rp4Wej7txzgO9i2c6GADbdFr41SUiDW3rbZQyQXZs+gjWbKPKzRJy9b2OzyIDVkh6B3p
6HGgAR0r+vjUuSj/UqqhGEqoTuHl3YlUZ0u9Eewk3dWUiCJN9VxnOUInWYCjel6NitffBH66M5Jf
b2SKlr84dfpui+LDomoYmCfrH53BPp3ckH+M7eBkfwdnynrvpXSEpPj+Cxotvyfqo8+3FMTL3X5c
lW0//3+XKtJSnD9ahDoF6pLSDthOhQsc5LCC62lL7BJVRld+XWrZOjHPQmfzia6AJR30IqHLGBL3
4Rvu5TcCqROA+RsY/QKhatrGNHakctmNQYAee5Mstfg9FJO1FfQVSQhwaSyGhuO08Oy2tjHXQ5e1
5lKLlkG6O5fQXL7liMwbig/JBnzSOy5hLYshYRNm2aFw/HbP8xQFa87wIUBtDSjBYaAUtat+/edq
bCXyhC+xhvKCa+nYEcciwyBf1D0hx1OFZJhYEEHwS3SGL6rsb1ha3gchvEk+uxtjhgwOJnVKxDix
bngeVURnxT/YvxhpJa8Fc7gR7Lx9iH/+YQmte0TXeVj5v8+7qvnW2h4beLeorxv8B1QHUzbNNaLh
m1ekBbJos8DGuO/T8XxVvvZ4iNYQWZJ53rNNSpSIHKSYgbv07mB42YbXEsuOlUp/ixKpev/1hbGD
cRIqHy1zDWarZ8eStiRskQudFcePV2b8x81eXgs7RPravX5DBbF2aJIiUrYm6cxcM8Fcq/5EQaZP
amNcXbWjEiF0mUGGRFAS34WhvYtWmec9T2ufMpXdpipfqDApNsWJ4Z/uxY3j76Ki4APw5VDwGTrd
OsHw3g5C2shYSTGxUI8eiSdRd77Nnwwh9+f9c3BcmQR6aa/UKPrV/avmZig2FGWujYrwodyjNtx/
HK4djFlki0QsOo0/DbNp3bQlSXeUq8kszGrJ9eK0dfD8bErdSKZOD4+RnfL/3K160HhdY2u0TVOR
PakVHesqOYBLnElM6AGcaWuNsxQsOjbjqGl0q7l/2x2t3mBKJwd8QIaQ+585LtSQlormAYGUAH77
Walxt5QkeEIgaaS//LLkGkULLM4GbtmnNbDeIttfDVwEWYqNTsgbWHxTVM2w1ajjC+dJ4VWYkU/P
caYyzd5v5rKzwTWLw0linDM7h6bAFibEZ51G/AVVq+WPkNpxDGjQShdHW3T1SC5VxaKoCfhXxKSH
1Sle5Z/TAZqOpJGfs7fMsaX0D17Ep4TFQrLcJBR7Qi/fYJ5qLsBRi0p9l4y6afv/d01jtDSlrJPp
NmLsMGWfAvsZZcPl63mVbgs9RXi1Df1mqY7TouQTNK2Fm28FSYwsIDxyo11Rx/Y94VuHzA9YBfFv
VzeGzG+uKHX3SVl423//DnYXaFKghBb5Vc0fCBZYPKWvl0Yl5J6WAITPevvWjIec5hZDTNfHxqwF
cnRBLH7NDlcgZlX2ZcamIH8mEFeque1h0ypLYUjju81rG0kN01P7qdvyyzOarIwFDj/MqZXIy3Wt
Enl2xV3kvQRViHWgsha7BhF3RKZWm2kmE+DpGrOYGOvvViujmzFD3XdqOXAMlsGi99f/yp1xGWtD
t3HmoBna3lu1MlorNV/YeJ9TXStvr5t3BmSn+w6GbPaxcLwvNmh1XiOu1svEIEHQY4D6/yv7JugF
JAkOc+gN4cFUMhrY30s/ds7qQH2J1tTMb+qQRKk4xGxe4FK4dVCYwYyxp8cm+QRdvAacdhqNq/j3
RyVOUv9bf+O+c71PvQSXVzD7nFsraDEXk8eWMVaCBAsqhlzJkbMaT7PEwnOb4bHMssvsPL0xYRfQ
rEQW+LwQKBM1XoWrWAYt2uGHA0C/9LRsUfv9BdVFzWaSdVUL+IpaJjutp/euH8R0XCgRt05US/pX
hO9oNQ832b71lcMOoBQma9s8Lyk4pXT7nFnzALGvKfgdToGnjSMx3ph8OG3fr8ITxKjQLe570oo8
+82+KOWPDyXx+IMt6l1ZfnvIuC9Qeu0RPhm/5hQirWvQ0iEVuG4b2iRwLvMEXoWsfMul/4WAWNiG
i/ITZwQ2fSEizU9xbULvVyWVTsst4jfoC8KQGnyD0hOtO1qqvdfFhy1D5o1q69frA6lS5gH7aBWD
2+MTXXRiaYJjUCabaPQk5wUFnAnkgbraQN4UNYMYsdJyL0IKI2V4nRDZ+YE0nuioDs8lki0IqChz
zs7rpajiQf1j6Dn92hj5MF+dwuib4J9JqZCJ9xaeU4Lv9rLkAyTUZBdaBInrqoajtNtZ/SIwsEwr
qpEvsJWh11g0xkdDtBaH3NOtZB7lnWcAXoS9yiw1TM4n8TV8i6FszFk58vMF7lweXl8RpwvU1gGS
WWOvJ2H38INW4yXohW6t4PgyfG7Ibh8p6/vVO7L3TqdCONQxmhFU6YBA13PgjfcCo7OQZHG07XLF
GJ6zpiI+En+CAoFcI4YWLrwnifyEACNW4msREDgUXOltZBdJDnFdH4qtMeM1Ek7CLvruPpCED3QT
sYK9aUsKGTe5tuhR4OFJ1O4DJffJtLVgPUH31WzRnJyWYI6j6Ddw/wv5WgLKtE+vXLFcs0BbPXGe
q3vvkC4owSdMHGeuz6DTWdwbgNR2pz6iS5FCxZ5TZahezFry1QB4sgxMnc4b0ZwdtNcW1m8w2kZQ
7whBtG2d7vg5yyKiSCV+Xll8YSHp/1ZkEcMFEPn/sRO6nh8i32XksnBmS2qhXewdZtW165g6+W9P
Q9tpqYcr/gBQtn/VFy4o8D/7QCSBtEJnoi/pKXRCJcJV6osA9D/0UGFbhRp/6e6TzFKmNHBL2PGt
cf93/vXD5USDZVU0ncCt1+RK0Pkhrf7oZkhtQqkRNTDggWofhnenoMh+QJBz2c3Qax5HpeZEwbvr
EpL059haM/u2CBcJRKaMr/1xS1YoVM/3cqlCVY/iGwpZ1BGx7J5hAdrC3IiVtiH4wZtM0qj9RW/J
3BJPX0brqhuYg/w/BPsbnyju4URW0DZBDbidn0m20iC8nZnFT7OmKuTqQsqZMR85a+dJ3Hwrjh9E
4zPr3ROefN9edpzvifD9X9RRhjw69E3PS6X5C5IbUn80qXK5kzgTFS9QsmHrvHPUMj+Clk/bR3MG
s2WAP/mUoSrIc2jqGEJFosenqiAft82COnaZmJtaZZHBvR54ib/126rF0+/F6OeRMzgWfXBkhwQy
1xdbvQKaWwCWMuxTAFHM3LYAeu6y9uEJqOa8uAlk2V3AZbXGuzlUj8GMDOpA18I+wzaW69WvBKqc
VrDGLkGG+G70VaAa1cGoswPDAxcCd3K8yr3+ytO6xFjo7kWVKnLEybdZT+R8phheIG4ihE/FAsUL
F5hr0uFcaxAOPVa0UcWxCfA9sTydnMepCHq1gDzh7zY6eVU3UXh3YsBCKq5zKWXIQDSnyxu/bT4i
pAoe2isTV+3wXaDwacve2tduQRDvwIxTIgEnQWNR4Oaht7r+HLMsHdhwFIqlzbozIqqfrmXOFZ4u
WqdNkT18v3ounpcrlOSVBLDLYMEBf1b12ei/UbIXAg+4hwU5pybFD/hloOiascb1nlvEdkZXbNUg
lgw3vlb5aIFCKThdlJCAG3djAbp4oYPIVtEKcUPx+9k7kydX5M2QajWDhtEhBCMUgo0yh53Z9BEA
K3k0q6gU3i8ddUin3iN4o6Y6Mi1KKoFKYKEvEAlCM7lsl+28KPw6DyeRxqcsX5swErlXvAVAbSue
wjHfmQukgaDxhiMBO/S23iLZ+vjqn7y/yqIZhRydH4tMbnIqaDaSGfdwgK/Oo47K4+zELSx4OvP2
tkK7JPUlK3jEtTyxY4MHULLr0K6qpTUMB557BoHFnNWmattYie+dymjPi/1ykRIsG3zhaBygo8w4
BDa3c6OkJoLngaLtGPDERb9y3RE7vsRy6VaBLamRtYhTS/YS2OZUeRzlCB7FLFg4tXuK+cDfwTLj
MH2SKsp1vwVW/gAVhzEHZOlPuNAAjgzSaZeRJ/VoVRcOh6WCMpRL17PH5ZpmPl/EVOQJbf9oKLXE
UM87TeQnfEYeqNaHi9fjepnakX3TcI1724jC/Do4JZcmBY1t92KcABTb5t442eWUaHHfCkhq932p
eN1v92QRijTyx6XeYW9U2shuUezSPkbUppFKHiDIiK7MxWbM3ymuuWIdqBMtft8GtW49lIwrtSXx
UoQXiHgttNcOGg4cCFZ8eydIyw3e9cdQixCj/wQi8ii3T7S6RNM2IhXGd09yU9P+0ybp0p//VxyU
gZNyTQzS9/zPkQ2Tm2rZ7Ns2UdzXnpJEwFWrHFybGy+MUWPcW7uhdtrmjiSAle21h+/25k1mt2Zp
ilFn8ptg9zsFhQtEUmDoqlIs/Ul00jLFjHEKxg5PHunwHvKTNDl+eu7xyx3Kdhcnt/k4MVD5Zd5w
Rh6pdsZr4esfXRF2oiIpkjz32OfjbmtHeRSSiq3soDwrvGQXRpSCHSnzwYlu+vqQ3JiLKsCIRx+v
I0Qb/+NKNzkWgw9ghS+HfTjLcUU+/HZIrVLvg9NzzyN2df3cdE+G2GrkJIC5nVWOehnxhFStiAk4
bMr0C5y5cSiDRXYvtPo5ecZ1en3PoUAwrsob16GKZxAapaSSHlceM4GM6EZKCsPlYKTI9hMmg4Gg
0nvST/xJskdiObb6faLKo+oe+nqIJYP1nnGXCQ3qxPxFK/3ZbOw4VfmodabgB9pH0hmXK1WxsfBn
HnJWE8uNywXLNJmuKM5LfbxgPHYgLZs52eggxo3SV5zy+7wOtwn94dwfaLB7fS2Wu818FWeQ1rqB
f6KSYvXe6d1M8YndQeIJ99PuggyOoxRR0+Lusfr9TgJIDhS2Nlyud2tV3JHhVNHqAMNjyMQjsCyD
PmYOLTfGmbjDOsKzE8vu6HUknVv+Sjy0d0lN9DdOlkQ170KmRkB9oONPDzTylpsc5GL9Ju1TWfP8
uvrsNpaNnWYURQp10g56FiN+4aCh1jpmlqq7caSHepF9XR+P3VyCe+gJpkQVLZxwGtKz+ZDQBSj2
/MMllJDBTvQmgxMQLLmCX2YSUwBOwZ4G9CFx59iPxTgAt0UDk0FqFBEJpA3tOULINoz5lRZqT3fv
EFrMkDFc2rYDyXYmMxhSvRwqZWS44dbUC75tds8P2MjODZenNC4vMDYi1ubS71J4iJnfLJT0JZIR
fK94pbayI+1wmF2XTYKzGJ7zNzJFSO17yQh9pPjX0L+6rHF786wTIGdMeiwCg5XFImf6lyXQLW+6
USUyu1undhnaThZK5m1pl4qsqZVFIO5YKkh/zv8mPmm+LndnMvMSpj9qzKq3o2tFaLyLPHeO4u/m
GhfAsthswC8WYixRimHZcUqecgTP7v1bZw6AAgx3gptGGKQrdLgcRdtBlXWY+3x2moJgOlpGk17o
qcCJYg6516CdQQHP4L03bzxgN0Etx9wydIrv50O0VVEPnWN34QEAsKAxxgNnu3BggkM9ye6ecY5W
9AWYtZAKepZudRcYgfUjISzhtxJdmlHHg8SmfsZuJYELiAQaei483wwQNjmbSevi/iVMFEgXG6m7
z/96I/3SyCgU4orl0K3d9eJog5mF2HOShyzeBfwJoWpx1bvQPWK/NxQQ4L47QeToOfTg+LkgD8QY
+ORpYlvIdGTMzJEuahme48xk9RD66s9gYULlW9G+3DgZ/vW2thbVPNi6DxXGsdOJt5tmXzOzcA9P
9HkeU0QKd/19TtjxuHWESVoIIqxNV4dN7GXlaxDdRYTtsgwGKFyr2qLS21SR1gBwjI0OQ56ICuws
cG7ltsU3GUCo2d8q5iIuBOhgjucWIusuDVd2reIMbtq9Snd0uNScbKxLW2UbKYQUlzmJuWdWG6i5
rveRk4jLp/TouyOSgp7CXKfp07+UBdGnfxpX2zyGJ+QWuvnkRHgxb3EKlOeRwCek/URDRZY3usqL
a9zhcoPbFQ4BSLBtc8jE6mUUtq+fbpdgsgWDKAboxssJPTSuhh3zpJZw8uyEgoOQgwgdOt2kRb5G
/AKSDhOIC89/h+P0Q6fEetPSZRevjfq7swOsIWDoZlTePRsXrgZJGf3QTWGD6DdeDNQPHTeNNowt
spT1RjoMYsfIZofX9l35NcA/J12jLhAcZlwnmHoiBP5IJecYBIy9hNUXZKlspZDDHUZ0iVNgv1R0
7EqZEM4Kd9uS1OhZvB/6XlKfTT6ukd5EHvPrcOMv3oN4Z+9C5XzVCjzsCk+//SPAlGFkJROCBsaU
FCCmuSTXxTEETIV1TqI5PU6FSQYetJP5aNgBzZWT6joxYwJujJAlQNRSXK95Iteu0uzMj0eZ7YRx
gHvYZ000TU3XdxYgjy/CXRmhaiFJQhKbhofXS6LISQ6lIY1XwQqtQ6cUG7etcrmORtBmKUWovadx
cf6F1caj6UgqGq1T0JXa1oJlx5jyCAmCM/OzvROQY4q6KE+xaPS7c8FzxjgLyb7qzgyc24+u/wGL
qyVEZlSkvVlq4QS66K91jdW+HkMckXz/iQUDvSfd6PvaId9uygPAmRlwor8PqTwJ087+ZYKwMraF
7VE9HdGy7/M1DM5TrVTcqwNq50YPFdKAppAlWbPQqFZwR+gLbgK912ye8M6Hf0tivrIyi7sDCXyp
PjczHivPIQB3su/cXcBAEVkJbu7bWD6phGBq22ULtgae5eoodQnvLTwCkoUmcUb3c7WizkfcfuJb
GTBsxOxdQ/q3ARCWKfuWuZcAsR+sx5b7aiW+nFbGzBPahNwlYcmoVIIKK5DOwuP6WU3C4ZF0nh/T
Z5xD1dYLwP3dRmohsSxRTaqthXw7+lLt7D8+SBLMk7wqbhvKoVGzVIpYt3LRoUF60E4zOqs0djbG
TksHl2wc+Ur1bQcITIpSuIZatt/MEyoVHJquLoMFmAaSWH4TNbHNs/dBjhgIN3vo2ji32YsmE3df
HZn6fM0zwB1qXST0geBqX0dT8VOt/mt4mjhFtm0xhiULb8DEU9ocv2EFj5Mk08dn+wxhqkZiZx0x
v/zkIza4jBmVPB3DZorx9ciipAhGH8Feow78tj3q37BkGpHS0MrU4NJbSaMgoQdbNsjYi5piPqU2
8J1hklTJpd4wCpkbOi77MmBJ55OfSzx2vJvD67+e1LrIiO47gYr9CroYFUqRU9Iu0a2TF0qx6CwW
/WBrpVMsy3Fp6L4vmtRQju2XsgD58tv/zU1yBfmYD4jjxZ/9R4zQmhCkD9RnDgNssiLHUsoTUgsc
1Y0wq6ysftJZQArT4R1Rig80x3MVXi3JsWq/1cOaqN4CigsNNuQiUjemFAbEpVhI4Nc4E0Lc0KDZ
Cv13L46sLY+nvnSqSFXA+W0ozsZL49c10TAuBlmkbhBmyAS9uVW+LtdtLnjAyThAEC0Yp0dHCRos
CBxjW7XXKPzuj6fBBjGhRSPohO8PcKf3H8V2l9P+1K3k6q76UpRmbAuu1Gu4uPQnP7ZiCF3S7Zjq
Jlwgdr9VLaWxzzls3DpnngLmIxSSjhIV7Z+kL9cg0NbiAd8ibzxkwWrf3QAu+KHpnTA9hxKDaq60
yyrOgkKGd8jbm/3GtaDME+DwPeCUimdRd3Y04W30pJvawWi/V3v+rh0PO24sPRI1Gpk/RY7hjvzi
0/VvLtIgkJNscZhgF1e/8nslGHntGwZy5mVvrIRjEXlhoCDh+NaUtcbCS7gpaPr4C1juR0wCcwOf
aWP/ArC7RaXiS6U0ovznT403KIFLCQ6TIghuRxi+p426RK70MiSiWuveWaBbZeM8a7soOzLG3+2Y
OY/OD6TljuLzvjosI4pnWr5z81vWdOLKiYD2oDVHfC1uYTzorq/BAZnzvrkaltYqLumf8Oa7Sh/F
L7rh/8vD8fEevgymQmWadVAvA6ffZj8COd7xaPkFLPaM+XASkgUDAv2k0spIj8ZdUQC1dz4lAWow
/c/RlJxuJc6K/Coui66gNO4fzLxVYUFQ0+vnC05e9iEPiaYyPsLgg7j5ZBrkMqUGdxbmRczx2QiV
JOdmFGbW4bOyNZw2lrNlPjjF1MhPOyHzVjaQSc8rcErGRJl3CS3QjYcCUqu3hxFx5/3VOFV0wqv4
cAWoEUld6BpPUBzaJDhqscZRAwNNk/Wl2F3TnqiPIH0wj7JwpaW+TEuA5YuFREg5gzzmUQ5YmnP3
S3d2siHKiuDhjB1M3US6ss6+2FjTtzK12mf1fMY38U0ZJ2u9hCk0oLCW4ZJXub/Qh1FL40SHqJRe
xKbnDsqZfHz26dK2ePldPuLW26VaJ9V5APv2mRXalFnkWe09k2t5T5olCLV/8Kxdd+3wf84AaR+m
F2+DZGhdFwfkjTBBorSZnnxL8Bd9TsHQceguVvnFfkld3cwuas6eZ2eJ1Bu5kqqPQitHXQ1+PsO0
jA4EDzyg9DFyYFW5YbGjDBdm7Y259tgHJhmhFwQ8tltJoFKrff2iOXqlHX/UFqVjaIa4eRXb0Ff8
DlwemazOelAjoVgsTMEJZ2nDLLV70/pi+IvkBQXwvzpsqyBA2CQ2tJwnWwhrPnjiZO44cpKiI+v5
nl+4CkacTYbZpdIi0ABCPIM9QJoQpWrB7HkQ8xJKDShU+A4go2H+VR8ItJHByfTD3263xzyJ/ecN
TmEVCMHCGLthZslr3+2Bv6R0D2nOkqy/KzVyN2V36AcD6unDIYn0WiUnMIrw/TXCawJxH/qD2aa1
SwJWRlK9QO7TNkpHV2RGa2BjFNDlCwGf5JZcB1DT9vs6akhoEu/pE5RJ0ZJoPROpd/ElfwxLeJ74
gfLfRwkwI9+jlPSLhint/Au3+UVhB4gREgfEcDgDVy0vkqrPrs3wgpJjL17Jo0uwUeq9YvM6YYDT
ttulrxIBvqb2QmwpRGnxuECH5PBz3vSNa4l4XY1IVY+ZH113vcH8Lr9q4HBOAESo6Y/ZI6Yvt3FC
xlp17olo7qKTfyeCxh0oiwNEitFQ23IxWgBpXmlaFosra4UX9copN9v8EeJipgO/0DMqAiWTvbdl
/XD9LVoafG4mPabsFqEOqZDtCW8ZtnfB3fbOrJtJaUtxIU+KaadhYig0JpeRteqjCVRHBdt199Gh
295X0H7gzvnUSNdC9x+8Yl0uWDSiCfv71sDBMcIPS3oQmBkmry2cOCYdPZhqc7cJ+UwQIT11kCYo
i3jfHUv0ms/d5GGKNOJAfVm3UQiJtz6+hazo98V6YmROKnRGysr3dddF5z8LDu5VOPpNGgOSN+1V
G07+OrPuZOO1G3Hb4vYQkUMR23Ywn8MvyLYtANHlsWWCpKhTxgZZx1Bz9uouuSkb4OBB8pCW8D3H
aLbNF8LQ54epG4Xisikqi48fHxxDo01dLB0YKyq+tbCFIx25LSk1+OhdXc/2Yqy3rgQDcYNlNqOZ
F9a9r2UxWLvzV3Zwr1POJnJYUozk4+yQGt+TCWjEn/WJ3+agZL7dmE4EqyUbL7eBs2HGEqbL/vCc
Rl5ql3yUn0BdPVLzFjBmNoP8c+U0tG1xXz76yHuGdbKOwtLk7nxaxJNOlAaI7p7mnenXZ1yNkhdF
YbJGKIpgvC3XFN8CXZuTHRDMCTAIIBSijhWz9GPk9FHSZbp0JFxrJ4JcDPrMfmnQUdIxEb8bItxt
agY/4DRkCwxzT5C9W4elcXS+/DzrZeQvtareq4iIA7qvw/4DwlwGT/fy4ynAvtzJoFrEyL+/GPE1
xZNi8zX0gazMaVGccgnMjQS0eAbj98qXJmM59ONGtvnBprDqSMbmrdq3eau2spwOaADn9oV/lOsf
tmjOmB5C5Sv8OPr5dewdIpMUDsZeR2y3kzg0wtMtD//c4zSc/8ZBy9KOFordRoi3N9nkaiBQqqX9
owF/SCUTJouSRPprq1KVPyNUXLLTzrbJK7+y1v8bFvrSjeGkVyfRpayaZ5OtB9GopNc/OdrzY7YM
/15H2FN+mQoMCj5w0YjdNE8FybInc0AejSTImQT5lA6uhbqhsdrP5yIhg8rihzYY+VefM1kmbws+
oMhg47wYK/zKylzvNp0EQU8VKiLfKnj556szcf9JQinSrJF8U1wGUTZp0hCImpcJxtdHivgzM8b7
QSLuSE5oj88bJheO033GKBw8k1OJPz50XEB9kWSjLs9cQus6Ogj3YQw8WLaRUSqbZiGNn0euNv1W
4mnxQVuYrN8fmyeYL2aej6Bjf8KMcLAiESZHKYSp2G/Qr+C9xlA8qrlT7WmKaRQB+x6dxEroqF8l
ItWdrLVKkUheMt46NpQv/l86r1Bswaqrso/oli6bbFokzBwweqPkDrlCVMHXWEBE/11bIyKsiPPg
5Cl92FQTz0EjfBaeD/NHPOOhXUoxhAnLlz+tFUWBGMBX6RDDlpxNpB0lpjcZLHizAsgKuxCeFcUl
KtrVldqWOyk32wFN38kzOjGcDALelT6PYjwHRymByrl9UBFLL8fSdqG95aHwtJQ2siAbkhhR4Mcp
tS9ei90jOxZdC2542lm0tVrRa5fQBLFJAlB4co5vWHPgWUaNB74m1jvfKacDR1+UHDFYNLdZUGTm
qAKgScD83v30g+BZAfa8+UHW32MFdtvwpuTrXfufYXs7EkBEnJNfO4Ytm2X5WUcgzCsb6ydLUiB0
jJuEWxAdFPaoKuD0TH/XA8q39+sseJQWbBh0D+i5YXl5aSUquQblwechbNrc9ND/TLp6EDguo78w
38XxeEHeYqRj18ys3g2jPt+ldu6yNGG1bd9LZMcCXDhyGMN+lFpCplcudNgHsgVXONN+pZHt3IU/
+kchPf1mV1Wh6mxL9zR4MSx2jhR6QIHbLrq6Fj4FkpJn0uKTDbUTbOU7RCun80oG6sppooa9eQFK
M5r7XVTB7ZJ3ExWi3g/Nvqnjju8MWT6IIGnzEfye/Uf/Ud0ewgUfaaGlqQ82Ia7d2KOq0sZ2T/8w
4pw8ss7i7Y4r3Vf5ogr159uX5QNU+NNcjER6rL5qPsES7tx5InRQnlnYTlpWYL6LhSt6iBPVQROo
nK5VvCbIWmmfyFBnp44meTygw7wYYjD6+Lhgv+Db/LG3pNzs1GPK/oFXkHib7bsgwc1jkqnv6rwu
Rv7FVElTrB/AiJw8d86sKmPnrjhCpTf7YR0zYsNcchvjOBFGoCkF04ONja59a8S/UeOMysaUlUKE
iMMK0bgL2ccdPdMK8w6kYi5FY3uDIEtZZqLzWGmARzLSV5zNKMo2Lrm+2bd+YO0/myGCSp/BE6LM
jhPBx2+N/57kD/qgpp14e6hRC3klcbrMdk5Gp3qz2j8WLQp10IMCPu9XvPG028QPdr3duM2jDuug
daZW1W0QPS2r267/M2ztZWXnPQYJOUXPYarsJAZYrG4DiIw8FNpMhjyjT8Na8t9QxMtVQZwRPSSA
TIdoTFyQ14eLEjtqP+ohK41qxfGJeA6DiBjLz8lT9/SS5tyneAjP+pMdXvF6IHAPXEjfXyhY+Yji
rqOX7zvqdXtCUg1glAxZvPR+7NIOyMdWBnWvEEX7a4a886zsnYyCJEgvXDfWIqPg8a9wiLNm02jo
mm8Sq5nOTCtRys0iygSHkgMHwYfqOSTTEU3toLBxNYLTpfRLr6AVM7OTUyGDf6vmh4f1iKCMQVno
qalYgKpdwXvYXWp/sntP6weUc1DrS+DcTKp7AS6Q4hi7EX8wJlDUZQumToQ64E1BJZpa0lDP6R6I
Wj6AWbc2J6kM/MSlKY73Jkn/QxpZ12X2k/U/F5hDNFDOTbAW59PKIyA2/bKj8Zfy6fTAiI+kxf9v
lUe1rn/TOcNm63sv05SQHJni0fNPfvdu6J4Qezzytek1ym0h6EtUn0lcKgCoA2/JcPioayLwvZXU
O2Sc0wYEbN8zYFOkcIZrBPhGUbpnOBT00v+mQpxglImeBvU5GdHPAP2xzSeMSgh12Ecu4I2ro6bu
02cCOeQj5qYYGeC1gsleeo0XWH8Y93eINMnYQ32JGs8PniJlTb43dG+umZHB9f1151Eu7P3Za4aD
BAOJDEHNJTxypVwGgz5gnfFNs2Z4AjGt9rGfw7COIoofecRxFAh/tpq7BkVvM15qM3iQ0p17UM+f
x6LD35WY1m+ZDSC+VGClIJvIIwSkltt+0i0O4BNpUsR8EPWR1wof1Wpp8Hy0mzHu7d3z6hTIRaOi
aygOOTSaDje9n8Ypcc+kZGTRhU0yLA5uWaii0MvLvfEeRlRjqpBPodljsM5h5buQ5DXLLxzxNvK0
rveNEdIR9sGE4N9k37F8FponiRLxYIID8oRbITsCadVUQXMBWerRj2mWk51rbcxnTr5SMg+P6Sen
1XrmXSQX4RlpxBvQkkjKnY/z2U/Z16HPxa3MXy0Es7gSQ5eI260G6Iuzt2je8262a1sjcIEmB7rw
Wyx3c/WyeZH2D4W35bU2hbfIl5tCK29kRTh9/ViOpSNbnk6ZgSbuNfhF/5kuUobSvMRU7yUsI1WU
/nzbrp9wms3Kc8ROwecq8yP3m49tfLiOBva5xMwox8QHg4otRuCQQrp8lAVsc2wAJpxRNub+4GGD
+7gX6ufZfKbE2yy0oJoF98+g4lrA0QA6KtGsfAG/Ws5pM1oRKxGEc4L0Aahft7ZRuJ+53j8/WsFI
uVaeW4whoZ5Ga0VmLlleCDt4c7t5+VwpEcAldFcJReBNhF710i2g/CQQtN298/sn5SNa6nbaudHy
RD9YNqMz/Xg0FW1QD2YILnzdSjtxhkFt2aX8b886+XN3oNJoDLULjJ0nsS8FXDJMOPQhmRiSLqyH
SzzIamPjX7yC6Prot10zNN6T2dkItFiwgKZcqdAfzFo0192zvcYEWn1gBJ4gd0yJyBWD8cs8k3k+
WNcPn7/zZTKhCydf9azJOWqNlVnXFh8aw3X6EckWK6u1fvy3ilcypwhZXPyaCDsYpQ2gGNkj0C6o
yjDEj5Euko3awuKDEarB4WWXLHW9DEYCy9QLhEo7qzaF0tY70IQllz8uRXP6cXrC0Bm7maik/hWi
5nnp25Z5fTna1qJR9VqAkkw8J5Y4ttRsYWfk9MmX6Ob2eSVjDareJobKWqZ2jHWrF7Kq288Bl40i
Em6HupSqKd5uKVWI5+PlYiVKBM7dSybADJzqTJzDoOpt6mlExR4BRYyZJwhHCuMyAWs0zycW0wlZ
FJ4gSVnzD9Ulnn7pQbcXz68xl+CcSgA8vkaxS0D9m/4VhYFQyxTNYYSyxJuYJ1ITrliOll+3SAAO
hueCxbWYBeAfabErBxwSIIB7h14yFKEqAodKcBM5wH0Da1ObKd7UOF8Gt+F81/nL3ZuEKa4EMZdq
wEYmixrSO/wNpefYbY7nmrSFicdvg51LJieeXRv4XpjWFWX6qaspdnzJkMO3hr7efKCqsq/bnlKX
pRZDLkwpGMH3qP/heomkrc6c4Q8HRXyUoVSf1/xmO/fCWD7BdP+tDmExlWzGCDr6RFEf4hnKmueV
01zc3GbaT8cH1AossRLioq13lnfdnpJw4/OMEC3zfVcG1CHRcWi57BLEQ7Z0bAgFNRh1ZgcOUd8l
dgiUU5ZUDKavDDrJAcV0hLViP/JOawnlAiCOjgeC6fos2uQR6mOl7dEedTefEC92DZAADBB/RRk2
jkyFrcra+VKAYQTyRhJCGuJoTaxKoF5ZFYl12LCTYjCK1BUJM4D/xGmDFnCWYEAowN3ACMRCiLLi
3TZHdliXegxCL8PwTddR3OTIanF6wvc7n0CLg3qmhqtmSQqzSgCTh6C8RmoHQgGwcvGR4pz1uWh6
zeJ2agSbSacx06il7GpTd6in7ucNaiBytoweYatxSGT6aEXfb/51Y/cfVedVF9QRLY1Snbzu23yx
mPkudPSPQ2eAUrMmlXs1VV1F7dS3KmtwKs64XfNcizd4aJbsA04b2IERzfCLTTwC7LTQodTW9owV
HKaVJGdVnFkCQULX/v4+IrObEShhiKR+bJS3TvsQ/QhhCf8cLY8HEdsU3BJ4u6b7ga2pu4FwtFWq
RiZ9x6eNG+VMKvWK/TuYITuU3Ohxu9jL/M4GQqcNrruaMmtgFxR8xMODEADBcF8IxItTlVy/UzMe
R+TEpQZA4irnvFffss4rlFtcDStsov9sEZIOk8CJefualc0tSKeEkA0O8eJq3Gi+9Rv3qXydERNH
7EePJ9H4QNeF9iOxHsd2xAE0tD3AE/0O7i8LKBkh/MaIESaiTANJcGd25LmE/fNkCvAjCEUS5sA8
q2MITqSmIB0e7HrJTQQYFi0wmeBnz74nQXN5PwKjNTQA64YcK4HuFD5VO/23JR9Y//psLrxYZ1NK
CUnTmVj8XVTWgmVx6nr8JgxBoZ5USjoQmU75YbesIi2CSd4g0xGHJbjiTZHCdn2Q4U9FBFVxC92u
WHyfwrT+rfdSFvpA4ZgW80IuLakq8vDV5NXREgmh+NsdF86cx5QzM7B1lqgEg3uYjfkd6/vvFVY4
ifB2G+vxm6vnSae1QN1wnRRr1aS5/8X/W5J6X91n6eRdXbpS+WCfz8/yYgePPKsMN+PHRD5kKIzC
U+1wrRlNeJ4LlB+7oKNJWr9BEcSDgH+zqIQTxZcW7N6n4tIDfV6LcxGKXsSGryHjKFaUszyT3DB+
vifiTdtlONF+yDBmiFSs7UOfoSewZvPfZjKGBmjCHWyVsSDkhKK18lsdWAr3pzJIWPJ1afn3oPn3
qctnco9mCrPhz44xeF27QkuQV9mMU4tPNSkbCKOGuu7kFU3MDafaYQ99xu+iw8BdumpmRtFyIIyl
PjY3C+5pVdKaPu4lRpnJyiI4mDhkt+I22Forz5QG9X0t6rrdF488W/GQNsxjSmA0y2wtc32qpyxy
TN/4VQ1GMTTPB25/U1aL/KZZrrEzjToisN0sd7W9iFMMpiLiGDcxhkDOP5WNMuIZVw3Mhj8GtQEt
6PJ0ajH6swDE9XomxAYMdWut1djeyrj67EompjTwumQtKAyGT9vzKajWkeGvMOTAQiXhFWDkfvkC
Y7FT/YPYX/m5wKWQgXGFmINXvIlt6GosgOpVADqTDqCIbH8vZoHmH9UyrEPHKCc/hGzPukiFQlBb
bPHYQ1BGwOgEmDPB8DX7S8+ZpXjEDCylmk0/VcZL06/2vFp3kgfgzlJ1K2VG6a1fkxrFFhLJfsOA
8wyWOs3fZUdiHZmA6npHd89ov20HVs4VXdzbIZUJdXCel6uD8zpB6T3nPli1j9ZnG/EwtDS7j7rc
zGtIWZJ5D08/uMCDl5qwCcRaKOkYkrUugTWEhAImFDUHJuiZ7ysbwM2UFM6KnmrKLmjluyBYBTMO
fLAfYjdgoWpXqbflvUmZcbg2MvVUFwm3weBUiC44yZ33Ll8HYFtH6foVkS4u7VT4YzizZQmPlapB
NB6Mr7stz0H+NBgev4Mfnx9T3+96sMh30615/W19kz0LB+w2Vq4AAdLX3SAvuhyo6a3cxxdUo1xk
aD0AbplfqiLIvVvReCMDHoI09fVEl7/8Tohfud5uqgaiERL6g0JZcjnJdXBYYo/uwq3+Rh+illiC
MeoYUSkPix87hPiaBjzu0YfKrVswdAicn9/MQrBTU6p2xW2d6oe4akAA3iLKZDbFDAIK5tJvjNna
k06wPR3NGrAdqOw72ERaOacWMt8VJEYor9LtJaqKTFmTm0F9wLtttDS+tGiubcqVFu4jfsOhpmBZ
tAiDIFA7m9P6qA3JvFEJXpgUveTlZXs2Zqj6ZTyiXghOeXZFiuaMry6jgm7BJXQeHEr5X/i6jn59
YQo/C4vshHMspmimIOqi8K2Y6MCLD0CxBG0Ze3AsrEq1zNQF+epempB7lm0Q3gfZy2aVw5n6+OpG
gpsAZlGCYvWyUoz+IS1rp8hlffI9Z/r9xMeyJMZN7XRy8W53v6psb2tjAkNr2Mdp6xDCmVGhcf94
Dm+ywOnWjyRRlU8/U8/iWTMJSJMLGa4HrxvkFWQSM8NJ/MjHRguojjxfVU9gkQjopFP8G1/O3qld
4QgsoJTh+jsjOVuz2b3N70pPdSEcOQbsy9kcQb+1EMxWmJYFlBgEODm/S2zz1t7mOOHZVpe3aAB4
Xo+OnaZdJGhNDZukIzCjINu5zt7f3ITzftB87yUGtMkZgBgfXFFcifxcZjUIpMwxUjivRzbRRlel
P5apy15jJymEQw+zKg2kYc4bmO9/+tfIJZ0aaHqKi/unJw+HMNo0AidUUfgW1X0j96kEBOX5tRAR
LMwICZF2sbGTw1Jq63q3M5arRol4d6EeMG87pbl/mG7UIkgMEivdUy8U+ohOBjZbtkPAi7ftMDva
rw7RxLLaewlGip5r4IrNssZVydBf9NM0iFknbqQcuSfQUXByBHRCfCm4cDjtzjICJjzIRgg0Wukc
c0c4OrFDCUVmpJ8UdTLwMXS4JdrOisMBAcAIpht1+FNh6EUnR22Z56Ace6Lv1klYyqntPyeae5ob
NCnErYvB4gmflZpZxwhDE/0Z9yafMFvwOmWxCjfqhi1UxFrDGGmglSrAf7k2G59N9odURc59o/j9
sVT2GBCBsTgOQ7dNNGWBM9HF/BCoche8TGIFtOYAbZbPdcKB681dz3bAdkKKpyQAgJ/IUAtLJOli
f1BWRMRWgwEPyvcbZyzPC51rL45XOmQoz9znuLIZ47ZYh9TSHTJkxJz2vXdQNb0CbaNd21ED6A2i
6aSpSocwnOSMN4aOcGMoswU2h99Gu9zq4t6HilFx/S6dlwNYb938qOz4uqf5M+qqRQfwR6MJ0qQ6
oUlTjFvxUdh0j2i61NyxPOS/CEacNhp62EFsy21aKKQhjbDRq0ervPMJOC7BiPuaBD21lO4hcg3O
zK1pKuKtnok1+RTPONZgCyvSQhYzt7vlv2prSfzpf/qp4xb4i0f5Mpm4bnFzmob7yZWTt+6E97pL
eYQTZ8J5bhGRThxg+GWy25Wwm+3xUmZb5ptjmBqCRSq+QEmPzyRLOE7UTBNtQYRWGm/DWDtUeSbR
l5eszBSs984tM2I7abQJQy+h92cd2fqXDdSA1W/J3AeGCiCUGow6yBBvC82PBg0OQA0QqEcPKBCA
yz7r8K44AQ0TYFeUGf9BLq3H6vXzquEAOOicmFugpuxtAXCoL7snuloTB1NfHhY9pYX6rXwzc+gg
+BIFLIDBFR91S6DxYuQyljI6UP+uCxxkdCKpmGTCNTyrY/q4IhPrfFeYXTYpukQU9TGwWnft7Oo+
feULjGpJnXHuzPldfansvsgzy2taX1PkW/A3nWQEGlljsj07ZmklVL3wg6NP5BL7FEK7BxOKRAak
z19xwE3P6sTSXSpjjY2wKjH7UJNydw5ehCAihPbiNvlxOBCQzeipm7VZUKEUkxVHHc+ATGxLMOHf
ONseXD70XVC4IkArucg0WdK2gUIj+3Npzk15T59cNC7QBsB4iR0lCnqllJcqoxD+6ysvt8gxvWrt
7lqVgBSqN7j/j9P8O7XIqPm9OrUH0V/Z+yPEXJL0oqMiVauuWWHBDGhmQictlFhGun/BFeFRrhIp
itnNtwjwi3puUHRDCZwssw7PfMxJemQffgzbxgAkjTH7dt+LI9tQq6vetZwOc2A770jtDl/Za715
6qffV3VW/DKz1gbt8hA3wMCLNPznc602PHkostshawgJPxnc7h1DnDb8SPgLupeVMNDUQA6JBat6
XHBUlL2RV42s/i6GNRwl4roeA3mj0Oor5BMm9i4EjQtTh3KrCu3vZmvQjdmQu1eqgWs1p9I9ypVl
IasRrIeyAUYaznJ7OIYmr2tBUXYK0/Hh4p/B1spwijUCr2Av5FkPo7NiG2h3+HNS76fEYeXFlRz9
5kJkbet4mZVTaBcLK7fr6VtunoZ6QmS+y8noB0erU22xK3eSnNJChdnkFMHSKSu/TGNYCe1RH5oS
Zoqk6dgc6YKMuysAz5Tnd9VX2/mFX1AoUyabmyXQB9U5aVdGm4SHLeccIxvHzl6cE0+reAjLedXr
PsmABcw/MmP9ewjk3Flqep7+NWVaDApi0FSPcbEN8FqGo/N51eEZ9ULXn3YRMVOr1nw6X9Zy6YCM
cJ5DVV/bKjVfiHYFHRqIjUuBE2tjwTsNUaO/GpSPjN7kNfdAf7gyCf49wP0Y8VFNy0dVFj/vhiRn
3P2VeKuyWmj6GdxPcR9y8OGsyRezeTgpw2ejtOy6m9KxDtdgaQTXukSx92VVauST4wRoAofFCp0R
Fo6UkW9ZYFchqC5GOk4EPgvNwk0Dtc6EvOlnvTdR2a7zynGHW99TIzv4tzo68LtK9v7h7njdr7Y0
3GMnVfYp1Ou1KbqEtZI5AB7OPbhqb4SNR0f9ZcrNc5/VsPxzlRGMuDV94JpSpLnJHnghZU3n9FjE
Mu4qoqn1DlLl3ogQCWm6CKYpDU9W/e8Imjh66tQeLRy+yEJ2Fc9k1QG+PR/oFV48xTwCV+gL8RQp
eMIr6cjsaq6uNpp3flYUTi5mdKqERUTYG+H6CYMWNDGqJj1/aovKaPoHnaMiNBkQHz3lCW7/daYF
htBLg3sh4cEvlPReYaISMLCe5HlARJE4VfaidNS/olPoShCeH2iXxLpDekU3V40v/KZsJWjwzbde
TEJjOaiXxA67xA9UyVRxfQqec9Z27StAFE4vUJXnhA1wbScJCBUiQqXIvNCAyx1Vf4VB+t2jzZga
OgfrR8y37njIG78YOa4N+5Nua9k6aoe8/SYu/xigL/VFPh1pFrUlOBzRJNLN1qW3jjAC1T+5EtHC
6gi+1sQgUfwRsnD2nI3jVFdTSCZc33cqKigxtrbAnbnhl5JTzUFp0IZnH0QKffH3nLbMSAlgbOFX
OymihqkOlDSZY1cAn5lzG0L8CZhxkhJCeTZpvg/vi+tAM8VHvOR4hXBQhqJ9inbDhrEJol2U3yBO
nqFhwhFrdl4NPSMtxwm84DlD+IGNRm3w2pVoEkiTJ0zFCSTrNoU9s/++Z7OXlQxwO8lIzhgAHXIp
+ytYefPzeeQRrxDCHkgSTN0Z7KyFqB1wsUSF7ZWa2U8esM4hkFb8p6UiPK06nXhDc+E1BUuRiWbI
zNmgTKhPUD+LE2s5ABMl7h0/oQLfHbpGd7r9BRqWFjUF5fnaEBUgn+rObj1GjopJB9ek4O/PaqEd
+rTlGtyhnuGWQDD0AHIR33JPTQmBC7BTe7gbemE2+C0JUhFwE3adJyJzatOvLzjYoM/IrKr/c1xE
l3MJaJCtLuqMvAx7a3SrXAHpGFaGPTz0E4Tb14nCv5NwlK++5CffxlOizxYTQDuedwUem6nMZvdi
Bp3WW1J4GtdCbRkonIXX10hu/S2eAK4CaNXRrZzSSJhtCwd9rUdb8MH7UEKl/rtFha7vMSGOgSxk
9NnsVD2+vTr2pJeCEZHa3nbrB/omGLq30vDw7eqy6pOfa9rTVd1e82mfmh9SNZV8QjyncoKxkq41
95s23PmAV6Pzg3IPeKhLMR6fVmo1u64vrLIOonFfYHLKhGK9MH8M0bjcAhdBzM7AnagP5i+3rKEl
UoLjhook3xYCoEjO13M8Wqh3UCqhfVlmrE+qkGPcL1OsGQV8LJC6Rn5zai7Jc+mWM4UWA+kplOPv
9ydH+aAvxT2Y5aRZ8jbOmzJHVE6KfVYfXDPcXcCqg6qdFX+XLSx4yxtRJEjiiiwUOKd8IxcRLi0j
Y0ApxSxmwlJ2zQlkkq987QXyuXvKxEUSXv16simE1PQi/2SM1tm7nRvI38Zjpn7lL9v7j9qrTs+a
YclAyBS7qVRm4b86hjsqTh0BM2BxhgpnMhRPMm7VfVb3yHQkQ38RXZr7OWxBFE7QMVNEMJdsNCAg
hVSsWgDm7ZVmNObBirFFhsxERzhqd7P7sSdvgxytMVDC3tGXm0IuaYTDECVgZO+7ibIqtShdpO7U
zUHLOMJNF1TtXcl46BSxHtwtkQ5uY7JsP4f6Fj0so2qOHA62YkmthMQgnwKxJrKm7ZuIXQtmezeH
HAxjSNQDaMCDfaTt6omg+VhDZPEH+rjqoUJ4CcEed3cSdI1rwBPn+2oyNqFP6pAjS7qFM0gi2yl7
bPKtOQpJLe0Q58ZyBxkoScryg1vPULnoXoDEyhN3cYphveMcvarD/xAdaSVrNEvJICMyfMuFqL9O
5r06LZCsEtEvkNUbrYFgTk7Jl25fsz4TtEA/yq1BYn+lBVAtzXM8tv/9WxoPWhmo9b2KPlVOGTZB
5dLwLzOnNCGl4KaZVyGxACjZ3UMbr+XxBYjbv0TUuoUU8GDZXyoLfwcXlpvdeUCj636iqW0Zrn9K
9Q3Ta37A53IsUWcVq4CiwZuNxAy3HSZGqjMEPzXudC3osSd3Sjupc53en7aH4/gyk0m+kIkrENHR
wG4yIy9gnKO8pGo3dfRVMAe9aXly5VGV3RlXV4p66J+uyCzayG51U27WFdgoJDNhJf9VzluyOE+w
83P5oA33F+Jv+fdQmBwK/FoPTB62GDNJJqnFOiHCCvEMu6c8I9G/jxOqcktEndP/v9OjjpoGQ+r7
BJFCGhX06rlRtTnxXzB2rZkm/wf6sUANPmHK4GEmIUB6LgXvA5Gl9s+e0Nz82L3GKHUnhV1uTkM5
x3ceavutB2W6TVcthWcf/ep6mBuiuyuLQPA15zFNrcl++2h3yMvZ8+NV/lqUaUghal0JUuKohV2c
KeUrAeM1UvhvWOnGs+5pFDpg2BmVt6BU9pCGoPX240QBNodg4VJ/3hGXWLpc5l2d4VCd34J2olW+
JTaavGEo17WboZbdlX+UWMHxcCO0V9B+Ztr8vhcs0+u6GK6czgHoe9Qyw7+8aR1hNHZCYJNUSrV6
rEYXBLY+UiPAB6iAUDaA5TFotW5q4Gw5Bcp51N7LPwuXicbs9psdLLBoiqwbV4jQ/K9UOJ4VOJqk
KRWe+obZM3cSul9vBHDOGSnT5sV1veHRgVPvoYs2MY6c4ZJWqCqXhlo+CdRNJmnABIYapHgP/xde
qcK6cdp2FU4kTGjJPjWTEIuub2vpw1rN+gJBMAu0oxxmjn763O/lqbQfK7lHubyaxZuHVeQjX13z
U1rfzfk8BCk9QlJlIfvKeI4YhAvAAY59iQif2Xyb8FU9/6sNQwxSdP1E7DzPbeKFzknEnQcl9AJu
D4y6prE5md5taYrYxJnAXg3Ob0ewAZ1X6oow39w0hgU92PM/Bv8JDDRFAVHKlt/Mqy4InFiRSXZp
8MzHkAonMgF4U32ZlT12uFSHzGfUwy21v0H03oBWt0ErVmwiTKjAZBljmSyAYXMIRH4MWCG3ps8W
pNXiQjDd3xPGFKAM6k6XExM2KheHFr1eAEcUN5XfIPNvBXQYL9zuV0kT86q7/xNSo7lbmk+wmBgp
8DbP63aKtjvd3khujM4QLNetw9qowqsO7maobNj9V2L5UIv6LWcdSQ03/stsbI3rWaGheeQhG9LP
dOp8hbZWJDLEVjkw46oQz3j+ZqorXEHoPAwrMR43Cvh9Wv3r/Alj6Osv5qim5QS4p1aKK24cy6Ck
r5NqrMlUzexoWIk3hhyy48erH54/ZTDI+A9a/ujXkxToKCYdMwfOd3Mkyx0QsZNhHOX2813XNOfh
B3uiAVMHCXZ0ZgqjBZYijDrqcFc4CW0vx++GM6CAz5t7rnut3Jff+5aXOf9mVIXv3SoDOEUKAJMy
vyb5D0jqI4PiLHfw84Rw26SgtEhHmmEA47k2IlYmFhBbmrU4At80WObYg7o208LYoFxbcY1rmq2r
jGtiatTdMMQuB2h16pjSAFYsWQ9wrfNexQaiOZNM8lflKph4ysIol1QB1GrNyYM4Tn1JypFZUS/u
SAJGAr5KKoG3ON94GuKQDAOKaiQOsyp/rsw9r16EIg7moEvTDvHkMO4k84PPnOG1Qx7AiA1fzu4m
6Miq/YmPmhNCTeYtMCE4gSxNZHisJ2BmnEjmd1Xs7Fl1JlmTLqV7FnKLjWd2NwLUkWv/KAGA6IwT
2gEewODlAepDyeS6C4Qu0xoJaPHKLzYus5RtjzDzGC2pTJY9D7QtW5PV8W0sjireD7DecJmR2SPg
ztS8mUEI4Rn5GkR9IAOlEVCj9pC4S6yStFsHo8NPk6p018IyYuE9uVaf0mlsM2pnLOwHblMbeYNL
AW07pO9cFpB406mW/6vxo5grCSmKgVkM2Hk2UBu3x4Q6+VoK7k7+VMECBa6qTkNss03rkRj93fQw
zTfOTLDekyi3HoG6Yyd6KNMbD7iXYG/hKcuFs5VzKpRMn+bqO3SR/OMlvOZC3QKXa/7kG3IoVxY7
dGsPr+kvruZ9onXuXHh7+9z1rUB4m7ZJvBN+8/1bjW6+MzFoVCJwTRu7EzRAQ5csAb2KKo1mbJFd
R6MLuYteidFbvFwGRjNKpoS+adLC3Qn+2V7QMqPcYwFyzsewWmmtNcdiBShZbw1LaqkCzku9gBIY
9f0ol7D1Ko9W2SATrmOZX6Br0KmVjUUj3yqiPB9KHDlo9/yr4G7UvvhmW9OF7L2l2XbhHwrGbM/8
sfwAzoO72kQ1FsBM7jGSd63WZkmIN3VM/7J+kq/IvSSoHORRgID/ErhYQa8/NlnjHrXTaxs1FGcY
1WO7b8c/5ulKGDDBnNZ4LTCyDcmfJpcsekuDjGGKkAP4M9e5tYW1nCt6Mt1arclPalqiKf7U06gm
J8uTHZQJ09VVNiNLxqOh/SsuoFI/6D+1QwP+188sR/ZDkzzB8NF3F1U4aU88tuCub1aSuSdjn2hQ
I1NWfh2RVebdOL75xsIaH3qvznHkdV4qbWq7ov82kDQ7kmjJUrxL+rHU/uNOsWQThVw9EEkXvbww
CeyfOSwlVGQPbjQVnIsBsSKNIcay2pTYE0+03UNtlj2aTu/QJNYyqN1FYzQwrX8XErgySG+Q9vij
5wjLaAEzEfphLTNI69xVRTaxC+xz/9zwmR3rOuJRcazPHy8aBM3hdlH6lyAKqGe1MNohGHlFvmDJ
51b4g1NHAZBbGwyH0xYIUVJxOvP82QmGAz3jIu1iFQkBiRAgwzSptUklYVDs2A9mzZc8znEgfhSF
EIH6RUZvO8dd79vg6rzNic0doI4EYrzVadL92+DSurPzF9nJkOG6iXQBx0JsdsUetVCQLRUHatPy
/pRVd3AFLi40n2bdzT7fzbc5E7BMl3dw0x9WKb3SZRBXhNDtvVDmPImafsw/U/6WOMclUnD23q+j
Tcr+L8dKgcK8eGDlgUmRVHSK/TcRpnBCuwcNbsWEdJnXrdbIj/vhRrlNQwZ3mFGx8ZpimYYs4fFm
0FNEvjqNbpx69/m5vdOq99Yxjc95DAR0oU0rKiVuN3d8QTyfxPt3GvoQep+FyJ3gCCD2Pkodyblg
qAEjFsXC/lTLakbabtxksF8n7Ql8oR3kJbhXm8sabcnGwkLFjNW2YegSGcl7NowhADL7BvmRbROQ
YNoFvJdRZG8hxwCAx1fAI2u+8/E/TzR3A+41xUgVMzN4vdBRVK+6bQk1w3LxjPZSZRl3Pi8+NYtU
7UovIB9Yt9vNZ2Hly7JDdylV4SQW8OEF9241Pic9RUL2BCy97TBC1kEIWuGZ/DFpxblEirR7gWBn
zg1Z/dsegPXd9YMr4xTUGcTyQkIuZqNxQYgu53nw7lr2GRsojiJNQTwAlhLg743k6W5HzjsxT2qZ
An6vZl6CfYFI/0Oeoh5MeHtirT8KZf4pB8DL+lG0S+UA7+jxE97tqMRFx9VrNur/+8IdjWjz9JBk
GURBXHxeaaLSSVAmySh6OW7tgP5b9B6f8MHwJc6RyTLJpRFFxYAKJ7evJrVnLgO2jEjAqqZRay5m
S/xHfjH5sAlI+xH1IHhmsQT4lrB+2wZC/eLvxflXj8kKuBU/5fl+kK+kZLVLWgrnhdtiW5xTNWj/
ZkO8paxrMcI1xLz5mYfJcawblD+9MUfC20tr7nJEveDVXavWrEkbkbleNTbGKcLz8cUY4I6LM3mK
M8TYWdQa4KaMWgNx+RMSZaedUrc6zrBlRhCeJ4QGpi6NbFD22ntOlHX0Kt0KW76pcpezOVc94q1e
F4m8kbYHDbhtnqnp+fWbWIc9LbA9SIixdkXBlS17xrKGdm2rvfLLV/adfIcId3UpdoqJWQmouqko
+Kqv6Lc/sd6E4CnlYoi/KupDHB42NqXDlzI31EwfyMN2Ml7JvCmDoRLc9eg97i5XIOp3a8Zo29/F
dB/e2dUj2JQtyPG4xB50kzyxPwGqet7Q9CrqZpCwWkdaXzayvNSH950voLMzAxCboIHUMPp01OF/
RRhEZ6fFlOUZGwPZBpMZPFVOY6WL5WsHtKTEFBz1zUPSYC7gJL0NYh27y/+dPLCbgWA8Ra4HmMVN
QeNdoavSVq7IXX4hyh5CGUuzfVWw5XTVD/7WS/J2i2rVpnbeZ+22Lts1QOviJysnO6KSOirFaHZj
wy8gwx00E2ngQhvY/6L3hzspCJwQAQnbF+xSjtmp4y4yEmlU1RyRbqGDNL7++EYRERt6CnTyP+Yl
Oet2DlWDgVV8zS6yVX91s+DV3pdkghrwQ6dyamhcmAemd438d0EmRORW+DbsckMHpH/aquFGzMOu
pzJxttK4x+LhpE6d/HzJAfqsRxpDA8f5nTgxFHOKcv4nioK2cxVDAzolrJ9W7gkb6EjI/VPyCx0v
4wuMSYIl4hvCWhEYHIUOMt9nq3b4H5yckIDWXqENEVjxLgRYl07LJU71Fh7wdVnfbCmyxgizEADt
5T1mt85yX7GNgZmvvyBwmi3jM/fKOyuOb77VnL+FR+TNkO6Ok80fMfIEmA1IkBSWhjQPFedbK/o2
jwzqh32LlS2WoWLgKreI3P6HBYY923AUdBR/1xh4EDjTJt8E30oUjO/FpKCIM5MwEKqgkFESiC1z
2ZdmB8j7uCDd2Al/Hwz6okE132pGNtYamERqb5amoq9f4aacZN/Akd+1CeKJut8gv235IoXGmHix
G+vnmnIndpGIEbyii8DSae6ZsM0eKFwX52ahYD3Dte8sHEwodO0PBSV/p8x31p4HNx8JCuAZPV3e
otDDagfEj4GI8hKlKGQZnhSl8FMkg91XQ41OAqEa2z8j51zTm1mqqcgkUPIN/Yiks2EZE6vP4IxN
+A+CqXgMVKLQpOXbomSLzqoLEQzhExQiqjsnchnksZrZVKj80ArWOAVD/S525CGlvoTfDVg96fzj
unkwNucc3kyMaU1swAMBaeWOmwKg/s63dxtNfVfmZcpA0sHQHcW4UtJriZBDqNWxIb+qXgxEnc5L
yQuYrYO2UbkZTd2ef3T2NAjRPPpWotTzBUx6FiJboo3a40Rz39KnoiOU2x4N8YnHGGFM+tyUFnRm
ZTv6yFXpDel+LB5OeDbBgrDfjgZGoMiuL+WXoELITE02FZ7dQUFTH0/Cv3e2wcM1vhfXnxqET9TP
hv3MaPlB2yuzB53cRH4dzga4M387HBGXTLd3P8ZF0fDC2ADZ+xVGzhvHHtmvDUoYAIiAsQzWJOxN
0MFa8gromIzpkMrBK8SShmdw9oltOLyV8uGvSJO38k7yYeZyfqCpjnMFBStjzpL84nNPxL+QdJtI
J4o2fJ//2uS8aY4XO47+50qHVAyQi7Y583YL+8H7CfoDZcBC+HfwwWgZoMOkNsBohx2zuhqdc0+m
u7WvTUGFMApuDQnG5YJK09EWty2q11+sRqpXsA/sNbhhwUkbtotFF0CICCrM+cTmic8GBYVLMk10
udg6p3tAgZ34haya3mURiRG6+pbUaDFPmbBCrMD5ZWejUWgr9BmmzscnVvzc3o1/0kiLYRBRcV1e
xlh5c9kIz4xAUf6ezoMiyW3hR3JsxgCiyZfmPY0zm6Sgy2hgeuQ66IpjjyHkWhoEAeWpLM4aoCLG
sIRbbiSjUgEvnsNerYAW7z91LMFUDLuOXpg/nGrxS+0X6UgFBLovDCCL6Wg+V3t5W4yj/GvFGXvt
EW7mur+edK2zIE02KRIxOdnR6b2b9uWNwrdifhxBk7RxXSUBSegk26KmZtxC1X7uzwHv2DYV3Ghd
AyCdwIxYmQeeVa8CQ3JXYzNog7ZJH5Dd0UKb14WPq+G7UgihL/6A9xk3Jy2NheUf3sHb8ltVc594
rrd2TWq2u5dVk3AOnbA94z8I4UmKug1k0AoSdIEoYeNWC6dKXx/qL1dB3tKaGDXAJVA/iK7oAhUH
Ic1foySpzkwrwCiopdRAwIgFePPWtOTJA/D8VPnGV/ULoyKkbeqN/IEUfEfhb6vl6p3kOXHm8wCb
Vz0+NlU27+uPCpBkK3R0sbhDDMrtBgNj3S6bQ4y8yonIdw63krExu8cHFxd7Fg2oQxStlkQKt5x3
jyv9Nv1mK3RT6r69Z8EheImFU7FUd2+AKHk4ArGRfbLiyZufTENJ/Roubq2GJr5M4lvTamAwqbAS
jEoKQj194SASdGRcPepslvoM+RfRHhyFPp9eKihpbx26XuBeHTQaLwHXgTqgTMt3Fz+BI27XIMIm
lkDZTR95jHo1YLK8qq+/46ZWLoXjRuQV6eadmGeV+cV404h/WfTOefqhqlKgGARIGxvaYyjux7hT
KWKalqItVmIwxNAe6NPgPV6JPDIzEWuAHz4O/3tuaZl+/LUx1AWazRoZdg08dDocsBOWQuv2LvSL
lCv6s0zZPXoE1FKInwEJhou0TGkWLecFga7mX4igbDKhghe5U9znbOJkDUXyfqvfx8AD6pIQk8XG
uBQlH+axuy1zTBlrLAUyExiVMB0KqVwBLvbz6Hic4K2hzffzGiAbo03TaTBOWadjti6OdEYcYQmO
0jrINz3LmRMcr4JVvlUv0+H4D+KVb5QWGqfclhfkAUBZ5zL3Uws4k3s0wMwmAoBERZBl12w/eP81
1CWL1f33pxcnt6ovo6WEmi7ScUACFixt1/YPEy2jnOkfkYNZMWPR8cw4+CVKMHVy0RonJFOlpeLG
hAVkb8rjQzdKAPhyPDFhYAt0Hqe4w+RX2AWGH0OhVyNPILKrv56jDwPYpHiNzSs8EVbjpUi/5d8F
iZtpfYq+XHn9Lh8A7ULJmD0ePES2Sd6qp+jNZy+R8L+shX8T+vQJbykNDorvr4xIf3pegk8pnE47
XK/1l5UM79xV62gXf4WJRb/Xuxv2550gBj9D/roHaPkGXLQTSNJ/bdqhyCv7vaWV+j+N8CllCvm1
CtAVBBGge6prfWjSbMa0XgIlHtwygvlBPePr6LHJU+Ccl6fnGO1W+wExfGBoCm+3Dn4x53WdZgaE
ltQYeebmSt77auCqW4O1gp6sng95o7CF4WqMpXYj2eBcFoKEe3iva+KcktuQ9sIt1IZDQGjmfqro
/5aI8k/eRM4+9FOspu4Lt+JIeR4kvFhJ9zjBChth/Q3mjvuAMe9ToExGTtPFUjWCWwBKpiiFIG/8
IASO8Da2t0gozxswINFdeCtvm9gvw7c9uPU4W+CqPuf5heDZIt59Oz9dY+b5ZM/rbg4hV3OsgbQe
zcdDlQvzG82bHnmNgS91xt1B/l1ooa/0PiiM3t2RekjyG2c2KZJ43Ji6EWXXNHH4X62F6pnmYl26
aFjO/NqWlJFBTiZhgCoCx4KhH6xWZeOzj43MnZB3k05Bd4rNgyOasbXJTTVhOHbK1fW4Cfhu63ze
/d1/KZx/zZbF/6x/177QLVfIWGa7iX+gIX5os8h9Q9BfQUDXQHykikiR+rnjCAyEy1kZNnI9unre
RMFwCpyyioVddrXiGhHX8UvELmSXYSOHymozBhAhlTxccgvzHYx+AbQ1d/6DOftvVNKGVlZdE9dX
WLnc4cyH4biucu5MpCALrpZdGo0PEMwWI/VKFI4FyG044LK3OJnWj3OLDdQ6Q2PpMIFTV5aUkKo2
qqWdpIqOdL6U5OLU0kLmfaOK5Q9SokS5sePumaPfbew45wXHWpFM1R21hCkHRlhhueP/aJ1qBCWG
92Kb1N30uZEOXN/NFL9NJPm/GE+IdZOdrOtLLhCOy/kilL8ZvL4TXUGnGSiz0ESREeIrSSDLtNCV
UJTBQpVZCjCoPmHw0gtXoc8Oer+wG6sSyac3ARnZXbMe9PX+A4sgEV94MXWfrOfBxlg0011VpgON
IdqU0KCToMTlwcfmP2jc1dyLGdF1v8SVMAJYwDtWZKPqOo1RiZT/qStNK5zdwtwDk20bQn3KplZg
UGzqWJdLzGkEq0wwivoUcgv7L2DzaBgdtMBCUfft8UmEqda0LTxWWn2ABTZdz9rTA9mCDGv2KHVM
g9/3Q7fg5eR3ueiAUZo97oREF89eY7ld+NNIAzQe5n3hWk8AtpaNsG7KZWacwkwap9foHdo/bUUQ
MSE6T9XlrOXKDsvUpGGsnv5IGQwDltUhvKbPKPpnbmhZu1Bc3S1W6o4ZpnL47bK4m6akcyswiVVt
WOpOuqPUuwiz2h2NisGeTBGtco8fb1mX81V+dc2Fa9Gksa/abMxkYPo4CWQDobeY/cWVnuzPKlm5
8UQ0ZyN64cNfuvDWGGgb+0Xr0QEJwpf27H3JF7p9RszD7C2Di1rIi903w/+aboUD53VMXebXeu49
GtfCqidK9iSV2PW8kWoJkZknXlXTmIdKvtd94TRJQXD2sMTJFCNRe3I5p03QG9pQCjsGUsH2QATR
5Cpqy+LQmjG1q7WRLbgxMEYfNKnUGJ2rI9ziuhfsE7xTyfTRYufjsX+OGkFDF9LwFD9zEokXk725
vnDe6HRc+7+5QiIez07TaxGgZbY1hw+rC7US6PrX/w9K3cjnW8kGFITr4DNuLyf9kni6Jwg5wvbr
Yt0lt/9XrZcLMg7DQ68ttJQFXsVKbE6KBvDfnylCqWCLCvQlZLnDwrIEm/MZEH58/WKTCBUTYgaC
buhAnSLTAbREBow0HeHjSy2627oCtyRLPxPCpFI/on2NJHbTG/WnQudQLPCGkfiASkAuCoFsbW8x
+TKoyBZEwueoo5Vadk1cMHZjZWI5R3GBB7rL4MOS9WjdwRpeFp7z1z3ycKoX4jaeAa1MeXR/uHGL
x0pwrrImLu9xw7fxqlJs/HQpb75vielbfudEbLfM1kUHAQbAquC7v8p61F8NtF9HrgXJywRDoo7f
lFHwoDNQcbVm04gWmpNERB2VD6SSi9wCbEJ4AVXRHGSA2v7hRgC02gLuCSb/RTWJ6GiE1uYEAamE
U6LOLEUTzQKcAiTecgdECaoWpmzrssDUgrX0yJSs0omUtP0y4WsEfEAn9YOIfHj55ZDx3uog09jj
EcXTsuUDVJBRmkkSUu5JCBdaIz0EdPHVQ4XzPU2J65QU4LOUVQEvJYsInQuQloHWjkQgf7SH6B0l
DAgfxGHaTHnLZpqmBfa2hWq/IB60i55YTPTIX41xMaBkj6UJ4JEyoH1T+LODNp5BQVw/vi+AmWl8
T9L4J0INVzUIBcHe4hWs/RzaOOpH3OP8Tt5f1kYNpTdnFD637yynbOEmoVnz9RoGzCKDNxnsOPnp
RBJz8bPuF0KmDqNTeuEamhSLNls7wXQ5DCtzkCxHSBZFeXauyMHxjvsa9kloYVNAJBYVjnX3YXkd
lyDItZxsaPfAn2/JywuGOMxLtt/hKYQrH2Uo3xCrKRf0Lok+sOoTqJ4sJTSKK0BbilRSo1kOPy/r
bB/xPNqqRfzijWnKst9WIPRh55MZyj3mqVtCyxyJfe9941gf9x467zyq4r0l9YgJrdQF+SkeNXip
i1Ho/AXYN4zCsKBUIyE78BLJYEA50tz1M4K7pQLV6Z1/qaqkfKeuGlwkTSXhLIA3YRoF2gedGfyb
d8OMhTxjGvpKR6hSVozhdVNs0OWJAZuyxHKZ+w1A7tQAIF4M2zB6BVHH2LqnNMLzwTXleXFjyP1T
wgV6KTV3+lIdoq8pnvS+9nR1MkV5Q2NUL6U2oVbHjCc2pn3WO0+xxuVcnnTSn+p2LnN7uKP8nEg4
vCsaDIv22LSKaGkA54R1famDNprowzjwxki6uK/fpR0Yt/ioQJqCDuitYKo6wtrtR0AmGr+I69Bf
ZBJltdSmR07s539v+d4TuLie3/xyL6s93wS02uRL1XQxxWhRrdT3WWJI+RrYabAHnlbR2qu4is1D
iyLusghwFY8QJDqgLjDG6yX7kIEa4dS1jHnQM78zNzgpW0huA5rgIk6ciAhrmZDDVRu5jGkoUnB6
QdlJEzEmJgynssw3urvcs1W8kuGVC+FZXz2CoKF965xJ9C/FjOLffWsIjyeixphyNGbDoKjr+zkZ
k1N7UBraEqXNHTKbQF/S4ugLxTraLjgmrz9yfFuF3LCK+NT1MS/H23R80ymhshn4EHdRC4PSe+Ee
mtLb0dTkwMNe9ceLo0N2OM+vaPsN00G5p808H5hk3bmMTHV77AUWCEOUxHWqV6ETiJozcWlcjNII
1p9MK8nZJW+8zzqS1kPtwtEvJC+BM22ZxUglfjqy6H6bGickDML6LCgZpcMw09x8EVmWdT0yCrtE
cV6LKfoHxydc2pPq1oWUrvqzLB+HFSt66aVcksfxsJ4a3cg88Hh29jUOVHZMLetyX8mnbX0e9o0/
QoAgpUqtHyy7ceJ0R29EUqZQ8hawi2dsr0P9o0JBsHNxFRYPWbUMyjVF+IGcNninlNDPf0dUeLvH
Dt3RhvFvVehKTh82nKqjHLqjf7qCX/ViD7Pj0ijEJcxCm9mJN7rMrQsNaClv/yv+8F5U6e3QxykV
0SHGr+7Pus1n0scPIKeu8xvLQiartdpCQnCH9wfaXDv4FT93xaLBcMMGDxkVoDi4CiZSK0sneFn7
RwekEJ7c+2Ij/uxC4Yc2tuyJYktHD+yezOprx6WrYaFuLxeNLmQVMg4o1kWnsPNM4XJbwGO+1pO1
RghOYI5KGCyCX1v6zwtDqtkF2AIDq+/OFhXKZtRCyO7YM09hrfHIcLhJY6E5Yp4wfCF2RwRtn24p
xasrfx9dA960zdVGH3vT3J/iYcg+/+jbV/YVUZ3zwSSx1HA6sr6StNn78pY7LkfKQw+pwuUJoL0I
xEt5tvF0XjwAWT18tCUsm4hEXJ6bCtvdFsKbuTBpj+hgpcH7AL3NaMIQ7ruaTCIOXzK0cIi3NW+/
4L008c7QAZBEZQgMUUjk52zcmLI3aLQaekqNu1MBPqJY7gSimwHX02SC+SLh/Okt5G9z3xT6KwCP
/jh23sUsADsh5n3ajanOZS6PSjVvNnDs/TGKIP3wBcCnzI2OZHQ7ZRq0vSz592IFGjov/12MPjN5
tiVYCdmigdvo6+SlcKsSV3Nf0cLplsAIFhQMtbN6CSuUhhFFw2Rz2mIX99diUo0GTW6tZbgCruUO
s6wBdOYMt+POAAkA29BnnGsxZOcZM+adOltL0LVsTN5O1de83lFeFscts5GtlZAAKJ2vBpQ6oDWV
R2NUFAFyUVTc8lz9PefXiI2giOOdY+Mpt5I5Fyx2z6jJ6YAnpff+Fi63E91acl5sBMC0CrTK86b9
rzlSmKDRrZw48DYjIDcgJ2rqoFzMdwnEgb6XGePSd56vc42qpwxpLl7rxrGrm506CUz4CPgR/2ZN
woeTuTHtDSeqXdmOK8g6lV36aIE79BbOAzlzLW3/Yuc6NVTVRMOWZw38insld8mA/O0ibDlbzfHu
AsOsJUs6srMy9nRccQV1VC+b3XBDnT/bpBJmMMuF7c4lAX/UngVX7frFB7Cgi5/U0Y8eATkGvcRH
ldy/syChr76mG1XpqeenfdX8YRdm7rzG7uhbBDy80r18uhs8oVwthqjO3fY++qPsfCXh+/UUcaGh
0iUk+0Q/dmeucpcfok8NdpAjNKuol8ic+vMk6JgBLqFmyRyVXjsiAs96h0PcgKcgW5/KMob8JQ1B
sn7+8mMZL5s2RlJKCjqFKXEXa0o5lYDLd9bIikW15HJtP41SsiejgnnhGpe08JeIYuD40Lbq7Mfv
eeKMJHbyi3XGawMvfflTIkoUMiZAY2CQW9qlvWbhkAHP4ow/bo3M1pijGBWtGTvVjXW9p+IEVuBC
6OHsCiMxBH5b1sODbJZ1z55MbV6sX8Nn3Uo7smAMZTCCN9WQhPijyj+aR4zpUQiggl/Pgwk73ezF
hNkMPXEBK316R2r1S8+wM6x6zxRDZiNRHltuHD73grmS3RISmqLNiupSaG2pJSQgZ6FHQVBjLio3
P64d2gfHf1EBBAw9kn1sJpisY6ZAX4csmAFAwItzVbzcdmDwmmlnaiTJc6WYkXQ/6mMHpjlZ71io
Z+c5gsOLsY9Me8RMGPl4dz5INLNIXFUO/AInY/EhJF6x/uh6bE0BhoJvaXqnm3hzZo2V+dXVW4GT
b0bjED1zHHv4XuO0ta3Z6ckZ6IuhabqlaqKdbAzcWqCT2XVmQGP1xVHqJx+XBAYVOzEwDFqmgV2L
LexAFBfHyhUHYEbhKFoy2AFB07yIwO4W1arKiMCkkzpPtrNzirx+D4wPGQwBsUJJxXMJ6s6OqeqQ
KBkfOM+8h2q4Z6GrblKKeXdeVdrfQ4yX+4K33hLrg8loTO4jKhg8Hm9NVVJFX55RLk8Fd6AmLbpU
yNaXTKlNHAJ7d8RsHxzhhnaXbzPAFhXmSbJ4XuD6hxximTUbhbdUGE7cL8uyQaRowtwDMKmRucj7
iXEdhCzHs2vGE0L40pjdZPDs8hJheYTMQSgzalXDIKz+8DKI2gX2DROC3t8NNAYYO0O2GbbNEThz
op54IuLI/okRE+MzvPl8my7DEZnz7iSZ1x0lBl81pRcR8nH81e+t/VAOIGip2VL87D2JVzrD6g+0
u4gFXns3SycMZvYpEf2oTjnPnp8EJlv62yBCH04rX2go2/MUPbC5JdGIGh+01NnqDAj9zPQOEvFu
SmMwXH5NBjmMGaAPjGwkPx4B2ugm+Uf2QN8rWbynt90Y3f5LfzgcfsZTWlLuLfjsk/OsLp7ap5Hr
bYL5fmoOx+EMUP0KVxM9oiYlvkjT9rI0w/2ZOU3m3K0KH3BuoRRbhRCD1RKsMd0hWVDNzw5ranp1
MfCOd2sXbBdb5Lz7Yc0wuDKnPR53hoEVBSYwwd9/R8H1S81j4RZGYJTG3x6fRsNhisFul8R5q2/A
AZNIwEmtRcWaMQx1nDV8CzhyX8KFW6t4xccLHTXyYgbqPhLFMGPtpnjonfJD+edNll95zOHkqo88
6JduYOt+344NBRE1qV7kwC0RW+/J935NDK4T4dHi0nwBjUbf69N5/FX1+pL51W2Vlc6naJeg6hPl
weZzkGoby02zs/g6aIQBgrXc5G6u+Fif2FMbo7/7vVI4SImVrpXEMcg1cHfNvjBNXFkd0SbVSWXG
0goeU+FxGX/uFzRv4O3NKhOZgFtyEZX6yAGtpgamtBcEW3qO+ohdM2KpBhFP3w0rW+a9/kCTgVh3
x7Gca75mj2jgFmhTaZc8m2ZnOsadg9EUx+p22B9k8VgFUs/QWrtA6JY/4rDsuD0OtEcHnkDlPrVy
BijvJwIF7XRCZ6hJrm/IWdiWgKWkrHde3Tm2IUP1iwzSd9ZyjBkJlBl92r1baDNZTksFaGW++y6S
b0fVBeH4furrADmYURitPJaxiwUIp+VkK2v0x6RZ4hPuzvlQZcLDRceQk/iiAQQL9Ks4MuP7Hi7M
aeAYmPhc/IVbn8cfEBA+JzeJU0RmYLczorcSXbNbcp6WGwSx3NVw9i5+yrhN1cfx6maQDieTmEKR
bA9sr2KqKrjPHB8vtGeVAwlvRct9cnYBh3fJ1CaT57aQoT1fsUzyBMYuILhaMvHXQZhr//HEab3c
cxxeccjIXK4QRc3PiOThO3k3uThyv++x0pabRWkCh3F24FwFuiVPsXnhxXblGXvbh2Ak0urIC4UX
fOUe1drFYjqk2ADCdfQ6SIx1NQq625zqn9DTWllU+FZwQ/UbTQV3l3jNXZzgRfDdmUePNdQ2c7WX
4y8uK2GDgRnwdhBBrOza+YOCW0+VvLOcYKmx5qCRISod1dlKtizcsZ8LzgdNwTZu779aR75I3R2F
VnNdY4kAsY+l48F1u4xlPUv7+1CJS/JXM3XTUvi2QM8rQTog8QtrxCaI8FJEnjd8CFNTjhFxTDfh
HHoFio7p38KbSmzafh/WaONx5/Xk0mga/nwq0Q3lp7ky+FPfJUv+gbCKB0HIbDiBACvjiieeTYkj
EeJglhHIpcJIb6CBaBDVXEIuDfdCdR2qHlatq8eHH9IsVp0xw9lKcbDJYlUEgKINSu7uolgNN2Zz
MHZv2Yrk3D5pepP576XJs8UU4kaAeCsWhClLMR8U/xeAnNTOBzJ27LRBAwtOV9HC2+ddnmYamccq
q5lb/mFrHiipofOkGDcRFMSmxzWZiCqHbweTZsKrNUT6B1b7s2ioP3fUR8j4WiWR0ABVHRfbBIcC
svyJgvFLSr0s+WQyjBODaAVqMZjSd76izMcBaeQQJJL7vrwWmZI6PNbQaUBXRhsyCBpi0ScBhbgZ
S7mL+8Vy1QTB22nkjcwkeGABRptQPMCSEHi5P8lnuCRF4ZXZ6luRz7NcAs/KjUqPiz6CXL4yTJQr
kyB4KtLqP8mpX1/BCS17k/08SKXWTyZ+suT//vBUTDmuZnBcWDXUOyPZJIcC4lxryM/s6lf0QbiD
z8S0PCu2e88PhH0zc+6S8HezqDBhL7J+ehKQK0VE/SoPxloyiE0YQMcr12KUHq3Y60pgfHYrLdm1
9GURzKcHQkzhkrkF86AP70t5Wx30tNxng6peOFJW9ZpaDHWJVI4JifNQQ4jiIdTz5a07TXLSFcU3
VYTGD0utIaD/xZw0aDUxR+1j4MiIHkumYx2i9q4FsbtR0PAqCNSnS/s5RutSmWCPV5SWu08bsBBC
4twX3KaK9alkI2HpWWJn7BOuK7dja7KpqJcdVWOrkJ8roUNBOj6Z9tnDIfIxVwMtv87oB0x/etrX
X1W1ItcLgW5YjzF22L0rQ/ce9+vGj5NMQlzkYI/KLsO1rUmi5+bDjxj9mvO+ki5tux1A6I7lGvNt
InYyS25K1HD95t4ZiW54BRhcRZSZkKsV1SaZd/xLW7B3t1jikXGYQ7A7ru3Ewl/nzokPXrWptiiO
v2jMHWf09x0yYK8/WIQ4LmZ0r209S+mUu5wFfd3LYvemubXj5gdPAi71S/zpIzwrKPWLlDswYSu2
BICzJhoBxK9xiMljqzFLmjUUZFhYtDXMuk494FpBnaSiULNHlytEiM5s/zWBAsd2LS0K2xssAQWM
stijmYXwiEZxvf88e3cHbpmLSWkW3ALSYy55WUTF0IDy6DqJhOPRt8O5qqbOC3iUFPyQUcU852Ii
0Eb2VhzFMh138e2YQtMoDCLWkSXssQE6rIwiYVvz8E+YmQOHpPKzlxvlSstbAsCryJ7yGl29dJD0
7VdO7cxDUEyyFRJPhCOY/yij7aad4+FC6GwjReyzvQIY51b5aLumbWCD8u7bN9Tdj3O5IamCZMtb
aGU1zmP4lneXOgPt/nf46vjTUMF5egctNyLBdWtvaNErAo+N8PHY6VnV7D2jyPVp7nDJAfJaYG1L
EEhw3xlZ6hY1YP9DrqOOvdduvEGUtCayCzLHGpRoUHvk2EtliAup60Pk1vC6Gi3FpAdYeU/006hb
d7e1//+JqdyTuu4V+GUzd32rgrHyzaAy8AhDSkj+37TTD0eLeTshEwaEfIKpZ/l8qmOq1i51jkWV
Go9QJjRo7C7xdmtIfO9Wi9oW9vlt/0bJdjOKGHbYwExG+BhB1Ww5i1/KAfxz6UzZnWsRfCtc0LtR
MmA8cbS7niwKql3uzdGEtPyKsbfbKkgKGq9+vZzcHANGSpDSBwfkn0hSjfszzzySdtii/2PebkhH
BoK8AI1IOByMkjLTlCQt9rMxYZNsYUR7pREu0FHaPNeGqTLhIhU/IcP6ZTR2RRWncujuDAJg2e8u
u1Qyhzm8050vzfUjOkjEkxtat8zZeWcC/jQStAwF0Qy6L2nep6aX6Glrdk24K9ovNdEAWdLN1tpE
NbE0NbD7E9B25SfD3X7m5/czGLU5iFzS+TGXhfRW15f0me7SZ4PoNjxeiz/kS2QesshHWLcs/oFw
DtdN37g6naVIR4Adb7aN0fPKjB9rSs2s+QcqzEsFVQWYoBN9qEhCcG1gFNVHhiHkznLY/pU8CVrI
tDA4fd85yZ9TAq3i1im5QVFJL+xZT/GR09pmA2BcH/VXQkBWAgxYRzpnj3iF1ZIeOF1XqBJiAVqy
Vwje8dQ5MpRZ5+1mDdBztHMtNuOp0x6yjIhuCSNNsVUae7SoDQCw4rRUDpyqezN0mo2RxF8m1CYA
BfnCvCSZhJYtCOTvHgpLtWsTA2eVhL6aLBmJw6OPdoNRcEcIy1RAbjXDXV81n07FvGhWgy7vLwZl
q56mcND3jQUxP9JZyE84L+xJURTkN/3Z5A9A/KDtnaefJz36iF3JdcnIs6U8dssmGeZXew+UrUDF
q/TeSRm3OCZAZZcEwveYYNVIUJdPV8II0N5EIopYHVEenpUXKU4Kb8AuQVVIzWOfvNnJch/FGPJw
FO3bG9IX9FhG3hDGoR9N7bi4L1veqNvQ6ZyeSYUKL+KnydLYSSa6mba/IWqm1q6ZRa4UC6dDfSLj
IQEe7I9x8k1YGbbRRm+aXHrZQrGZX9DmunKFwxpO8yyIWP2qv1K/lB+sS2Bwi1U06J/C/T+reWix
bstBM1NvXjPO/Pt+3L6VLoQgJn8BxWkurnlW61D2trGYjv3H8+4NyjxknDH+PnuLi6+Hj6L6Sbfe
+lcmLjzM6hw5PyYxIsAa1sqgMkJZ1wsqTvhNmcB7ImgusTzw00QQkjqd7FekFrwoq7TsSub0syJw
MLKJduXoa74SxsBqsRnPpvUuamohHYykXvzU4XYE8dcEeVVWxDQcENl2evkjLeeH4J99q1xJVj4u
Y1TUTRTiBeAfwIsNAVJF290g1Dp5Nm/ADC2cYFpDdjfFnarZhfbrR8lmGdtUqINOUpmyLAMBEsCV
25aYK2t1NsM9In0gBNgDazTmAB1CAQWK++NIbNYAtrJWmnyQcv5mQrxath0aiM9DErQnzh47SPWq
fN450A8kYwtUL0+j/TyoIZk0GwLxHcsUuYrN4a+tfT1kXvgJDg6eQQW1Cg3hnL2hnIWYzB3smyG3
v5bmmJpQPg7nNVxej6w6hTA+tdig0B7OPuKQZSA5IZn5Qsd4WsmavmIxMIaW3MRUGLhNY+j+6eI/
5jFRyqhQV/2c6QH2chP3Cszqu7VtwbhqZXvE3/WMnSAOk3dB3LYdDpG7/iTfDoQVpSfBaLMqtwqe
G4qM2rgkbDgKTLj5AU4b+ojmkj75X+LWSyIfE7bo2tWwQyLXDyzv7dSevMXDIHS9w8Ith5Zzlt4w
iaZnKtnf8w/dqPrRTLUW4/IMLL+LJCkYvPZzsmuBIqH8cK7M0cK23X06gtuOGgdUTsv0EKi2fS29
iCopP+LHHnxBpAaDZRHz3RGibFZwVRNeHon7wISPPAPA6Ha4EhYDQ1C3rHFFy/4Z5uw5weXA0A6c
7ZDIkAsZ/Mt12uTgOIZ41OHdQgJOE169lddy1vsZJYbtqKEFK+MRzinW5XWlZsyVzgHE8rH6SKQq
elGBSNaICcNow5OmJCqH1QTwQlzqEdzUCuh9LIjVt1RLLLoOXfg43thyjZmc1xXSuNoDwZzShgza
j0o1SsV/xZD8W5mqWRKVewPTGsZr4C3lUbXjM1WIHE+Vr+9ALFaiju7n53Nx5saOX6fO/VqpaWNa
K0ZM0ZjnBxcKUHV85q8ni0QP2/LYC4tuTZ6vScy2RBIUAyg4l9cbPaPH+0u7Mmt8OqnXaimaEUx3
+4EQqUu0gWwVMrsVJqB9rM0OO2kvKhxtQmg1UAsPyCIGWcfjoN7n+COAiZwkht8RdF1WKGszxfgo
TrnugTsFdJcwtfagcZGjLD2KFtlKcHyi2wsQwdGLCI+uvg1/eg1fDkACgttissxY87Y73VPhBsAh
iOPgY75h91Dv+ErgrrEBaz9Ewu1oLh/EJ/iIe+qBCNWLz5pxuU9/vlt4L2zoPfT7BFmGFuWL4IHv
Wd8z+R+6ApnjwpNMyjsEzGiPKMo7JT+zouXpAeG7sT8YlCJPq/fy43qqqFDl+20LTQly9bIuiNzi
0ytff693n6xAcIHE2DrhUSQal5eWgYTs8WNWjetcKVKHGcniHAs2rgiGujk2GUGd1ci1kJ5VpMkq
WwQEGGYZcB8O76tcAiOiWk6OiqsTHgJvi9HxHyK3wEY51PtJDb3muYdb0XZgV4qVYyOKgb86n6No
3w5uFIbYCHfGdW8mKCwIRKAFnxEXuwFjeqk8c6hCn7chSAHHJdvTIteBfILR1mz7UCwpOGWJF6ai
cSFmnzZ8fRw7PAGBcc7bV8w6757PBhJtJAJ93O8emxaJThggR1i1GXA+M9OcnEFI0inickiADwAP
OQQrwtOtm4s92pg/fY35O1Z7zh52elBXHrRg8sq/lpgfxoSf/Gu/AI8qJlIuU29aUd6dGYV8r/CV
N395munt7KZDRtVJCh8bXs4zYF9R3YHSMW/2p6FnMvnllqnO8XVsmxJ4Gw+36636JsVhlP+1PFmt
2rB0ZTH2sz17/ReJeq1CPPsGRJKFzMhtVVqdzVKVU0VCoi19Kcht/H20z2mWCcCFnzxi3zeG0a+b
scBFFg/ZjVyNk5lR0m+qdiMuZy0IO7WiRGFQJXvXnM08IFNvAi0pDCgISYkEU5FH9THkI5cwiRrD
J494ilLgRC5L9CSBJQ1dCfEq4y050N+0g4HamfafXU1qGShIObghABUoSFf1LLq2CDg4W9XOc/Rl
jzNOQ4UdocdAY4fT5Os77YG80kVv4mu6lXAccGMJXhqwHTFAcdEgvY8f4K/vp4fJ1yAJr+92TR4n
3f/LurJXnGaP9ia09gHiZV6M4ZU00cEcnXJ/zlH8vrLl8yc7C9hsLo086W4dEN1Nlw9YGtItdJ2w
CuTa1ixzoIx+11bZ5lVUY06ywaBHml00i7bepDx3p8tok299gb1evoj4SxicZFQ5VeoA6OO20FSP
SAhmKZM1I9DIOr3XRm6xKeF8PvYJ8RqFniOiUBeCbIqJwetwCwLYXjTDzOmJ6z6R0O+6p3NFLg8L
cFnOtrmOZbAqqdBujhzpGSINl8Yv2z8QOJa1wnJmcJhEe1twvnlRV6yUn0IJXih2ruWg5reVs8DX
ECLFujbf/yclfqZUkU4HLGoyNry1ZAQh0CChMEXACICD3pYOIxvADPOBI/Wk1lgeuP889Bc3Z+V+
OAoyC+WmrfB4qBN8tJMgiUbQ3jWSWgQ/K2CfzMhP9LWsyL6RyK+4Svi4JzGE2PU1eiN1QFI9W8io
vt93MQys3aezCm3a2ub+h+lTlRAzSAt/CLf/neCLFX3LzplpLdZ+GbMhofUuVPUCYGE7RADmTdTr
12z8wKQRkfoHyh43wvkrVzv3nk9H03IcIQEoC/nYgOzYHyDhtrfAB8M2z/VKFPQH3SKNmTq5iOZv
5mkLiLtZgjllX+8jujytMN12kraK3Hcz6Svst4xxhzk5EEEDtt/g+T/n0gldESWhyTFEy0Njzhan
pBvHl7DGjUWfAqZhuNQP/iT0Lsw3lEV5r8TcbDnQDz/wycvIqBqDX6SPXhxHVGpbqO6OxAfRQQQC
ayPgurZ4N8tYh5WXDOONBoBqSyLtYZ/FDPFShnTaGaw1p6hu+gCXOUZ/W6wcXb6q/kmM/wEm+ANf
8tyW87CtmEeihZ+1t6tR7XlEOlfN7jw3thoG64VjGfnlRnTA8/IWjc9H51U/3ONVQ+iOmHEQoGat
+0bFXvT+kLDVzj0nrEt6Y5WeqzIVnADO47bcrmhQWHhhHhBiCC14/iwU2JwexXk1ez3j/bm1eE+w
2f/glP6SxmwyBZWeFxsnAkwChZVtQxWeCrTxZHzSiNDYh/fKz1z5rXQ9XgRZX+NJeDr4bWPyHOQ3
7rFjkQY5kdish+EsYngFnbFEOqzDMA90X1UPhr423phoBGyuP1t2mZxUMHX+ZGH6wSWu1w1b5200
JqedevmKAlsWGL64ZfZN/76bxcm6tIdMRzXDCFfF9twLSJWXnVe4dBno8dUPYwLw01NDxFqK/c8a
fpsPJ0ZLSjjhitsv+rjitaVahGp5yhyyhSSJSg5y/reognxP+zxHkk5Ys2diRDA9S42vxKyRiNTL
sclVcrQObCsuITWa2wbPgwBcRlFuMQGSBNxHmoHPOsgfIor32kONT2yC0i5+EAD4qlhZ+r4+URY0
F7y1TAviPrFrWYeM8niu++dWPD3/Dwdczt44IRUjqo6DUsRZDvgfd+//Mg63BTXIaKKCJSQNEQW3
qLnrjacMhvtC9szrzb187EeX0iB/rknOvIGpO+W3CzvaQ88mHf/MGW0w63+0jbvfBxvTV4JrOCQY
3JP5+FdkyrmJgM3az54oDSJ8lQJseNPVmMzxHs/5QWA8BPrSJnRxPr5DjdrhwxCe2iJyJkS8DrJ6
7PzwBsV1/Rc5nExUMRRjj42kTfFbBaqFMuLWXLJIWb1W1acnJ53Thj+DnoyxjkwhIBcZMXfE6+IR
oYhcgM9JnID3H7+XTjbjUX+QhN/cj92dtwRLXKvj+pKKWfp+FtIUjbPwBPwAPCRRn8j5lDYgevph
/wD++50L/9na/7qHSz2AypJxS+Qk98WzyHFk95olgLO+jUZkd4M5m7c9KwNWjwJ27z4JaiH4CtH+
TMYaA4Vn1ZIznWDOSO6CcHL2DZqL2pXfzPUSWXNDbwLAk+xAuVyBTF3u+AfN3/NqndgpMB32j3je
5t9s1RkepUq/6r+SU+JUQDFphOPu0tKLwmVCcJkUTkZNUJd0tje9mnL88lbo3n+nwQSEeHdiTLGq
TCDDloXnTeII3gWgHVJIpHt826m/R5w22GA9o/IdW1HoYqF5pdev66q2m6mzQ7RP1lPdTO2hleSi
s9N9nklxhuydxfRWw2SbYDyPN5RvfBgkYNrJd72sUs26ZiOquW/YFvr7VsFpXvYS1R4MmbzS5xy0
0KRxYEPPTKgmNHnw7Nd9FbVW3bKHYDu1SjB3Lbk4E7qCThYwoiNXL7Vj1mqLl5kpjkz/EXb/mXKw
FtgRbyQhgHZ/zk1UejqS6k9oWNG1ZHuoaUmx1MVgtg9CZJvr8SifQJtspLFSjVbr9pK4lg417NHO
oux4lxzoo0GH2mf8oB9nB/O+82rml9n4bz9b+r9/hi78UVYxhz/XxqPWw0UAIXFONIXc85/Wj6VG
ekMe8aU0YMXfddWcbQi/BoDwpXuZTLtsHaPAX69s30h7M6ma/yhoXk4WDyYnnqRpyX+7+wHaBYrS
Lucj3KjLCOhNkHiTzioYkJl/D6JaRvcBq3rzB9QoYa8h57rvqytXtFsn3aVW5JXdpOGYaTjYQaIe
R/CxllsUcL5GtpJ+B2bjxv+9r1ZtY8Ce9bfpZJCrzqxfrPv1/naYyEuQatLw7Evb743S8ibW1zSx
sBBOyupmvbmb2a4b5R4WUUPjFeHodOiJubI82sxJ2RJubcVqHjVw9/Vi8ccfNiUa5fqHSkzQIZ0+
/sq7qAeHjYhTGexKHGhEiJ+dVFrOFjCEAyHxVu59r0+ri4qg7jCYao5FAfnP74EYunzGgo1PL6a4
fhtsT/2G+OpLM3o/iRDyBPDusAsxZjV3P1zrnZBy1VaAa/4nzrwEeX+F97yuRAucq3J1ymZUt6Of
Ki5kHfhJX7DCg4W79pC0/Uwi3D2k+2sJ3qgtHzzLF1OHvWdolB2R2mo69uXwKsjIH2INNCuqYMiv
HsxGO795DBHLRXWsheyXc0NLdp0LiNx87AC1rW3RkfosXMmiFRH+7G8ZIi/qDMutXnfCFkJwmeqJ
e0+KHR0AhbIzixBcqq3LI1X2RE44my7gddIPYBLdliXg56Om8scsIzNyYwq0LLUQqYX3RpJFkrT1
X8qGjcoHCXf6N6N4VsT8UNcj4TX35MffDhWu1DHspD9HAGqW57OLyc76kTJw45oDwmbso16cu6KE
q9fqJQKuyV+tRHmecIZGiaceHX5MTq3MPuwPjGPBfURQnlOGB9BchssrxqjYplgBUi6rxGYprBeX
Rjm0s2SdbQfjCSz1vjOSdYoTuEibeERvYnwMtznix42xWNI3KPfpwyIZvuxP2dnfE99fPkVsCSES
kOpG54fDYDiDpQYCfbfZeLhAZz/fIpXiQQOqtC1Y6rss5x8aa/ZbUCUqv9ofiFC2sYUfbxkPmO3s
wum6yC05GHCY8clnsBVuBRg6feuaQMU12Uxrh+MDm2fL7sBGcBvCiARESnMCDgXQgfgPq13CoWvb
4MjXX8UBdPw8XmqFqJDcS8RKjoT6nbsQaan6pUTLAtICf/j8oH0d7IH3K7OQLCMsUDIZbrJ4iwgj
7AC5XMsiEayfibyf/rtAIMeWPjZ9hxNojAGK4o8L71+qa9XCIUgGrkMNHHKxFdaPPzLzkNOdof60
sDoAGEM7gwsuu5FTdTFhZB3VLpmdu4871M6CwwgN0D55RdNF7wyg5ItTgAKzvkA/OUO349HkG/ds
sJrtn5fizX19Otb7gzfzje6/OI22d9b0lJ4n7r9iLT8aTNzT5Qjj/pfV1edwGECsxjy7F4cMX5QV
AyK9iW0IdzJ+3NpC0FOAMXBFtXEaIxrIEDvBoZy3HPRXCYbAkfMmG/Jp+QjVqxbGvDBX+dnGJz+i
ws2XoW/UP8d6pmzr8zKWcg/wvaCxOA8e06F67zW2g+MtbnUni+eo+npWKXy8PtdS3tr70daKo1e1
CF5kGPFpL0XO/K4OjmRDFzL6fhvww+bBSRxFvWsBDLOdq5sH3oK8cd0r9o6NcqRfzq+DlKm4Jipe
q7yTcmHITDF39qXQP1dN4VfqF3koIel23AQnGvzyGTPqoIg3qNe/WI0I+wYNsl0UPfP1rQhUXosR
9xNt9I0NRHOBpjBvLbOb2OmM6ivgwYBd8QzQtJZk73KpIOGG6TC3+/os0P2MjqqwzLEceAM7RHvL
QR/xj//Moyi/MLNArtV9fSTut7nUlNQ/xYEx5LBnoYohQ/hM9k+qNu0aDz53WC2B9hf5Pwz1Eua/
OSEHQdVqU10HfO98sWP5fFpQ01I3BaS3Z4ktGYcOx7VLWUBBCJI8e7CZyfiz5NedcTVzRyHJqu1O
eEuIz839ctfvbBZ6lRmby48GiUfUcL84azRM6VfCo9ngGFK47jPYRU9EAVOJyhMluzY5Snk87H5W
OE80PerrNPqlwxVEb7KmC4KOnY+5daryHjEm+kY2MXVW9aBunKtQnxSDdzmmHGQwoYungM6ofFDR
C48AWsrZSW73ZQ58x10ntRMDMWDaOeLyR4t7b/AxsVEE9bvvhPBUoLq/OCFgut11i/ii69NCJNUH
LrFybByrywdsuhaWT7Tudz1KZ5574FDYlfQLNLO31U5soch/5plS+x8bVCLl/nvbemBYm+LAHcVL
bWyCUHgXCk9tZympZdFFa/hEdTDeLYM0QfssjDV0acNXGxlh59aKG2ZYGPBpozkGd1DKBCiPcBQg
h4powkLFqTejOLcXoilpp61Rn0umRmZ+t+ZYOPqTqZm1qNB1LN/vs7dgwwrUdYpZz3hrvk90hmZT
xCSuhpMhlJ/M929WAN/BcIFz6cRRJhcemPHydQTAmAmHF+NlU8HXAo44iIhzAlKUVJtGNIJvg6td
DXFVA5YQIyze2jFK2zAX3ZqyIeYfK+aWx0gX+gd35FPcUY/yILfeIIbtAjwobSiFa9bJeXlXdUlQ
GOocAl7/5PMEsI3gCH7hT3BAfCNW+WY4h6yTVflZygPC+/DUtMfaldUeJFSQ+Zy8cFMzBDLy9Uud
fpTg9IbNWCfX9gpD7l0QMUywxCTzLpdlYyplS7humMZDUTd00zeXvyltQDBCiNvn+iRY7eS2r6py
ZUcVHLv44a/YgDfz6rk8F1HBUagGFRO74fbEr7YZgrgwskH75gFDd5uTBfQdfO1cQqZd6PNKW2zH
x3KljEyunkeTYD0aqeXVgua09BH8tYdt0OBEpEm5vw28EMlUoJHBJYIaWhftWzE/vU6zrUPDnLdi
dDaIhZ/CQaQPi6G/TL1trlplvE6jZHE2FyX1DctEPnyrxCJzJdG4hS7iYzPmmvbW64O8jAyAJpfl
ne2Cv6YwtBpCMI4PJVHaxhJOwvgu44JUNd8BvCfPztX7T3tgXzn/560l2IPK3EGRUhaNvs1UpgxE
RoHbrCS/kMbo9BxYVtBiso6sZaHjeGqivJ+/9C23ty6qjn+3pglyuzk2Pn2VXJQYixCrrB6LPrLc
qcwKecDx/S/bWJmgzyXc4QXvEvJlgR6t83NmknxER3X27XbZLJeNEIlYomjdhywSbc9mBevq+LRm
cQH8xARaB6fTvIqKHTj2v2CV4SNYgWMplD2SnvOJaSBLT9upKUlb229YlWRfcbWNBKXKB756LvnX
2bDZCGVjaSQdfpbQhlgyBrjJ8XJNoO3kdfjx5aLfCSIMvdougfRtlUDMt80ctg+dznmtyjZw1yOO
C0CtmE0WUmJuaaAHpDuoxeUcANMj/fD5moobhswGoC5WYb4xc/QuDOKQd4t7R1XVUCKFteK3lQZS
4G9rqHG8oBrLUkOcD2vc6R9a/N87a9UeXiwRCr75KzIIKaOBxZlz9gjHgnPaIr7MicR/iwmxH4ju
OAUg9jvgPO6MLtwcLifEJLKzInXqblrePds+tXriZTO9jVLlNF9wvPKm21akU5YpeVPh++O7WHGT
321s2PWdZ2rlyyow4qPps6FJWqe22sN7VjsEiR8PIXwim5yuVwwcsQn+nqNgXFyhy84pG8n0RxtV
qphn2LEYD0fbKQZA5QU06QVFVjpgKBqya8ZucDX2KhnROPHoC3tOSnZEUqBBaIdmgTy32G6uWASb
W5D+5yt7MeZXvzRp07QpknVjKDXIOLA+buVnih8+WDxa6HppqDhyLamWAYjq1rzIm6PbwJlN0XoA
JryBW+R3iAw12NSTEWUil9J/f6rMQJBOa1/nYZ+EW1pXGE0zk0nzILfWKPleC7Fg1Q20yp+NUx5T
diybKBdhcBG086cISN/qlmET+vgiQafQWd3jzjIIKjNyPK0iJxRu0pi6dJxJP1fA8gV1TwajWzjL
7IkjeOd6cI4V154gLaSvNHBwK9J1Q5xE2GrTCg8iAzHTo4lEOh2l1gahfGFBYgRWsuFVF9OAePA9
drNGY+keMpvvhmaLAZIZMsnazZL0HgT81dOobRkjDxvFQTr1y9gQp8TfPWumNP8gD8DQ7InNSgnU
NjpK/7QsnsZjqO9bVn/UEDIxSnQrz3A7gRo8BkMpE4jbeYtMfFRWLNPzp78ejKBOUp85AUU6eTHB
NKVnvVETWCCFC4rIC3C8lTVBiBNm7wHRGsllBqm0lwAH0+rpgnycQ57h5W8eZwjFmXmW/CYtdDIq
YAUbpv5y+h03B+6fz9HbTN3vBBOKsP8ET0O40EeEeNEJXWamdYOrjLCg1ELkO4D3X6dvikhvYLUV
uuYDkTWCsQIeLu7am9cG1PX92iP6I7HnmpTrWhHa5y1GRyp7UgXQqf3kRfbPL+Am+8uKWOH6KIZu
oOObBzi7DRCvrXxQiLixxyMvIfJ+UlcgsIaRTTS8hyoyjmOcdYUivPKIDTLfFsn1/sKgyxH4jmDg
pMrrg6r3+GM+vIB6hJkBRvB/8spu9aw7uUUzxxb2fE9rAb5aMnHpAv4YqVeuLIF8lcgB6HDTJxuC
YYVL8X1tMdM2J4WsNj/OYgNxcVERK0fD2q3WloEaNud49yCaiVlthXb+akBR/ZIl+ArNfnoLGAkB
YGsinNJKWYWGZUL2El0caydxWgE+A8vheBPHuzqFM/KuRCk3AF+KVmf5G+decXHSeF9CLeGTFT1E
QK6OqN0ogjUbmi1B2i4z11xu/aVNkwIkbG3ZUvbLm3PezDjSOdFX6q9kRLO6nQanvsRSdYfAQMQi
8XQOxXlvj0zfrssws020kUzOpB3XGEARYpP0uqnuw5FHqTZBQCWd7yBSU+0Ka95lNB0CU+evtXdo
OnBHyqR1fMpWrr7HumfrGYG3omyz9LCgmzyKUq/NBEt6ai39qpfVo3nYmB38PwFrdAkw/eNIFtrL
TSyoRPynqTP/7LT/lZIoKpxRgqDXyKfF2hEYQ3lWVwTVQIkrJsPRV4RxpSJQMixc4Qzqymcy7vcL
S5nGMxyCCHhsQPJx53qerDxKKfuQq+oeLkUTmxBXT7G5eeKVDDXCSe/oPm0PUMcg5J/AOX9aZ61S
LZ5Ej8LbLo+1+iUmLtM8nWRSfRqTeuSShEX1ivdHSZq69CfnWvBPqiWoOOCiG+QIaXKFBrVIrtPG
wVb+ICiprr8Y2XpfRyOMrUPHnjiYRK1lVmyTZTZ7DuIEjMi637rOEReAbWARFTFpWPWmbvAO0q3t
jlK3kFRwSQRM4egqIS69xHkDzU8v2FQdQ2SAuZniIEhdegd5uDaK6V3Fhm/rWkumiQQrDyTqilXe
XOoHRx7tZlvL1OV+mzR7pfVwyKylp38eJp7v0EOhJJis/BkrRSZShN1R2VY72QpzGRNBDVGkOxn7
wWnBpGLhw46UlPc2xqv+UN7csbffoTbZe0Q2q2btHkZqPftm5hSUluF+FUPYw/LwJgogxM0CkndZ
Z21eXA4wWt/M+hNJjkF5yaTTSKz/QZz+vzsEGsWh71gW1fE34bc6Bj71zs4N69pdaDqS6t4AzLlB
b7pAuVGKvXTSjk33fOHQEkgJ8vCbYNpQRCHTtyAmPNCA6Xu4nxO88BRoHEJialAq0MHT9vo60OhI
i8d5HHUcNfkSecocZF7KxxaoJ+Iy9wbfhLvCy+2OSJUjRGDWe1TgeVzOGiPzWmbvXzc6lJXPjb9u
sNti+CWYva0DoqB/DCioWS5DF+V23CzSkeXMXDBNNDmaZbQA+BUxsS784zH8Nfv3j2UL6VPZoKRc
Vp+zGKAeff01EfTSznOF/BN4EGFM3AoIeL7WhFGfgjSNhPF4+HVyXX/7PrOVyXURdBXngOhitJ3Z
Us1WfLqCaIPyYrs/9w60FZIX+k+ApDTkTz1lSaRO1bAtNpfaDIC+XFtTzyKEPKWM7cLeKWChtVKu
Kr/3Xd0TPfr9h7zMNO4Ug6eVWfRjVJLjqUzwbbUJ59QN1vpF0q2+51wCQl1xWcRh6wsaMwGIxoNE
vNafgJZPabwtwnczwuGpbwpRQI2e3NzitPtfGzaKWABrpW3UlNiQ6fdO5BqsHCAqkSiqMGeCTCIQ
1gDoBGSOuhofMEvuOKLZfF1DvWZr44FG0s8Wr4kjJP+f85ZmjLEPUFLuc7FgbZnpgxogQSYAr/q4
8mZfm0McOWHZisZJ9FtAK7Segz2KwtUVICrtNm3PRpVH2ktJcnBS6bglEqcCpK2A7de1Iq+YBAyj
QUSTLoL45UiG9IzxAsdqNwxf7OOJRqtErb77gxjkibuqy2Rb3e7lS0ozWkHdyUmpzLphU2KkUQxe
vizNWpIkXFfG6nqhYE6yfMSOoP4Bfnu7h2rG6vb1SxgjowyEtWAzsd5CoZUBlv8DCj8mIQ8++KSp
LtXw5WlqBytGfXPIUW9c1kvKa2z2ZmOsJNf7lpDKAZclCsIPhbA0UkRFbdfV4QJTArH/w3VjYd8e
wYht9TYU39joJAAZR6dwpG6Ntq+kMSx1EauO4YO+GjVLzTBSnBcZeguXbltdEBoi3xlLfvwByMez
tkjJqh0qq7alm9fm6XkLnPDweThuih15Q+TBVQaUukOveyq8U+YW9/8i1iHSytRpk735bH35QL3f
Raswk7FDfcqCi3BHvh+7YxJvX275cAxK+9QsqFyFB6iiR3DU2z8pebKaZbOY1salxyaZSXuaHFL8
TsXzHgXT06rsc7X2scx8eWMLMV4uv1iv27YhJ2nQ7xPzXp3FewqZXQuT4KDsahVqdiLx8jiYqTpW
1Q9izqiOg6s2C81aWJl874WKArxgRNN+iZThdkvWDG9qkyqKie6t+NCauHEnUdexxYA67BHmnWJT
0vRjNyLf+2P+sMk6x2b1f9d//pPnEkgO9hohwuWFeMeOpw8n7D/xDnmEUzOgN/mDlX5TSFzBkOP6
6UaWQe8AxXRr0kk51tYy8fkxeW8nCV64KlIai4vWqNizPhKpaPVGz8u8l6Bp++RhLK2tMCFmUqdM
HcJbEkzna20b265ZLrOji2kZU46uXBOJvbcu5RMgrlhQzv1ApIptS8jyDcuSsS0/No53OkN8cXPc
e1aWHAgvk28r8Oyg+Cs5B/vd0AG2N+5kUgyz/yQyAn1nIEjEDpw4eGbVr6x+jWGM4/udsjwbkB2a
pMbovqizpTz5zyul8eIZQO66yLQtJVkarAnY3Zb+vOBlfKKd8G+etM47y/gNV0g6mauD98BcIB4M
Sl7kLabAYocA07p0PlCFEldBkBRkBja7LCHZkNRiUcANdVGWIDWhXP6URZawyngzdXCcZgj/D6Ug
9Q/c4gR3yY6zUmtsZZnd3Bq7ItDw8f3QWjCXEuq5sCboYwJuWpJR5UsV4WQ2w9QdL2eUuZVbcYKj
HZG6EIR/6cJ1loIjrHNc1BCUadEOFj9p0sgEX99Z8M4nmYjinukfYw5nzQuxjZ8jam//65g3DoGA
w/bSCZ89Y6SyAdzyQm8DL6uJJXLVYHg7n8HMG2mwj9V1jups5aCCY6Z4GYjmr5mFZxSyjFiNh8hA
29rWY871+toIWDEk30M8Gbv24hTlzlJ5C13TjPzyUuWuTU3jkN4cj/+Fjpyp25+///dWVn9Qj/xh
C7t9cJsyj/RDs2Xo3lN1JjO2eLrcecZ/A0CvPxnMDOy3qboa2w3T5Ent3O5q92AS472LMPAjx5j5
fgJVO8ddA97hxZ4FF0n22l+0eZAhE5bjylu8N7z2Y9+4SJdmGY2GlaBjIP0R0rt44Q615rDAqaoA
xBz3TqImd4uKhRV6eDbJlCI/SqXh56LhZFRQ8ZCHU6q2Ozz+BBvdfvhXPkUDIsvLGlF3DLhfcYZ/
lYVleIbfcc46XlwBFxF7WNQI2MAD50oSRmFfJ6PPfPKPRpgjLty0iPkEmDu3WX3u7CBJ8mdsiLSW
jElze1X7d8uWlwVzYs5U+GXuHGxto7MWtvMWqdq0dl6niIrOMY8yTwaYi5+FIp4X+KzyEV8cPo5Q
HqccDmb5ooINwXfaDA2IM8AB1X5QjgpnIvnK7c6gvHF6iDk7NQDH8P+BqTtvVf0DiK7n+Q6zzYuE
u6ELjVITE7H06VuravXlLI0epfNErEGPePuU4TlvyZO71/uvtYDBrDQ6u9rKYbWyNWR6jhIP3wZE
BO2sT6obq6KiLMmdJR5PqzEvfmbt7CYu8yT6la8uPB24ji4KkSle7gNmgoLm5irNRB2HATczHCcZ
tLQKMeHv/rWoZJBYV5r2dNclTneJhlAaUKYJrvMkWZfTWt0ZOesnT0TZSVnGBvuU9vB48YFHdObm
Q/EN3MQrOaHyvJGRxXS/Yl0/Bdpu2rvlTFU3AFHtSsUWx2EKnL8u2r+ui1GXrtmx5O1Es9s30VS/
ClIAHWCXfrpOTfcwJWklj2/HUI478k+vVbQslAbrZw33yTzIUaXNrP16K1IuGhyYa3vwsDjR4FbT
86wNQrRrfhjyW4pbA/8J4ypM2uOJCnbj8UK56VpMuYPrU9WReAXr3fS1BiJVQAfH0CMUAFte+ne1
peDAaYBCLVQS5nAlX3ZepFdILKsQEcYYBR7cQAx0aumUjhQSyFp7h3Iohhkyetz7nMLbqQztWs0w
kAwCaTAjJLPIS0tMhH7w1zEfJdzzlzt6nZcJVtv+mrgz9M4Wj1JCicCwuPfTbkzUuMHCu7BSkLia
c79wwOfXqPuAD1LjajSZFj4vO/m21XdNCslhpKhjZwMmw/Jjt0eSBpLzvYSkZzg32IbL3FRe53xF
J6QlnFz3IMVYaeYNEm9YtcRq00GfjZmWyVFQzK0KiD28I/ft+3XIQSbVLJVbQW7PClvYPwbQkSj/
37dk1HU2rQVszEBzV69MCDrDFijoQTLo+sRFLvdAi1RK7bP+lRfMLLv5CtVyJPL1kJscCs9JvV6e
JQVgVzoIG6go3ficJNSQCGEOpCu/OLddpbyNSaZgV21tewWeqfeBFyE4SCINC2FhF1dCYo+mnPAz
zPnLY+fhGQRalBvzU59NsJ2mQeayQfyFWmkaZF/hetdebbRwBFBX0ernORueHtRGuPkEu105KWHV
Guj8IN029Unhm9MYTtq9UMVRtOjFmu9vrc3acNIj8AOWzqcEIXyH9RBowH6ISd+azjm2Q7KDMfha
Xyeu81TZUFr+HSCl3Chl06LbtrABpn3rg4w8Pxf7t13OEyKg+RU3FmnZxwsjAGB0p5ELcgGnRUPK
CSl2T5FPMHNa5Qvvt5vU32OMvAnqLDycq8NEX6hRsIw5O7EtxgPGrrjdwOBeVG4x/+Vyk/7sZU4J
wQ5GRqRSFW3kiiWUDqkRvncCs8sA8lSWlqrLLGPX8I5BBOibboVJzga8L+aXVF1ycmoDhyJVbSen
I2Rs0VK/NpgErHy/llMe49Zk6wJG0/Jn3ltVvV1t/C5ez2/uvVOp4AOE/xnXFe/l7djILH70a+kb
oUUKoDevLzyfHnaG6ixtv4e/GhsWybsLXJ+wH/nGf6gyKlra57xhLULd4gjM/HnIuFhhprXOGpQ6
tYbAEM5sExrszGNld8VvZnY0osUYTnhgJsF4AgxHl9c0xsD68NU/0DQsBJvbuVxy+vlt7eptUXOZ
iltZSW+OTCIz1ZjTB7wgMJ0SAwf+YdNEYl8MoS5YJaryNwin31I5VLD5ew1hZX2e0vOP0lQiYytz
FKx9JzEjlLCc8ZAfXx8AYrnnbu7dd7+qdNTnzMbgpK2Ij19KNiQh4/IM9OX4HB6teR1jac6ZCqfy
QZSyYJniJos9woHoAoO1uc041oVLgjhrx1fUEB5fgU4XI3Oa7kiHbvDOwwqGWHX0aIqGwysbggYq
E5Mjv+XIYz0c4ZJTzfaKJO95x+ib2kBjjQVfadq4P+XZz9jwRaB6Q+/zQgdoSXilz5GpbQXVP54a
l+kldCDrXuYEtRhA/3IaZOYFOymifrIPJKHlvPXAUz7RjVQaHl11kIcxNwHHeI6wxpO6apNpytiJ
OG03m3vijOb5afbh3NQDBJGvEN9MWGh6FCc53L+XE+eSSFsGxkIl6WmTCqM4oyIWdbs2UMH+JJgo
HK6XUnprW4sddlJ+p9vmlBDjUqD7J/kXsEUyMW1fWVkz1bOqg6Y7QGKRnk9hrNB83lJBVQF9a58G
ZN/COhYmjWpnGzg8J1wf/EGle+kn2rKTnUjzaOQsenlm5xX/WHspyOvR2Y+GoMnWAPfZVgOe1kn9
0uTEZW0P/d8H84uKMo9QOLnJUnBVEBtMg2pfq6L2t5VoemsKxfz8nT3YFcE1ZUY3rFqkzaJ6Blta
3VR9v12VXDZYbTURD8ly5+LKeGgEVh/Y/aYycPeEVsZai8ULlRRfBKHP6wSxASvKxmluwXs9Wzue
3RlOSSCTroFb3Up0BRk6SiHsV2WyKyW8362qjT4KY9RZsmqJX8npK4dgAJp6tgGTnzN0zbieMrLt
KjUjYKI7lFyDpBKrY178wyIOZ8Fy4ap5yvXbgvMci41Zuwr6n0kffvULvyjaSOK4PeRkKf6MX9C2
MFBOkfJ/G3PVbLSPBG7I3UWI+BK6XMvl2stiWIHQd1vK8i2dVVsYG7yXKZQtLS3dIO3SVelOKNxX
z6bQKJsQ/BlBPcglIjuwinztQAIuAQzNWYrl0H5e2oLOPnubc1C4B2ZJbzNNmZWiYufs1e906QdN
JAnApLID7LR5pWYUFmvQGn2r7w5cK+qHs/qv3g0EdgciMqqkn0a9+PDv8BDGSlFbDoYYQXwUmJJn
qjOO2fENMBcS9IRwEic2INjahgYmfArkIMXVqPf2k9AlyE0Ie0OEQTrVVS36R8nv3YGYIpIb0/RR
UVzvQ7DUJtE0+i2UugCORubKXQpIQ09X0r5OEJew7t9oVtRgT3tD6693f04k2ym0geIgvpiRsEv2
8qrdKJjCNR8Y/PuEiChm//4plHgK54MI1lrkhXycYXFBmaYD/Uw/XUQ2+nqACXh4MmevYybxU5wt
vU9Ubw7paXy6cN73KayPv/SNawA0p51BLwTr0+/n0lUdGUV2wjxIHQH90r9wL5tHSZnX16W5NVf9
fzgZ+9sviHL9C0WjHIy8akFkfwqx/7QnwV5kzVMvFZPgT2biW5eQ72kM4hpm9DGh1Fe5cvMez1VL
WpRhwJGCyV4+LHZgHisiHsRjxFQl3fAf64WZ1YvFKfpFLWkj8qCkI84OKGIBzQxF5ZC+NXXxuhx0
ushyR/EQXMFl6R2FEYufy2uF28RDXsAjPqd5aCmv+dHz5CdpJZB3zy9UED6PkZym+63vxMR1+OOd
hXWyfxpDo9qtPrkOLZNnZ5z3AVVGRGnhV/6Js8wFd0v8cGokZujbWlqQOoSl7Izw0eTDh6Nirbme
Y+jJmMAfS7bO4y9yLDbqFQgfz/bfH4vV2tUSZceLAEFOjnMiVWefDHpmwRIsjAaLOt5kCbSu7rQk
WVZVnMAOwE8elcW9le94sGsO1rzXZkAKcOfVwikbrCmXsWkgTDDrdEgz47caKzvfIx1m3FSqBcmr
CTzWjnLXB++slLeqRCFxxqtZeBGLtlwSfDQaQhQofB14QlHJrG/NCcLbwCHH35gCKuQb7XAI98/l
Vvs1K6hHAyDfN5PArk19PCh9gzMHxLG1rPrWsv+86wqc9fyHjdvDZvlPIwd/cn/qi0JuImg1frWs
4FIWvzEUj/Zwkht732MWHNK7hAKwqHZnjvz3ycOxnA1fD0MvhZEPsHix+Xxb9UVo/rWgyUxMy9bi
NAYVN0G9I0Cl2gOyQtPTb2HZ0AHw0B1lcFLPgd8sD1+uEgOWMz+wFyyiFOqdxrUmwLU1nDoj3NWl
cGHTchwMxHaZEhk6/58VaXvBbqQsUPI1oe1V85XEbOrE1eJ2SbKOHcTnI9aOSC+gADVJoJ/H9Rv0
ZHgFJrajw+AYs+n8BkA0ijL0nSrqv5/dLdsdWWddryp9JlKS5hSqBmLu8mtN+lGaKkjLlK4JZsf+
9gRtIFg7fUKwR7EFHZh22bGV4aPiqMXKnH0hRCxxexr8Dv15Sl5Y56HXsoVPfQBUp7JyZXGeFyDp
gkjlhLPhwyFle6kn70vxRlHUasTfSZXEA6oBTUKRMVxTFi3F1zoDV8p2ZWbgKIyi/KZUMpkhye62
6UomjOFuKlymI3h5keqJUafX2jegpdRoSqG2awty4T5PjkZCpsJHi4C8ayDkKogjYg9+R2qkZMgP
lJmKselAMsrFyKBTI6nzdzDHQ+ofk5mpyrAG+6B8yLDs+jcaMSZEtu3wPHhNpxTKa2DbcbZWahN8
dpzU4pyZmZkob/mrdWg6AFrZnxmEO9k7BFwAEr3NgVcaA3pKACx32XeRV0RE3i9kUl0eL+79Dpnw
XPnXsCqAH2E/NArUrM1oRSWGs81sMLGW9PapOSdxSbe7mRDHQnm3VY6Z/YKqX6q3xtG4jhgD4Ksc
MCF6DwLfHOeEoZUWHuaO794q6CL8ItqkhVASVR37sAQCGaJSSOepFYhsjatYsPjk3L7TVbkSr0cC
bzAXqSba+5twBj4AqI42JhXYCzBO61juKqB1bokHfhDgXV7YB7RImO/+WOuuf6ZTkBaLVPODIgUu
HreEHnf4m4aLokgNU5/ifqZM1ylij5jLzJBcF9hHOoNrstP31iU0j5cunrK6V+t5fbEcu7LciTVJ
AP+grNRH5je3wR344F5VdO7g0L/xSLip9lBD8ZKFxbNkKqjCJ4cFsSMlSlCWsWW3vFuLbhOzXaU4
1l7x1EM0gCJjntV/g+9NcrMHsJgYMU7DIzaRXtgWoJxsgX8iLBPC/2gEVMoW3t6KPqTlEHfTdN8A
ObGxME2E5KmXIY6xJ14U0b/PlzAuKvoV4R8Dba9h6RGeo3I98OGirMyNOCL5PB/hOQ48/2G4v+kt
SczGu822ITCz3RYDv+aBlzYz/uuoWxOGG7WGj8mstjaihDE40oNi0tpGQN9/F+WStb7Pc61X/Y+J
Ns1V1t22vOA+t0nYCw5UvTPw4nKRv7T2o4JykTsaAH6RcG+gX87rTVlzm/kh9UDqwKns4KXNNasw
wFZZFA7rH2dL9SrA6a6E9UC2D1GfK7Uvw139Q1koAySJtQYFpiIBSSsmgiY9wdekMMtewsDLwxTU
JpFJO0SVd8Jp5DUocloZgjj3YUk6jfK+n38koIhi4faYuPDY2PUti6ZLPZHVx7yaql6Lg8wqj/co
NDjg9H4Jwwzk6W6cZlK4lQu+mxzWFTYhHMUln4AiSX/lFM3qW+oHcD7HcDBHmYekG+mbDOSY5ffw
ByFDNi91ZYse+oDbdGD2oHzM2Xnmot5roay3PslDD48AVDAZOZ5onZC9HyADakTLEX5wTZLIxto+
VHK57d78OK8DVlKl3O2rEB3957eA7Dcm++5dDPKZ0LifUkqap/44IeNMOCyNq7vZMBMPvYNNVG2p
tyvE7sf72xht0KWzWElmy/X5jiynDLnvwBda1dSUJ4QTniwUYRDpl3OdPGpzO+MT6Fjw8J8v50Ba
QWWosC1HH3JA/zP0SxBoMOTEXRCgHyRL3LDGOX0rID2QGq2m4Dj8SvQgJJgXBripn9AHoXHYeveH
zkNubIaS2xcsoYcWZw1HvLeDsryTelNCchlZj7Nw619QqdD8IGX6CUL69A6ib7KDW7Rf9SQ5HJgc
ESanuiRXtDtaALu/63JaPxwTSnb7PFoAL1FQjcZ4/MZ+gzH611A9yWE1IwH169NTEJIay5g3tknQ
9cd3RrymAKeSoy7VUO0ajlFMLbki1KziXtJ6+djzvQnou/okqGUlN/Nw0BmOBcazxymNnNOJmWje
fKRtONSkaL0450pB5lu1f860DY+BKhyZ6Af0Brwh8H8QWF0YXat1FqKP3RGfxYGgg3QLbVUAxubf
f/rIDnnrhIA5PRLr3UizVoydctxLl1XAYeJL24UOweKUMgwg632TzEbtwp0tW0Iv30zcpuUAPlpS
R9tU/Ixqq9ectA7Xjex8vW43OHR7Mm6i5y00SLtP+k4szX2U/z7bTgGqfyLTfW2gO/hv4k7znd7k
Ed5n4614QJcEgdLTUdPwGrfZMc/XA0qtzl0MM6IAykeOHFMlD5BVNQ8OgYOkoM42eax2Q3ylC5oZ
59vagfk/6KulMamUWRFZRnsXLVnRLxnO1uDaHwhmcxBI/t94NRyupgKPPrGq0ClcdvvEMdUHtG0r
MZrXyXyF6lOJJtmCyZw3aTNuBWugOLPGSjll2MYwn650S7MDH7ld5If59BgnSahcA7tjal407YO0
VFTjxC2x22Dy7o5hK5n+O7McsCh/63on0OS30b5OJFI4TvGAUAxUNorcwjweMH7xpekzS/uoBdxp
Pm0dNEGkgq1igQ8DBgCK2TGoa/4PelfqLU2+qffnCy/Pa3ZcdxTVkHSBvKZZEUeHCMbH55Eds55h
K0N+0nd4h0yaSpwf9DNzCkXdKn0P74CRcP35g8mnPzDetMd3Q5R4pIXiNsV1xtYTcuZH2OPOgiCs
BAvz3XCtKLlT7/WHV/wIBjMXoyt8MXSygxsANGCZYH2voPyAkS/aWpy76xwn/Fy1qcILc/A3NToX
aF9qImkvn8uUVbStl8qNvovv/fg3fomxEpZW+jHK/CDYi7uqPkiiuSmicqFNev1J2PeuwmxleDpu
q1ynHVgtDnGRPZ1FT6VI4/cMN9fVl1troXtKRYyen4HVGrX18PiX30qNXCWCh2VtuLGNmvaWbjNL
uxX54Z6NOtAdC/dukEpl+jJa53vporwzKvGJmrTBSbBSTkfLb2zphzeNz7OundAV8LgUrGML1RuB
65RbOSbsEPtjNRD0ds0WoJ7828ywJnB0O0yH0CqFzt8Pu9+No2YqDxZVzpnrE8JzsCFi2XSikewA
HMnSsXHkCF2EX7cckTyCmkrBKxDxUOk84GkfT20/buWChSjAHAM6RMUmmyFD6bcZ2+4ad9tiGolB
DLpfrL7NPO0lI5jwhVKpgP0mZmcLD/vpP68/cFWslsLebr6GmmXnZRaw2EsLIeauLPaO3FRr/rlo
qN9KEgMiQg8A0uQleoPktTNNIzkzNcgjN/wjUWLGywP1Z2X0GELuGoTU6NpVFr+zdePb7iJXdIcj
zEbOKSA1ftgo+SUTCFIGiMV3U+E5RVjJ17dOblgDqoPU9hCrM/76LXazjFDpClJk6lLYQiXbAa/x
R+uoNbw/116gFQFFwA7s1IGU4gRlqakFkbLl0K/ofv3S8H982cMxgD/c7VwRZ/1ZxBJc4/azdn1T
qZiF38tzr5wUlw2niBp5UAqFNd/QU40KfD9uAhWwoKmY3hVTugvVATWQ4JmA/FluCsNWj34v1ehu
EIWTHBpmxqDMhF5o1JtGICbYXTd3wk0p3m+qPngVQe2d83vVxNfD3qXlZteyhTyXUPTh/AV96WuK
vBS7DRksyyE+Cl6QEPq5ljDTC0LotATjQhGGJufo800ILXoJvMAyxV3IPijrR7yqhSTyUqCDYdgb
KbNBo6kK7NgWjVK/5uCGRj6Tjy6XsApMmnvTVtZjP/Viq868oCZVBN6LJOsuPHp4EQYy2/K0R0UM
L6XmUK+ch6gyU377Z4sasnxuviPpdnc3gTVIAqnN7Q4gIgMF+9F6/5XDDMnWsksyxV5dZieC2tGf
j0jcZ3HxvOIdROKHI+bIAeIsI/v1j0mF/pwwhVBPfrxpksIYqSLvjyYTRjYgALyhjSkk/nYQ7esj
ByQrEjGY76Pmp93V0997W2Hlu76gMLoFK71AcWaUARHpMcgCsES04YV+22dvimdiofdlCfZqFIDs
xvV4RNoI3oST2JBkDxjHvGy4vAhI1hcVJRUYANDlOL4hOD3eEIv2ZK783pEpw3F3l+k47nYs4HkY
M6BE69s7GUlDSQCgTNPOJmC4EQq2M3QAhZiMrOVULT3ti7AFYhgv7zlnP8aOqIfdq5JTuFlZcN/7
3J95MGrzxP79W5LOyCtJfajhTfdmjngsZjRcOygaKvzNePbHb0jQqd7JnzI7hyPdweUFOYUl2ok7
fRICDSIIcVhtjrntMfrOedbm/sWWt1nBAI1OwsKSVEHo3pS6t/6QrFmOyJtxJytXAvI8OS6HpxiI
82u9Zs2ZZJhOcF/hMM4A/o4M3LyBuOcvhMKePuy6mNZeuzGYMPZ/8+qY1W5uNdfng/VrT2b7S3aK
bFnqLCu1wvhZ/ZGEO8jkVuDcVw3SJp+9ea2rnigkzF9B9mbH1ru1S3jOMRHkP+0e0aY9v7alLzuF
lH4PH5JwjZUwniZLTqat22KTelHfFdoqvVfAvYUdflapkURHA4Cdht4FeW47FtcMbRqitmGzXtaA
sqmTnzxGCxKjFP8tfDXsoPMhvyD4zg1A5i3ovvSrpqlgQQi5/jmnrMC1pbG0cH5yOhiiFd+IrP5f
Mazq4ggYFhg/edRfuemwIemP1LAGXyEJgqItNdx3jFN1YXNU9IZdqLmkyNq2x01mnCdbbItEVcXg
rxtA1cbNu58x7n5uvm/cgFf0R2q5JLwiDfE34UXmwPM42cswCMpGm+pML19GMeLmwjgJEOZULBNA
QfiuXDjVwp2Dk9cCFrYL9wh64q+l9II/osych1KN1wi6bHYDGG43ttkamGfOXRDA6PLBNg528vPL
LHg38WweaO1/Y8PWHedCCRGOSmzP9+yMlvG7vsn7QM0USp1M5nmY8ep5xWP9+3nEBCm2DaGYOz2Q
fsofLoWeDUdnIl/kdbBnEsVUqBuziPEX4I4AU9QLhX7WXU4teOqHt7heeG3H5iQqWxtdQUqbpKy4
sr2+5EZTwTZvne83hoAG0aCtXthBLt8SKMzMxGg7cuxXSUhqm2oOVJI2QB8tW6+l9FMzcYyuGQLS
m9tnQ4qLvdFzq6/73RsHJ5mIxO31KP7a9jhb1uaz+HaSoWNpDTRFDcvLnp/sUJRlNIUVO/1RegqP
G+vMzQiFWkHmpvETxH9o6RRuEnIFajWjpwMoCMC/u2C/l1TdRbJKLUxpoE4ncrD+SWPwBbfLhJ+G
EkssftYRClnMAvrIDmoMc5J343IiDI2u1C8zl8i3pfe1rSPZZgBwcdx1qcEdeLPuQKq2RrHa7Ta+
e9rmlo/ZXF3IIUGJH4Xzs2j5tXQXh4XSUYZQNKCWnqSE3p5RwO0pDgYKSX/Ubky9XnQaAF9qOu9Q
WSv5JrI+NpH9NvpGZ/sm7ffhx9dIoTelOawh/JbTnOvnwvJunJIdbEekVl916YSfUmax9dY9jWa6
Vewbq2BWaILnBA+QQF+i6Satcu4bL0HdtICW4xsfxTOnNDocVwuEZ3HHtn0KuGABB/uoHWBp/BxC
NOzhkFmRxY/21Bf3PV6cdOkt3w3W4h40LjrEyi2l/hKGuthsrK+c6tt9cmboPGa8f88NxEfMtfSc
mC0gKvAW6zdZXXoQzlY+DtFtgP/pTqG3VfTndxiPo6Ws/YOhj46wujsWn366xdjIdT3hGvfnmyFu
YiHcZS3ocMALEnhD0+E8BrKKlaeFEpE0SispEPsjd+FT0odJ1uGukpQH85mrPWDDVjlA8yY+fGp9
ubojx/NmONpJtL1ZI82KEXFjiImDyzh76Z35sloJcL5OFcdJplL4+JUaJ1KuNYYoVTh3lQboEJOZ
5jZc656heDAwsljqyUZEbJT8X7TOc6GzLbXebAQ/gJzMFyFB1eKA3XVHduEWgeboanF3xRD3U3tz
EK8B/iPXgnzB4b6wKdBTYevEgNC/1io8lELVm5uB4AkIk8sgtynrmx8spG8nAj17dMZtL1vtG8jB
jm6r3JCR0Qckl3cOqPjHcPScOUqCK1Ag/DdEcsykdLb91WSgUtfE/FqPTB3hc0X9Qqotul2scvH1
YO8hHzjsn7HbU2X7okJISfKdab9p6HPHLosXVg2UeFXk+Li+jPslMVKQozSa3Zdyoo6K/bBDP3YO
Zlcm4rkrjHlyhLWS8HPgmu6GD0RQo8v6dBmCKEBwbqNI9nkN7JIhOzBVbjzqn1dtOGarU0MRLpNU
GL2t43K+zQ1/50YSRtGktcW3gtvYjdUXhCoUiHdZU6XXI2PYDYINHQkI+k8i72IigNysF4M+HEGP
4dE7QVo7aznHMEiw0GIjNh4A0oxaxxXS20x0WCFA53UlSG+cNs+PRXxSIcu2m3PQmeFjkV3I+O3K
Pv9VXEycEGhkUaBhHfdSMTlnky4WeFscOBsZTNjD3q3UBXaPdGsDLevj5BwRBN19gsgwvR8Q15kV
tKNGBkp4UZGZw2dIuHnoOCLvFntZf6Er9n/O68TzybROhZsAv1VaH2TY123s3dvxnVPjry9e8Fds
h3SGvgVL0LUjzHJePyk9zF9ecACOyP7KMC0N5v2jaE9UmLKy15cFUJnIFjGzJJ04YOQGLLQWL44Y
2yd1LPzGLSNcYUf8EqIEOSd+D3EiC1xxJ43TWb69wal8Dhju3DPHIvvkBL/ClygFs4u8GexWE6ue
SejJhh1CA8eSnj14k6WBEcjzTOHjxvhGBOUPIGXubdU9s/iWJjsKos5hh7f75l/plVvIlrZiDXjv
/iLvGrWiJVdnY4unzFRrK0hRWdwsHNCa83BLv7Si7CRPnhUOQBiYgq1Uod3kRQHpoLCesfJkKliG
BpXDvfQYrzKcR0Lb2vQYt1n32MqIkyoLB8CskQ8gJA5+3rEqRyvctKAaQyMm7nQVX8XEG0lPzYbZ
oCZ//DkWV2O/NTG0iDLjcZJej/8cW7zqclIQjtKrmEdlEYIpmDe9QkgMtjnyI/K9KpJZUAQvc7O/
pI6ochWiclgAOYOST+Z5cs109pR5ZXujfza4Clw5MfqJXw5RpbT9dv44VJL83ogoCUM72y6Gj5rS
8bLXYKP20naD9vOtm9989jSM6/okS2hSaZu6STBiFU+bZGpq+gFrca+PO7RD3HZtgo2gKtwNm5Z4
FS68NQbdzk4YGJwHlTPmVuuSVfnDvC2opIPJORmRwknGyxjinAS2g+wL9raJDTt2YoM2MfTcLThl
mc3eGoYAr2wLDbI+asDzYghUruot3gdY0NXQJhOaSJJXYs2y/k8uJLbOFFEyUaglwWKUzMbUN5nn
cRCHz4iElQWfNpQR006TtcVIodLGqzrQplKsEo5tJW3nS7b1ZJ76zrespTJ4vrjsNwCYcm6q9fw8
9M2LUyUuRAVYpIUo7Rj9DZd6x1ZrkUlV/vkLrBaarJP2iE9EbhYkWwNKGby1CmGuWTifZWri7Luc
FEtEcYA5mQrYgGRNiNL9cAzDc0drRRrCf4iQmOLJXMFsBA2HhcunUj6CcvIE5voBgcghrvpU+/1y
14S7T1iAu2kZ2x0LJi10kAaZPQafvqroHvO2uO6LNB0oXsVibxXTOwC4w0tByobaWkb0kCYLj0XS
uQsgJSu8Fy+qKJBkWEpAS7WNgrKtq4ecBdGRORxh06g165wyemZq+11FMGdl88ty8/CjscpfvdIY
aAxPb7PwLWKQGCemibIpK6l9mmN5/KMDJaDK41eMzn6G9eNmfVmPCc0BJx8HMCGTgd1zVKhC5GbG
FgSw8vCmY0HVT8jRKigNCn7cWo8g7ndxKa6F/6HdAofxyW0+3S+gyOEyW/T6MpPHnayFbgYN7MSV
L8wS3XE5lMG3yUM0gk/eWp0q2Hpg7hs52hrEyypLL/N8vi4Q/0M9km/8ZxrUkw9umJmjpZ0bJU/V
HKf+JGIU7O22M98qU6RqGrxcxzXOgdUkn4/tRh53FSKcmvKYB0O1svNDrcykZSiY5Kyi1CTACheZ
V9KjDkOZEzSjnIJtwW0XkTeO6r8CjOUIlMpjYfHpI8dGcAkl5Xkjjv9SjRXaLonrqhKz/WrRdIdm
rWjLlOms70gP5NJunCf18NAA86bB8pZZ9nWazyE0aODvX08zpUGFAb88JBKOI3/rqzGqTh18fczY
sxoYJvXeyGMWTTjqbBrEeZLNKgkKNd0OEd1SmwQn74SAw4miTClFu+agOIm5rhm+hg3RbaGg8q58
V74sOmQ3V1bRuIZ44lk0Sfd4hSQBlz+jYW/sh0y4Vp1ypYwaIT8/Jbh4/ra0RClcAt3KnN2rqznY
2gA3pjyGbF22SHAEhpfbRmCA7dYHCUpOfZV6SXKun5oSnPLEUu14hsotPPBsQ8xry54FBryoS767
yRIX+4Qx0rFPilSL6sK473O0f6mw9Rc91Fac+b/B1QJV773ZjRQgH1N74+1xOQJOKbmeM3qdeq/k
c0hDFgMHf8pwzbGjE2XBKo/kBXe55urnkLBDRcoxsTgGMnNUxGwyY9xOreIC9w+p4d8tGwJ5xBVY
UIbEsyibn+063lB+4fcLEbvl7T2QTzFocj84Ay0c4QVxa+dIkk6QApZRQ3BLr48gUD+7Iq2Sur5+
Ok3K5U8jtDOmYz1vtlDlesqz0mgFSZZJA8MBH8XO3zh435PSaVkzejIr6bH0P/OTHs8KR9s74Bol
JCOW2W8TpVrjtqchy3KtV5AVIaMOr+IiTy89o76KYaLY3Z2bl7yUXtCqnlndAxtrQQdN1DsS5Gph
D0b3kfmmlYm6Su6rSVKeiN8ExClrNx3JCcpswb7DpNsPHO4klybGWlLlZqWOf8uVqX9bAIkq+0n9
L8QT9wdi50tPNG6WSH+SDmgfroUwbdiDcS1QRBTese2RDhqkircVUniMJOzTAXAjVMo6wb0xyrwu
rBeIQw3Ea1pK2MB4C9LglR0aV8/ySFb3OBMG2oSELEn6JzCXjaSRVTplCxOQJN0QSaYU7VpT9Ph4
2WBQJxv6jOYUMAq8hAtiw3C5UE4qQewyq+ur+DfwPdJwVsuRn40X7hqokaJbrO/fQcCnWoJ1ld7Z
+c8BXoAkveJ/14ZHiH3XD4k03nnQKyJbQxyD/W21Rfg36WBK7cdf8yEvpRBaM25YvrdRs3F1km6f
XGibvSDMcsv80JW8dwRah7Umnllu8b9uWKNNrdAn5gEqm6k/qWodgkHKDzMSSLwSRxmJATItuSqA
yM4U85mDWgMQcIow9CVjM5EaD6JrApXo68ZTkv7S47r0S98y7wihciIseuWFGHl7jbu27IfUUKJ0
uHANifVq56D9YBzoJTkn1iFqziR41uejWMgyil2DSLJzSXMde4o2kyY6xOzBPrxKke0g+FCSRN6l
bk4OqNn60p2SeOuXYXWlXyXKQk1AB57CwW6AmYRyZpSRQ+mQkJybzQGyROqUU1q+0IWH49mdDNmq
W/c8WHgHq5k4HetF3lixt3H8wP49arzw9eTMrIbFGcz97r9Q0CeGpjf6U/JUhdg+tDYe6F5d4IBQ
0efS44j8WD92KpkRvoFOjq63/L8SMN0BLd2/Yv6tFzMQFDh/sH+zegL1TpelqmzeIHFD6O4hKWaD
XtVlHWCDHvd8ny4wLsipfrln1AiMcaP90QAjVmY2PMf2xQ+oXBqguPgqTfZbcG9KtT2hU4dSdm+G
GkUFY+cAwxUxjwaRgxITy/sSNbYc+F0itI3tlh99oBzw/OAUaD37D7Dn9HeODFv/RNodREQ1mk6P
d/U15K26Gmn8thhlTNnT3zJ8GfHgLeTtmJZx/YWD4DBPSlsdg/qKpg2KahITXFIBt4vCsb7ihoUF
4xgBua1Izw2aIBA3+bvoQ6iSbAlwEDDkk977F721s6IRx5Ya7MeQPKLzqM/3Eq+JnZmzgU+DurC9
ibicxly0DiBryDGIV+2+rELEE5jwZlHqv5SearWGzUSiYtHTtdhp21Mq9ds8CLbaP1AUtzwL+kUk
dXLjjeoawMI0J2VFvMURhUXWuQPzSW83uTInaA23fEG4cCoNI6SmrZ7PgrgiLJ3QaNiJgFZb8a7D
MArf8E3phBwhUo7HjltkrLQk8MT8ODAeRazh+vtA4wIMDD1hBwF1kmiKCdlD2Rgd6eQVo+rubwEf
41RBhK1ceqLFdoqkp+jzqtbI7UeGkI+sOLeoHz6gSGTTj01mP7uny0rCr7rMKM11kFNM+NDbHpmQ
aRVpV72mWrur4aYNa7gjtKowHX4P4FHtTXBDPKiCNM8u4oMZOzJe+XEp7U3D/fO5qEW5GSaWjVMV
BhVgR2FYA/y0y5OVK2y+82tL2x4ix3jt/zUe4s6DOZcJt0rv+EFRnNKL8Ta3NY6L3Ys/rg9wL4in
L83S/Bqhs3ZWqIXS3bRrrmVRaAafqWMOAuKjVTb+4nssfyCSXIwYYuhnDN1lzi9mz3T8R9VEuZyS
hKshCwfoF1f78Bt7XpI9SZ92du3JVIttzrI6zmXHK/GX6n0dvCfzTJHWvwf5t6726CK87q79+aV+
+4ExgxLBV39xu4pN23USFT6OVrzGb/giDztJ5jEr1EYpJIQTkZj0fUeP23lps+hqRVwY9acQ88SZ
T6uY2zs87zMP7fm/qiFIDKn6Hfi5ML/Y9vdiQk4culC3HF2Qnj1i45dRwpZeu6g9w/dCgKhoIXJ5
EmuVIqe/i6aWP0L/5kuff0GNBKA4+SSUPW7ugT4ijfN38ckv3PSauZ4lCS/gf9dryZHNU7bED6nu
1JV/bs5f54xI8RRKUpzXmWDNUUBlMcJ1jEKEuJ7b5Nif7c7FC6Jh3Pl5CmIrGlrwca3yytKcbBfz
Qr8U4jCZeRyPzQX7WRqIxrJViNRvnyUrrvIuHeaV0JgpPWsb+U9wc+0uBtM4M4/rHcf/Z08oytsq
Kk4wTGGo6V9M35/Qrbg8IzoTrjQ4uHsttSYZn65gsjBKTSnUZHCH/8v9VKGK6wsrMhoXVd/HTVVN
YVL/YRYrGw9ULKPoPJeMT2u7vkDGPinFqh21l/o0P6RhfHHbgCDL34nRq7epX32swYRZiu9W9dKE
qaCi44KMcilb6eANCF3kI1SvNlqn7pRP1uGXCJuaYXiZpkkNVl0gyoTkFTUNelrIQRTESddnkLVq
lvyEQFLUEuc/u4SJlzM29Yo7BQw3R4BmzIyV/ouKB5pxreUByvlz7e31K1AsCLaz5QN2ehBNg+72
gmJcSe869+3nA/wTd4xARIk3pK6fpnKeaUCdaUlWfKTliJ9SI4bpE/6QNz0A5NXxaZDGIoIkJwxT
P5UNOzWhevGxHAQNYefoUJFHDEVPahdDil8WbUWMOcs/pq47JPO/5AU5jSrXpkFtzOxKyjtU+NEN
VmnUGd9bEobvRZu02JM8O1rVvXY1eGifS1O1Uxso67rRrwNT3Ode2ueEE/OZVv65eT8Q0bZNlg7p
sJbdCFxBPyVAwpDIoHzLsTGuX056Mbe9h3DfN+y6BTrRht/88pgFCfJwy+JNBQQLPKF6j1cS06z8
QeGPvaB5nio9thubOsfynsXt5QThKN2+xOl5D1/RWItNniBXP7GbvgWBWMky9aLnJUqm3kqchBOS
lG2PuxR/r2Y6qF2lIeWKEkYW6zDiW9g8w69uPIBiCcAvo5tbmG2197IAnB7bBcwF0ad/x+A4NeS9
2NNoHHt64RrWndlzhk6yOOKswgJ1bBbgpKYdapTIQbfVh5jRCICqSDT8ypt1FcFQSXSgnQ8dSZvL
5YaP8GNPwaXEK+FErc/eLvQQUEyRe3GUO2WHQTowIbnjJpOwbfv4dVCkHyi1XNlqLdBwR/bABwKS
bYcKaX6tYVzwLXoJWgW/fsKX2iPqAlLvGlTYso8HbLqTyP9Jj968Vfi3frCWx2ZxIYaVckm4MPpf
xFajg40bNMHs4wU5Jd8Sl5MwEabH8q980uqcfTepmEtTLdKOWfm8SzzhBKWDq+MS07poC1plli60
a3G7YKUzP6da/UNlF9gNNr03ZU6C3vRG3t67VI8FdDndyxRX2qbkgfi726p1ShJrBKFLIIT2hMSp
T9fFIoE8YGVJKhvxfOO9dDuSr5pdRIX9maRhrNnhEEjW23DhA8v3+gKG16XfUZ4KckByeWuIeTU4
l4strzvkv3JevOPW9O8n63YjRtTHa6vIOdmuGDyWVwXWZ1qHpJLpZxuZLS5wm5uj439sFiEJ6bsC
MdWuJn9RDWzBcKVuJqjwu5Dpl90tlfWKUOkl2K7qoLhvfuBki24+fScBSMy7fh4DR1cXejLtIytE
nAsiC7TCnAHgxTwrECMFDRe+iu0ODdNYzaM5my3FHAt+fWv7XSNDRy85pHUMl52sMZObA4kMbf/J
mfIk+qnONVhiUrrIn451AdZWN0TIRdjxtqAdfvK0Hg9Gq+6oMAHIoKc0ZVqYWbuno35nmgpiFDz9
YamqSLZHPsfl9SVEkKMzkBUgFpS32fgsjZZf7JD35xX+Pk89/R2Yg1t9WCbZPSwKnIZGWdrywHnN
ZDOeJtSB+9dNq9XuXtS3+HdOcQxVbO/ThVK1bc5e+HwD24ObN9T1332DX1OGSiC+uQEJUj/o+D4/
FNHjNZn4976apN7+hW0SITonoZIiwSUPjMBx7ZvEv027HI7AvWkNxBFktz/QgCoNqmtoPNIt0Zlj
p8AavZOTByPZqgstMBL8CdnxtRRnWChXjNazROaaNF0A89qVne0FYoV254WcAt24AQwlFZku0gwC
v9GodILJ4r6Mh2u/3Mi3w3Xh6asCwgI/xzQ39lVFmq3vCB5yci25KHH518qfHYoZ0OPtggOZ8gfV
CDQRS5zGpLLIZ8rZM+I+ixgzQcf2GmG0B77r4P4/ZtdIBWqUw0tPXzXm+i+goTNO0lcWeaxf21h+
cq3rAL0IHlWIHkFIIMIek4WgNf4wwXF7XOPYv7Q5O7YXYdjpT3GLbQn52xWF8B/xrhuQfPj1tv4g
ZKnxVUry6/qYV+lHUdxbi7SoEBaP1ozyLWMYqMPgJm7N0hBXIyKwYtq+E1B3hUbkNmovQtr9uIMd
l+a2GgdsgGAb0ROx1JowiU5+jNI1jNql8G6O5nY7q5s8jJ/xjALcCwSiC7uOnS5UM0sqfnozojnd
hHEmZB6oa1s/2c/915YVkQi11gqbXurDkZn13wbHhbQ0Z1mx5oHrLAk68t8oHpVrtHOlou0/1Rol
HzUEfW//L2j0yCUl/H6ELlKn/s6jlJoVHwzpOkPeGcIj+Yyk2UaoanyJeIpB/1lW9YpldxCkcvHP
jMXuVZhdP7CylU/xLSutJWmLpmBQ7uUwcbK6UygdMy0d1gppKMoxJMCTD+yBreTcidWpvH6cRRvf
SBbj8fzS3wJM3g98mQUmP/NQSdh47ndm9L7PNO8gnoc8dSRA1ljSHkHrrhJE8nuB+4B4cx1rtihr
TqIcWrT8dLo9g5vZjCkEEGDgJdVcSd7sDpvy4UuK19JNLY4DhmYzvBZ5fqyMkNyA1JhCRV196dqU
BblWcrGUop4LfdiznYYh8103xQk7xdS+CpdPdkmsMPu1LYy9Zefot3/zmcVLBOAbBGq0B+pcuxn8
J9qhqKPGS/8w1PdJJ8nLenx3XW0jOyuAOLv1eEflC+Yn9hf/tsIF+3AxIngN1XdBsustrBOW0ZNH
UEgF5g6NSVBuFLnV4LOwVz1Jpd/wvYhIwJiwUVGFC8pFsAjy1YHTRX/r4gRWcJSRxpoWl2UqAgC6
0AE/xpmB1g/Xj7KKlEGGdOB5h4ytXqtPUTeSH0iVs0Ci+abVotTXkymGYYYk0r/3HhryFbPsQ9zy
etk99i8Zu84gUU1lJsCNCTRoqjgCGmMUa3d5M67GfCEZLW8cYgyrHeDSjzAHKY2llkpsm0bI+j0q
2cMBusLIW8ue0EYZJedezZpl3qmjJ8tbMELLeunOWNf96VNVcZLP0JqSiTnaHB3VcDiG75NzPnzu
CPgc9NuGOzLFWg69kfuDk2bEz0KSFHK/E0/vHIpzTTdottHtjlISDxznPQ8Zg/Idcbk3lwIWbME0
Pis/Oy1AtuzAA867DyxWMsHGhEIOo8AhmrjArS4pZPSmLYQcy08OIAxQoPxXJQorOsxjYF4LigxH
DWV3TJhQGXJGRKo744kZFKL2ZikherMFI9odJbc0TjngXtFot02UsBNGkUwfNqJiIXqJpYm+xKJ7
BJHbncYAmHh4jZRMKk0rHZqNSQ+RfASgQ4yA4k62pYjDpjw148lUGKmNAJf+gwf+wDeEaWr/mh7+
7OSUkKaTcXD8iuOLJkkmWuDOnA2aSBQF9Pu3EZgt5V9cBaVw8NBKOQYeto2XvEhZTC+G0ZQss5GV
Plglj40L8vqzjAQ1Ovki9jfszjDg7AJw8eL3NZwgbCK0KWu9F3n07Vf9G2boiZtahVMoeB+NWJaK
+Rk/yQKBuU/noE5h1r9UEvc9ro1axe3Ecz6eol3Khfh6OfSdl3PRUyDPT0z/Tl59bhwymgiDthtz
ihdVf6KOUis/3HOOXgHRsnrINgOT4cqRr38ggJcRYSKR/1Gj1Jns2VMnX7gudFv3NO/QxfTeS685
dhwbWpuWwAk5ZrtNqekzkkl2BU/E0oPKJy5TZOuJt+n6YwQUzAKbTMJem6xf53rS+CdsV2tDR+UF
PnRTtZyBAD/ixwJ/y/r4QN7oB40GzlY65OGBGRVJXT4XLfbx3aCwMXb4Tk9pDslICgeC8xwDPN+e
ht0IHEp1WOjxdzkCCbZmGGblY0ihg9CAIvYJx72xygmfq7cse157WrirJV/IzGbxACrHmsOa03MJ
UH2TqKGMjq3NV715R/oCyh1lirnx3NeLkVwlY9FICAFIyxZkfN2FebvuwGuAOF3Lakgwx0T0afr6
OTKZ+M/KzB3cUMPDGmQ210w9mtizxJlYXsMpxmASWhyEYKFNevQnrekh0UVy/QZS585fA+ot5F83
EeDQf2dt1gVReOs36tZigJap+WyLwnAYzV8EQCyLJi6BYaGhtIpwGwdLHmFcG7I7Pw/rO7YuUuk+
Y4MMgvx1F/5ADjJ61IjiVUPP7QRb7doHH0+Egqn3Ymq7qMVcxOnEWxnmVE2WxKPbPQVcNZWROAin
S3WCV2TgErv75qMyAsNVj6G2mjNXu7Fx8OGnqThg6sUkyYNhup6geY9wDUzSlv17Psfs0bTQt0Xk
J6h0Kc6iC8oIklke7uWVX20nqyF5EWfQkp6Y7V0M2+jREtrtQOsf7F2x9vsAmxvEzuv0C2Eg1SEK
YN0MEKexiOqJqREI5sc5x+h+ZoW+NMrg/V430c8NaNYvwoLRTjOoxh2IdCUS/krXm7r04XXfl4n2
pQQvoK6dBriV08btZXTk7uXxAr+EUL/Re+8LWYwzDERKH3oko7Ip8x0lrUHGyjdZL5EsxX3sHCtQ
MAhHzP/zxgm+TenO5+idp/u9UOJ9wHTCJhXNSGtEFMpH6ZZEOISooz5DgHAFEbneKmbNAANcYhZa
d9H/yPpcm20WFjDKlrex9+kRSVgZ7rC+H0Ix2Rgcn7QJ47RjAYbQJnfuvGQ8BU3KYC03o+Nyk/oR
RuE+bhcy+b/+ioWZZ8xgayRcRAAOqGUFhVxyMOcXMd4C54SLazs55djpHL5MVEkpPOQ9TvR1fCXn
TVT34oevlbXFDMvUTQD6PVcY5mTCxow0jsiN7olN3Bcws44pGVA+NzkjGzK7r/czc8ellsMmZj8P
zcdv1oUKbMrxurjpYGbltQ75duhYoKI+yY5RmtI2KaA9s7eCoRkMoyXPdYFUSuTluwlFPef/YygZ
7jhCNPLn84oLUh1EbIv6lzrURb4FGMSq2ryOnlvzjsVQqzSeH7i868wZHB+ONCO5XlrLG/cAbJkh
K3OPrrNCzt/0G0aW8OOIv/E713j0Q/FwKVzWPNPu1qASl5boLJjFhztLDGT0QQcWEb4us1+9MOe+
E8j++2fYO1T1qpkvhVz0sfg1rghVScX0jDMk0WtJ8YiHeLZL6bygJ56SNi7RHh7znEm2iIbced9q
ZguOBxzcXHrwpKU5SnV1glxLEfYAoZhlwme5Fc/SrI7FEIhWAq5ppjPHmLZjxx+ScPnr5HuIkYKI
ipiMwGhyJsOrm4bSj4IdNzTL3zE7klh4Ms2Sd5E8aIbDc9uZoWpHsTLMil90kRGdbq2WrW0Du+BK
5uYPQSKArn0/qOOe0kLf0c4Z03Y/nnZeO0glHAcUhJqMMhdyBjHbMEyLfZqVAK+WUshkkp+L3gyw
IncRNrqr+duqENfoVANs5uiKgCwo3vaoBtRnjHlABtgQW/8Wm7LrTBWgvB+vSazoj6rpzQ8IcDEL
hZ8r1fdp1/iIJfQ+I3N1+3OZji4kcxxA0C5KXlElXCMzkpoJbrOrdJWFqT0sAyHr135Ej0wwwJ4x
vohMMZcvHBPDzzH4I2Aq7JTKzefIWR72jizXPZUDcum7iN7GHn64PS8dq9rboX+uneHDMCaHg9gT
SUB15F/ernUzqxU2cFBat1uY6F4e0LZ+cfIojSc4wmPMSbU0rpmC7/+sdQ4AUL8Oy3m39u/P8vw0
U0XHCWPXeY0fKp5JElOprPyjJUR1NYXo7E6aMUvv3QeEUJxpXkDvudd67Lih1+V9g3TT5TUZw2+n
ND8hEbHsc1wOafcFR5SjaSZNnGUBf1YnaO9YlsDmNvMr7S91U9ggarjk2/mn18db+3ZFpoy/3sw/
un3vdCAbw/e9xs3L9am+NEdybSThJO+X1qiv8OoAWEYRklJl5O3MiCw4LhFfkQvcNWM6HXDhfNMU
1d1/BH9R8hBjixcTAtKgLzI+gLsnMsgl7Xzg98oW3pIkDO+MBwX29zWKgTk/PDLWOnoW8ipscIcW
bB7HD4dZlzB4P57njvPv7/Tlc1gngWcmOj4sQjGV4VIVnVfNKWfm61mKaNHGb90yYdAiVcDfw80I
vs+DFlnnVaoj16z+PF6O90srl7j2ruqTrnp9D+cpYtBHTTXnFsS7et2ygVkeI/sFHFGK23Fph/M5
X5NsYl2CpQq5Q/DY6XVRK0QAULQLWcdP3bqewtoVUd1IbGREs6lsA/IDhhuWN1HY38P980aAR2aW
D3iJRI/umTm1RfChKpQLFNx4yjPuNn+0u57VZY2C3QdhPz5+OzJgqimrevecubV4JDNGOrOuRXFu
qJVTrZLEPyDScs2cgZC0rQX90N0qf9NY5fC645DNaN9+R/XnpG+ra4ySh+jxnh5h4u6VYuEz1vL5
80pHwRRBZJ0nxc5H5csIEy3gGUqngGsXXd6DE7VKf0gu303PoTWfQieTsZ6WWHpxrK2vbf/PvDzn
0vJLJjY8RPMv0W8uomSYIr45LSEzponaR5B4welGWJj5xoDV4R53jKG5hQrovHvs2jd70WoM9a0d
f/4US/CzviJeJj/S161RajmyX8osLsMcR7uMahWEIhQz/gEsF+PnjeO3l/cV4Ms8fxBDJ+8HEzeu
Dtr4CxEF+CEth+KE8T1SW/INf9m5B0HOoynPiyDf6+PyHfiZUoLzXSs6BdsSSpwev4rbrHn4kfQn
W2XaTVtvQp+LYnpYJA4e9omQCoUC2z4x1sqMD9Wa6lLclNCJHnNtE1J6KZ8VjwAxYrS1vUX9PWLt
lqYcDJu33KuaRnnU/kqCFm3JmKqUb7cE/StA/cPQ7JkGVxaFpURnHKGMd81GqqnnUHtLeH/kkd6S
MNxhnje5wn+qLwTgZJqERbyL2QANJ07AxcMgtkm1C5ohy0kb4DhhN7neUCOc3HSccX3v36BHtoFw
14IXkP1JZv6SMj8X7o2Dh9co9OuopAvYlt6tF6UUuWFYBnSiJjq8CM7QCcSSe2bAaD5lxqUIupyi
K/Uh1cPD0CcA5n50iCgRvROjYrPNsDNNr0q2IJuzllBe0DPqEuI3Wichjw5k4JHr9P3oWgUBDS+4
ocqLfsydvMrze99ZAwBVGoKZFS6DM8qyX5XSSU281fYlCDsJ2daGbWANYODZyeRIQ6jk3ZFgr7xL
FQYX+qIdNjk6GVpKmm2RmqO85xqgw84xRU+m9b6PzYn5sz32LoVvtE+4MSA18sWjTdddNaM7Ju9+
AH9gnX6p0wOdqOvdTRnlfcvkF0XBfqfFNbyQwjIudTiLDCH5jxMU+FZQPahIPd2FGxKLbjdRByAC
fM7Qknbn1v0qYJt5nm8avwuN+WwuvhYbu4eaTXxTf9LyRZJA6s4YeMTKVkpEvmdSTxi4YvOZTgT0
tjYIZMfC+hmXlVkaBSFYbmmQparL1KRatnTNU/HPEy4i5h0VNKSZWAAaWY6H+wkewY/leNFAfU9D
SlPCsuoPvDK30mDkts75/8UhmcPmJaslAU9bDpEnCy6GiNm40PANA/Dq6eRazuOY9d3dnMA/7YLo
zdqE6nZ46P1lutInFc3G6unr1JrmFrSycNrqmWwST3rouDr7Osiz3JfZeeqJpBe6A78UryTgC2zT
I3iCBBO7AeKHs5FSH+Yf4tHY20eHxkOG4XhdjinQy4Zgq8niLgMI4Jlxekz60llF9Ju3p1hg/c6Q
iSEx6y/r9eKobvasY4RU4BAsS9aqhFJxA12Wth0L+2jP1sU8t3jvGTFjVGwyzzutqLSvck/V/dGz
oDElH59UqqQZkvh5aG0qo1h5PQcxrdP1z4zRMhbFnqUqmB4JUbiCVeyLxja47mxjJ/3JmpgV7kfo
4OJon1Z0NvsQ4W9mSUFGG9sZ0utG+qGUxt3745B0s4RjKjAhnev5uD3/w7ri+f3iJM5ZXPBBDiKI
yRlcMibMN1846j7ymy10D7ZkGvhD9+FQqldL6tQgZjNjMfJlHta6LnLlYurX2hwYjxxOqQU2yKJB
1VxjcCvzV5JGA8Lb8nCePnPTUCli1bLlLrxCsUJepXfSV/ucMQVQMas452fHw13pziUd4oWmVrNm
IcGBK7wBAI+1+zAJONN2iwpOK7VUn95Ne80u4QhQcQQvy4tf08ZzJM+00ltOemFJ4gc3kRH18v9y
Sci2gV27DZQAgowBOW+Ls8ZlszCMUoybu36bYGUd6zuKAhw2IQ5mYHcCCfEZGs7iqFiRQ4A5ixun
Pe4CNOHbFpREMuKVeKC+InGz2H9l+A49G8ZYixCsLTOJQbSN6h7vFvz3O3q90Yztw+QomZ12Fsqm
XrDeuz+v87zLoiOFCRV9VzNFF1NLSPNOCbS4GxADquzLlwY8xsIxsBqj5CS5EzHOyC87WZzu5zvj
CjiL8RHNNcCGWxlstVFO81933SYub4rZE3xQsMMoViZccr4slJz7u3cHOcOKGfWeGfQZAtHt6ZB5
KaSZR/xc86UmlbpVYNIYy5P7u8I8S3wwbCF2+LNjo5uYAmTz9miA9jXPRgv9WhNUIg+r/r6rmogw
z3LTq4M+c3EULMoE7RCnlLXaaeuY69Lp/dQ8YSM9rhXBIanGRi4XuRtYL+uItuQmMyhCMncPPAw4
8n7r0dx2dDNbkQl/LS4BDEg6VkP9I3BjfM0JXHb5rfxLDUsyIkpmjakkX4Krx+eEy1PZhwo+K5rW
p1/rXNESnI7iIB+H+ifIU9ZqIaleg8hpa7RLo866qWjGARqitgpcvht4hyxvlMN+r97gKWrBX5MO
QdJ/hmt0L1K98YHD/DeqN8mrYODr6zhH85Pw1SvREP7mVEW4XI6HbfkdxyiRY0CEsJjGSfGEiIxd
Olk3ps/7K+pMi5fD9eBMVBxng0+t7rwdUcfc4fyPVslu9SU/yhY912e2KsKHXSGcXkpBSWz8VInr
FK8hJU3vaD7B3r2PDcCHxTVPUL6615iFT/oRuJoIrfzbxubJr6sl9NqGVJMAAfmRM9NdEjStNt7h
R1E8ZFzwu1HjQnIiiEOjR7hgLA6aUXbsX9lPqHTMv809BXzQgz1+b2Rl4nW+sg2DcGJTrBeYbRzq
tXhYp/tP8w4zhnzFhYAQ2JBRmZNfrqd7/P0iHbjux1fMywdnf7z9W9zl6ERwOY9WTYzTi2DmWJ8u
4OaU2Cef/k65aCjt5uyN7FHR5mjSY7R2UdZyiS7sUVXqi1eC30z9QbRIUboAU4AdbBzHIQW8tfMv
ANV0pWhafIxMORVTG1PLDO3g/6thAILv/fHEuurR3TKLs37PbHO/GCPe97OIhYgXxTsBy/7KZ1b/
7tUx0xOQgXgBiZthtiuWIju0b1zShyz3cZS1i0OFAXGIPyHPl4BANpJhfjRibVfLsNXR+m2b9mSC
7I7dFH7gXcRbFwIxHpYa69JWBAeY/UIeKFENWtvRiAlK0SV6elMvPzRPsLunNrGAHnst0c4TOoTY
77whBuqJk/wLDPVGgCtPX6e24ereRKDMAU4h7izs3BOyck3LInlnDkPlQ+PmkxZuZJtWV2E+N/aZ
tH8j3c4hMuplH1RV12LobXSTiRRx+CNyiX4X8ZUDBi8YGTxpMxj6tZncXYRInHaYgOT9GWrYVELg
1YTH7GI8Z6Os/+eAZVuvi598vi7QTQN0V8ezQ/c2mRMU1mZfjRHJmH0CfEhSEwrgZvxLH6lRR0Lu
TurjOPJ6UxPqtuMxw4N0I4wvHIErenC9npGaQp9hZiGV7zYKCsorhhlISHPp+pqbEa0XQtsJpOAm
F59Ca+NrANe/UhSFRurMH8ga4qoevt5jq3cT3HZbGXgFwRNrnjHz8M5MvEHX9RL+P9tLKd613B3t
5Cc6jhqx3xo63yO2HXd3VkftPGomJ8R5/IA1Chb119F8BAQdsM/5bFmWrLP8pLiQ86vtCx3MHTTA
rC4vccmcX18liZVt0KbakXKKa6RotHBfV2DdhA/a5QceIdR41h8p3zhePF7qa4VY1t5W+hv+DhST
oVjWpH20i6U2Fkgz8IeaCO+PERHSC+Ftn531JKvO45dcuk1JaAioKtSbQbX+zHNGczIjRHeqiEY4
7eIAdwUFKsO6DSqlOJTRfuacRIS/qoUSbduWfJTUzl1JJYnq/+ipxgXZT1KJDZdXXQtVsFEKXwWa
U4MbUFr62bm9yP/xbFB6g0KOFSuj4HVJeaZ8HjYUXjDTcM4s8xFGDl8WFkSk7hTOGVDNedDQa/Lz
vkFgNeEp6ceCXY0CCRK89WnJ5Vq3TxGo/BeWU0sDVRACwMq7XoE8JXeqqvyDkWyFiGsxj+6uPmuE
lTvCAfzgQ2uNMgQf8cxnOfGau1XKMQ2bM9YZjYxYEFTll6cBVEOabPR2RP2sL8rkCS3XdspSQAlh
PejyRlnoLijHu+vMe6W0obTgHM+sJXwq2iOLInNCEkDQmQrkdykJweW1joflI4zXSzQM88dULDGX
stT6hXlBipvT4DZGJ5vyINTkticFPv9Ig4sPJVyiQaKqnaJqZLzmJKT9jpA13eslFWeIQwBgDi94
55rp0AOGl8aW9ftqSpD+GEWh1dcYmJk6BDuvZ3CISUwOjubfuvlbthocaFJEXkEEW32wkQhdFKXy
btBlp1QvH6iYkG5jsNrwUW2JtoASfffnruWRB9kn1gAMCrWutKHY3X0fp7aF9sE0e7oam/JqjjZN
L/081KXxY8pAvwTQqIH8I5jT8BVBKQh03PE0b3eOJ5DoavsF1F8OglrMGZcFjsfZ4LZte0f0WTqR
FH7U9uZnG1yv2UYKRJ6VFpPu3EOYF0dKgDlFkOEtH+RS6jfnZYdiSK50tWfI3C4UxuLazPHw+iGl
o/IDG8Hqb3oVHjszzwDtOt23GQK4ChrllVJV3EgMV9HMMP4W333BPSmja/LqMyJqVx+cwUXFFaTb
dxECOw/XjP/KC6j0EwFU3P57IqHnHU/OQnmfItRi6nuJ3RJ6yEFx5yi9MXFzplQ8v/OREywW6NJH
hPerK8GaL9qEe0A3yVcbzkvhnGB5qwsfWAPT2DNOycfzZhza5mzi5lVPUyHoLmSIvxJCwIEaCi26
bgrySEPzucE5jdDWBvDqvGwUtF5sDDRcGke7cj9Pzvsy0Dv7jWtX+0WBJGfWhfQyIcIeBnKjp51T
8Q8K2ZEPpNubismrFXgU8KPBJ36w+/fw1gRjK5nObSZAMU4ajPCjSBZPM66EEshWsvNR28j7SIE5
l6BwrFAtAxfS6FH1j8nwQisP4wqaG3BZCv54ImCI0p0DsZQx2CDbgeedVbbVnPeScUqI6luyJCRX
18THT7gVkVnifVTipqX3khvT0Kf76kiiXP+WSXLj1nBQcOR+L7owgyjGxQx5qHx2vGPHJtKe32Nj
45A6kAoXKquLDQp9IVblkACJJ1KqLcfl7/Tb10eZhtgGKs9sPu6xT7BmECENmLPTsI6FcER6yK4/
OWSHqG7hyyWmYzHgSeYdo0cDHuNNtAoQ+ayy5gOM9dlM1/7yRojlXt0+IeyQeU1qXD4Rf3rdAmxq
SnS5N0X5jUq7z0kt7kD0hAF2bx1e1Vq5m12wpSnwQJOmXHk8Ik/BpsmRPBGR6GTmuxomEsr8r9o9
13v5dhOTBCdZKq+mMPu3Du5NvOS0URuLFCmnHoRwG1ULyJsEK3TR9SDmljKNcDoTyAVV6scdC1vb
Oxj0ZVMNLVTft7ysZ6V+iHaMhCjTyGYEYvJcYV6t1dln2kihHZyu3jri3GDwzmbDlngdhj0/N/6f
iRm4tmSqYonqeIs7z6LCUIFu44GlYxqXbUiOvAbXxXiLzj/cK8TauoAj5qx3Y/RBZYVmwx0abRbA
MBBFj+ZOfYu0+ypaipUw5BiXCUyhuiuuAWVMGM0RZnXu9c1Ia52/KwGYeAkjHJf837rqIEjzDUfm
sAD91S9uTT7K5LUVxQY3GLkvjmS09EE5BN75F3qjwjMp6mUoF5FNDC5qmw5/TQ4dZzxZ46tLFik6
psOzdsJCk4zXlTe84f7cFk7NkTdWEpTNO96RdKvylTS6ZVb/YvunT5tEAfsltlwsbmjX3tX0z/ru
m39qByQX091XhKyKanZC+YyZB5JXBKNEuyPsTcVJEMr5lDQ5b2ihVbjCNyQ6V/UTiaS+2Nsji4Nn
BndT+nZ79wWo1BmDWEF8Ut7C55QHlcLlV0lnJS4aoiEUfwvK2By0ireJ/8XWcm2pfXjTUPf5kYnn
eg6s4kiUDpiTSmiztjAhJoTx8bvXIlIEREMjSyXczBGtaKXw88MiAmfJ38r3buMkKR6nBqDAQ9/S
6Ws+Us+NLOF7JIavjyjzVO3ajNB8GDMbcxsuS+Sqb6TJxo6Q/FnofF5s6Fr98vgluU/mPZ4lAcU+
1OXgl1sR5cjPGX2L5VungMoYitTCqbTATSqFyUC3BPdXJcbJrtw0EAS9UIB3lNbQdEnDJ+zJMOR7
kHjslbMGXThjrO7mly7ej7d49t8N3Z/e1ryArO1UebRP+Pama9PsGlJmFPNSVMBZJTm4divBMAJk
BnjpcPPygTbRpG/QVArEb23/ptgUCAX7NT4ujlt6MyHPdl53UWrEbChdjtYyxeTH8x94JTbDxV0d
mpWZ/mJ17n+hrHxey4djRWK5dphATfS8Zo6/zOMwFB53ajru0bcdj2P8c2WfH6ZVuQrzWgZYC3zL
F3iv4T59kXECmGdOHVVg82xZTxf4N53uN451RIdy1+Y9CBP0u06wqVbarOFMf0c7/4n5w/oCM66N
bHzqAMq5dR1++VolYQISqcIGTe9raS0uoCZW+172+BJc4BUSlMdNfFWfCiNOZT6AlgWU7dqxw4hd
3KeDw74RVcCHtHXJG5oPMIAyC7GolZe0p1Ofaig3tIanR3mfmHEexfqIo1nfh/wP4+z1XCtXt++3
zBZQCme+0NiyH3UWt0t2z9N/Ee9Rkuo3895YU7Rx+X2T3WH5AFvRSy1W0W7NBDIdZaLyTt2paCwO
Hi7H41h9veAp3TB7RaNjhEFJNv/WmRtQwUpFkYHsIV74/WA26gAuEAIZdJlLHlyi6cqRG69jzMF6
JlC3tXx8xzh/SioXCmKxmyWMaSNN6nKqVNRSKzwc8Un1TBZNFwbyd4pmlAW/mfRPMuPf0+IKlM6A
GgZdlXPeTxwV1s5/t2u26WNDxbHkYLZp8hAflFXMGJSoOpHtp4N08mcEPXA1XC8E6AUkIVlf7QcK
kVgYqqgLBmE2g2yp1MdVU/6Bxin8tZ7oKO96mHT1NIUOYaYp4Dqo/AOm7X2+erzhBnZC2u03V5XC
puQyWZZ5BIYBYFNeooFROHjz8qVZkaeVfSpzwE4qCQ/j/aKW1z3JyeD4qRQyg+u5Q84g0jIJ7uD+
Q5Ab3nzFyQ18NZlmeWIaTLpf/fcKHFAnrUrWy7pnfmF3AsdpKh5ZkKMJEeXEvaGlsoiHFV1eYmZU
8YngPW2IKxGxDB8Fv2O5n0Sl3yth0eqXWBa9bgnxdjEhGqOHauZdTTDaCKMDICCW2Fvghxj1kvae
Vx2wo+DRuf0ijccjhxepswyWQ/MHMQPWqBgQcBl4/g2JbuCtZPL4E7kCGmp2S0tRsEgIfQm8ZYFQ
YrB9UJvHuLJ7VKUu49daJVZUsBCOViaE/jB+LYMaa21rK8dBxO2Wm3LYnbhmwwZ1UzsuAfTGnPs/
WDDhxlF0/SJy95YrdtZ0no2GdsHBNueISP/cu6fwGmyrzwqlUFaFw8aZUCE5cyqkNmNrt+9OdfWW
bcSvJs1bsHYxTBlIV/GsyaK7tFRjcH2f4ua+6Jy3DOmOnOB5+9jcdYadIZm+10VaeQT2katCFKMf
yvUV/JQKbFnoe0/Qw3wbfanQuNoGuXdAS+9y5+bD0PDXSfmESyA7KK5vNDf/cOLzlcawqWzsRvpf
CUguplJhxJXyQSdeI49/M4o+xzyvzjbNlEK5dNAUTg3UfSJMiQsN0UsDpYVTzQvZ8iLaWntk8HDZ
ZhYtQFy7NRoZqgz4xeLGIf/Vlvcg7al0E+hs9m9/r+39nLuHUxNGo9wOJ1OVMZzLNyON0j/azP+7
s52/z0pkgP96vXrGY5RdMMezziixAIDVdOrVu19diBreouFAcVFP2n675CYoMn58TwZPcdxZH33g
CxFeoZr9mwY4v7XXSzA3GRJS1eCGAyzzTlO0wrT190yaLjqCQkROb8XaWMIkS/30/IsGicWhDxu+
HyyusYeILiH1xC15PGnuOui7tcLvbLqn1ZBCukU1zXQ9W8kb1TTdqsol030VgHbGz62nVnOyrTKT
4UEh8eVE3q3piZuVwTUYK0rCTH+WqJa9qbXUVkv+Czvp5DeYXVaD9PhN4vZcVFtsZIvUpbHUgXSZ
SVz74HAICqu68Aj2r9nrLj2Trt0jc+D8RvGf9JxEuv8xxtuKf20R1k/fa8cnzqlrp1G2HfqKh424
VZy0Jmp+LX4IIemZ7+wjDBmLVP1LpemQE2nWtA0WC9tUea49h4llURElXdJOh6p5QX4m214377ww
0vQTFhC/fcI4w+HyyN1vm8zhrGn6kMHub2OPctCJM0UdIvPjpjsoKBnJCvZBZJGcdLurdVcwXI7K
exzLcYvaB+Jv1kBZW/13EO7F3P+T3FK9Rjdao0x+wE3QPNjxKjim3KX9py4L8aGM5c+W+EakpSw9
72qjXwhuGbrU1PQs1PVrZu7qbKf/j8++fIsI0g1tm4qW/taufrAJtxdtaC/v9bCkNW9YGRhc76Mw
XknOeUgE0LL2eP8fYGlxFBJ6sxugZzTxzmxgHgBzVqZeASbrKQsSyavALBBpfgA/FS06IKSYkqHC
+cp64qoq4W3SmFMfHV/Y8pajJCp69n73pr7msUNPpsqClezMfTBFHJyPWrzSMKu14uipgJhabpqr
d/G3Fq5S3J3FCBTQVCEuqAFinhrnlI18D665OfyzIi9CpyWWVOxYrp9ajR5U4NaabZ5sHHsmgxju
ytRo25ddsCbIwdAZ+tfFXoDNj+Z35Ei4Mf4EJ1MijS8LB+lG+Rg3QlLUF3OTJWvfJN23e7eF8RRb
qQ1sS8JP25HIjSPBa4lRUwJTGxMk+HA+ymcc2c03G2v0b/7++jO8kJYttf4venbulQkIYyJWyLLh
ZL3sGYPSC0bHEvf4pkRFDo5/N0IRz7cT2qWqf/YmMAE6PPboTacQlKynGve2TJuz5MEPSU6oP/HP
yzdJP/lMAZNF8LgEsIYaAOWKuNG0ZPc8T77BMrGlNIIIK+bgWQuYM/SfpXZVy96h0T61cYRju9rE
Wcm6JvbxfWBS0xPYepmK9Kj+SQDigMHrzyEapUziaKvU0JIptBSHagO0mXm+VO53BJvg6W/Tg+/7
O/UxngWztpy6eZK6Pq9nNBM9Pp2YFu6Rn2wnGXMvLUVm98vAuPp2FCY1eUHKOpNFDNkMMlRfZECT
hoH8K/4PSxFudme4uv14wZ8yw1gUiz0azZsJpop9o8Oee7yxYD9Ax/EsOy9fUxvB8mdcSuhBwOWk
NcZdqCZ41yGeLDIOJuWlggJXpHyYrwMOHSocrBLW4Ps9r+zAFUDzwN4e9guHpC82J1O9GHf8QtWQ
x5jXiHHDgeITmbRX3BAMQMinUkEIHyux4QJLhzeGmNwJaaJtMKkj1TJ6n/TOZJf9y4LtQzQcQ7GZ
SotmtidHvgOQ3F7IbaJdF1SrN3Ajg6kDtbfJ6IMmcXbEBSWR5h/LuRrWsq4MBOoUSAZ6Am9cVMJ/
1YvcIlDG4KnxS4Rc0D0rdOrF4pHpRjo73TNg/uJwcAPY/zCTNXCZEIhjpnw05YVDI2le8y/xYsV7
6P9ls4VMQ2mTroyWeKVE0LtllUrm48Zgvql4v48aJQnRJ08nscvViJdGRmFWsjJSipMS61yRnUHl
2dFRKfOox6zWy6mcE5sc9doFyfNXT/SC3PEiZgsExBnyJstij8R4PTOpuP1u8K0m0shxbH6LjSp1
vlQEyrgQbZnGY95cNTbjohSnE6GM991X+DgicFPnQ2rYw8rqTnzt9M+M/n/ml+E5R7NCxxD7/7cg
bKsCAuLpcSchTWSE/e/FY8MGaeF+xT3/Y8wSGfoN6HdDlMAyCss7J7YYGJFt/mpj60ob2fWiZGIv
yDD7J9XZmW+1h/GneAqFYyhkuATGQ0u212k+12NrkjCwI+wxpB97cVJzSFHcpfOXWZQcvDinEX0y
3eQinmmZRfX23H3sUY97WfSVMWPi6xfQvqLyyIvDsRUk8yKyNBdyQVSvfk8wQ/thyqPj9Ocmh0/L
MGKd8rvQOZT9N57+61dl3ibSQl1misDTSI8q2PdT3p8G5j4lFW8H6+sdzJ8TpRfWOsMe3GbjRqzL
ITqYm74yzL+DRndt2z9GMq/WFNaQpNu0b9GKxIom0qrFaFBRnt4ISInr7BoHeHEodi7kJdrHbAOq
8QWRdsaYihEz6Us/3/pbFYIUgMC3GUK9kF6N95GwaJJ/2VnlsHkUXPkXeOVwI+CROo/fOFraaAd+
0C55rV9d81t1hgUFdIFQ9ak+IPk/vltJcKhwJd1cL22vv7m3XfGFlmZiziCUfHgHL9js768bec+i
j5kvHda2ikXtG0ODaQiIQS7zcrAZYvOYzzcNP5A99nGiM2tIQOpJogiORvl7Ookya4ElSp9BOntF
4u63T9FvXyYSrb7I2Z86g/a7X4Lfs6pW+w1xPALZusGmjvMURkpLhXxWfjEyRY46q+DbkYqlFTID
qZhemBG4c1r1N9vYvwiU0B+m7Vq3kXnUr3nvj3xV56JQ5fdvu2suCyuM54aMVEf5rMZX5ABA0+lg
KpLZ7MmS2lDaMjsRAjwOiYpXGbxVyZvwhRxiJRgx/5Hc1ANTOXBGGhK6Rx9CTG3iv84ApJfxEhiF
ATrmxfYCvfVD3nw5PA9R8cAEAWSJzK09GUEx7nzOJUJWBZJIwmRnmWvzE2DAYEPf2762mdHkO3k/
fqoEJBn7RuLu1sxtQApeddcCY1Zefq5InArrcKGVr4gt4FkRt5jdRX8vus7Vg1JWmWt8S5RIPjum
uvd7eZ3VGRRHRifni5CizEw9/XdVdlRiowAXhmHBnBvpYe8lmZcvsgF0XpNkGpiZNdWOfWtlZnEZ
hRhcfNE8nIVRBA2U1eCGnaAbC4cGCMIqF0TdJtcL0mKeKhkBlmrGWy3yh3llG8vrc8YQ/UYFofJf
dL09DO9kusEHgdzcfNzq0TrH2dNK41mtAn3pdVR0f+VBYWpPgW3fyg/AukaVQDEjiCIbrZzBi+2+
mzJo3MUgcfte3u+f5UnySVlMDBJumXaOLj0+pvh6mFXa+P7irLGilTez2affka5Y0BW48ryAoq/S
nrShPKO3y6nFp4O8QnZhiuQ9Gqe7Tf//90H6G3YXtIh5UUCq0NwcoO2E2CFi4QmPN0MLFL/lb7Lu
CGwGBkIqNJTt3WbHYUWADaRs59ReVt8OBWpE9px5OMiEHG0iLjDZgAHAiJxlNjIv9imbjR12zfcw
TZfgrePRFwC+P5VDNlLYGf1zF+qVy9kUEm8eFi7Bw/M5riet6yGXI23hNLFbs2w0Lzypct5iKxzx
us1KNkvI8tgqjhy7Ld7m03wTaV07zFQ92hNh2JlQ4/jrAFbcCIh7y6YEicFoG6aCUH9GhdYbY4OE
cUQxGCizYHQCEZH/UyO4kD42zGCkv52L0oi/2EM86qjVHLivtaLMm+f+aecusjXmHJebKZXxRQDr
ZLh9NexcCpyL/U4btEFHWBMIjeuZFihgHa4xp+xwsPM8D8Qp74fD+zrSJ8Q4yuvgst8o3kGWJoX7
5E/O4qH1161hHydXGm2mBfQiSs/GmfcYA7XE3ijCjKIk9UjZr+3E08vkTph3tQUdu3oYoBlTPWao
9lfnWj0wV/BR7pxbocKA+LmV1o/jo6x1NB+Idl/xkqyNhnDc3bKfd9tW+L7Rb7NJJQzvDjz707CY
wLtWJFQ3AwTKBWYb1UewY9TOLGXcLoEL65Ny5o88aG/Qoai5ftPELH//6ZuANM7+kRceVyuvTkZj
aaYz0610aC6luenLHEEQmxVA2Bl8IIEbFhL9gG9tUjkt1jyCkyzS521/2B914u/CYnyJTwoqmIJv
/v0P3XC40mGhDX/w/jTp/35T1IByWoMRF5+VqP0zeWvJ4khsOzs+pdtz753/0krJ1cyIE4bKdzrU
OJQklJ8MOT89HWOXEQGPROn70czAb8NHzHV4hfHQBT7ZurR1fMsQAFXJ9RgdwERb86J66SNltAtz
SpKkxztVTlwajzu946VyRGyOqGSPildy7zgyONXWFuGV0qziRvPu1ScPfqXRoNNGWVQ5eE4m6YFP
c5OWvEAOx//PvEnVmeRM/zuVhxD6hAQD4Ii8iht6xfMS4smBeS343yQt/iLWWBPkRVSmQyhuepQc
bL18tATXPOdRHJTy+KI3U8u2NJ1dd0kfuw2FRNJiB6gKOkaS/Qbz6EcTVnBjqcByd88XbvIElaDa
ceywWhqWqq+x+5IskMvZUlJqxV0SawhDt/NlrGf0IDbk43EZzVE8hEG82j3IkXfnMtgrGD1Q9z8a
XiAN5f9qOQXwbrnGJ8djvq3odBav1QHMF34x4M7etOL1gca3TsDBvoq8TA0wNN7smyv6duRMZYM+
Cbp2wjTow3iu1o6nu699gUfu6pB+Pj/eJ3pCcEqADtKBtCx+4rrMr562GV2ZXv7fMs+4rxNSe62y
To5KL1CicVqACdSBoT8HIYbWe6C1FCDqGFKDeTu3atWgty31aCjq2MnI53ZTSsM5YZyvOGd83P39
nHAWo3wS/P+i5l4PK/En2SdpF2SwAc6b5OhAgxI47VU6vL/lMUrsJY/4BRjXdzTwhOUVxplYlbBi
QXxlih+VInaI7mExZzomjShzWoLA7yHjP0KQzuryISPHllGja2T639MKQMehCt6h40za9dZvyF5T
IbJjsVKE7AFKKutPEcTAhg/IOcCNWiuijoUKt5Rv/4I58csSfUJ6na9uUAS4nGU5mb1ZUZJkMASm
jiHsWTi6AkmBKUK4lxtf1SdLVjYw60Y6E3+QZUpYpY4qRwtA2jtSNY/lUCpMvuvd8Bg6Wi4cgT7i
RaGG+ib4qbhmVnpXJFqDAxuE9h99fHiDYvn2dMVEiH0sQ7j4XUllM/+BXolByhV/foSor5Z3+CTz
OCFva5uhlQt4HGXV4mMZIALWLhgHKliCowAvcKLXnXnVatzW8XXSnMu7zKk+ZKLMwdkOK/dZwqiW
Qz2y0XEKOBLlEc3SCa0/bnPZBXOW0R592ebd0+x5nISjUuAk5dos+gl3QQhb62AhEEFJnoR7t6he
bMJbsskQWmT9R/yQGWQsaT0NOKrv4pXYJ6ao29b1Zegl71gBUbnbMEglbU9gmVrfrcDalPAEcJop
OKy7hZIjcjd8O9PVONM3/NAEOaz1+HEEbB+CX6O0wDWs8LWKL48Zak5TRWl5AQPDcNnJCxTB+Tp1
u1psxjkTIPLijOZLUk0R1XiTPJ6n7EZjD01n6iSt8olriITAZPcPpH6qfYtNAZSj6+HzUEUX7IX3
7AV/DA09xlQo1vfVTnAXz5ax17Tm21ysAMDzgLvsZJWojuf+GPL8hZgFIIr4N83iBpOPPsgD1qHR
ueo4awFWNS31F0LgK1PIELU831qaGU3ImHrVKet0+J1WJXQpBxUjrSxf46N9zNG2WBTZDC3/DbCB
xl7EHU0Mdkgn8be9QqyJOkuOKpVbBJMX/5vscvEhtsNzchTT+NOb5ppoR9VU7eHMN4fMdMVibo27
fj3Q+Hogp+zu0rk0eAHwJ3w66TLOzIeaVIzFqoreTpxLNv4UBaar2Hxqsf4gV5gX49RBX94jg927
yqbiRgWOc18cFIYIu3Oez66PrCRvRFscOhIS2hTlktM+yLCxUY9Se7JP9HNmw20+Wj1/8WM1OqB6
wjT11Y3PIZztnW+rMjrDJ47FoYjNAnBsMa3eZ39Dss6idPWipEhPw6VHvn7NBkRG2z8MUu5lQFIi
1TigxzQjASUPywjVUGpv5m98KKDikZvEX3D37uuD6ss3PuPYuMApbckBfSltAc4FwLNcgKJCRhPn
5AxOAeBR77T6jzBxuujO0QyqhEQDs8fviv/JZKgW5lI7LsLWGDVbRPqVfcV+neN/DmMrwLYkit0t
6B33BCJoOZcuya3ML/vr8ZByd+a65C9dRcBdjGzJitxfpZFI3eezxkz/44iP0xxPznLCq84/PL/x
k2hKGyPmPk3koJ/bDRMAVryY13qFsZBHV5UNlFQCqNbT2GCUbnRym8y9UfkPMVLpWngeD6DlL5e7
DIfeVLMYHvL4gllDl1i8193B7KXh3Tfv8LK25sNyBmvHKMWq2kvWsGDYeUweDCIYhjTLf33c9pYL
Q2uBzbG7+w7hue0xjlY37M70G7wls7FkGaumwl38+BAY3lvdr5UFLmwcV+BVti/1/7jxXkDxsPh5
OxsCR6ySGoEHpVgBIPUApmzvykssrSBOifl0eSi5ZV8rBQ4nHeXz2i5qHW5lB8wy2pizO76NT/Jl
XNGoI6vw41LMj6EfKlPBteaLBiPBcvk3fcoL3RosH5H1BF8UBK537SiJ13dadSeDIxax7mHVO0zt
e/DW6+mWWKjsL/GX8H1Yc5cRoqPvnS29BozZwRA+Ps09CpoGvsF4Rp5hMv093rf/lbb39kUqnGXa
mYTTqh9UexF6lbgCwZfT3YsHBn8OV6SoLEvJerpRJTmCj4mT3bsGrloLXfdNjWm03F3YaMrIKAhx
CFzwELcydWGSX8360gQ6dhD83OniASK9egsGevxd2by+Gjv+MgizyTcVmYvutfhZAzHEoAADZNjG
tvw0B4yFgVfHwdlvaoMUEF6WWeHaKAKwl2ieEbDjv8BXKjvEmaTru9JiCbFuJHvnShtybn/vCRhB
WDr6Xq4rW2XUckyyLFebb1szT0hvVlr2tcaxNmJX74JNE5w4PZg9j4OljMVmX5O4mBRHytR8YMG3
q619gXxF2fjVDL9jSqCVqHy9AFxMnnbhGUuCvHM25lkau1m+btebiX+VsPzEpqSPoo0vNYtA6jbD
pe6fT44KXNwdtH3C4qSeStKquX041vVvAsUCs16d2GHmNCKqObEuV3pcTRrAK7AaoDgi2DHXz0Wg
y18FLPcdVnbu8BReyLjGyJwEdPtN2OHtqaZmQjbZ5WdzMzW7z+7p6fQJakXEmbg/ualKm775pEsz
jkpP/gSJ4GAR8dhFHTlylhrL87yst6eqb7eJJuwh7U7ktKzyZX9Qebr6Ct7LhPUXvgJmv+w8J0vt
937PJ0dFKBBqUzJlEkzbx8gMQh5dqN25hv6F3wGA7KlddckmZ5Q6JxEDODEQJlOPsC+H2oW2AWhQ
uzpVkci/wXlNy9zfvmsoX9ZR+QDFnOr8JvmHzNd7Xf3J9D7wGVM9YJ8VJmF82sCwF43JH3ZHzzzI
2WeQOZ3Itbv0zFpYaayUhTx2V6VxYCIyrOIR5rwPZbL6hgl18hX1ZfJcRevPf9wFwyxJhkuMYfoO
8hIxXj1bCwMD29dVb/bGIQPkU+NITUD6wf+m8FnhtjtXGJIKxV5aa39FK5XTEGTymnJbPDWU2xIK
7Fcis3ci9PSXApq0oExMzVqOZRJklLGdK7Uj2OZo/Ku9fWWOVLh5iLzWId49XlqU4DMRlwfHDH1s
FTVtWtNwV7AmaBsQ1izYaRQvkUGG87H4gZEC+DArGd2a82mr4RUB/tO9xKcyA3nuvaC5QAiZjCCX
Me6d4dqXs4refvr4dMbri2OwaK7tb9yS38W6XLCTkL5dpgQ+S/IyjVRIa4z2T0Bf6QSgYyvKQUjl
9YOLj/04CNXwbM6fYbm3/s0I/+CqNeVyR50uhmjwrNHzFum+3XyjU9/V4jUGHaxTZwBljNuYWkuG
mec/ApYEYOdHmsb0cA8IjaopcZdlLvv2SzoNtyV9d3VANaosaPv//AARNMWCYSLsKSB1NrihLoJg
oP00PQfgc+4DMbitmdZi0rWaHJrD1lH6B2qfXZuwUR7JwdbUu2/SyxDrgMEHKWyUp8XUliQnSw57
9yRXXdAxDrzg1A3OzmIAhMa1JMZa/PkRPyA5/YNi+IAWFj8u24U0SfGegZxdtR4L17zihsQW7m28
hoysEhlle/jrcx8xI1VQe0KTaTXjKddhGzQn9KZbSsPUj5UlIlhg7ssMDgBktPrfnPP+C9+tMUoQ
rKACS9x6u1/TgWiehbIBKDAYRdnMs6wg36/TsaJ8aMIhpfiSBDpbrdGkpaWdrRf3OOZ/c73+9vww
Iot/UxLxj3YqOgWVvAqrpkgGu/btn7Olit5I0PzDTfAcnrHspPrtqn32WQE20fC5O6mxPJ/iwroD
FVNFXXkrM65B9OR2nZlBbVBpVG1C3DVbQ4XSlOT3dRYQlnuuqH9XW8ppHFZdS/NLYiDMuL44GSIG
++BJgDOhh0FIKaPirzUhG+jvfUmqsLjlva3OMEOk80+ASQ7DLjiGrupD2GIZQDwJgHHTyxz+1Tcv
pZcnWGhOQnpvfnk4oBN6kABg2bs/++Lf0FiMC9oe0+itg5TfHuoCey9Pqz2aMqi66e0+qe1r+b0X
J+SSaPUzUoAds+T6fgnZb6jvuYJP+kRUzbgLFaJXmMbAplzOs9Zz1xINELx68QFuQCIHJdQsKjlr
zFo6wq7xqLUa8x87lQYE8KtZlqu+zCL0MgkGSrJ2KTi2qMBfnBDmhH3mlA8p30VW16oiD56tli5J
Q1sjTrRFSCewKya30YPvEfX/8cM80jF3stgBJejeNWxnbCM1NDYDqmtEQVyjqzcM3IkgRSJTSX/+
IRFe2rqNHNEkSThNGzSrvjXvDuqbLQ9UdwqRfnYNUGutHnUtTXT3J2LlHPvm2POqHzbI5cCTLmxM
hTqVk8RVHIItlAojvEKAoL/e0PE97FTGyrwrktFzqX9D5jkW8aelk0Fy2X5AUdqR10VyFu5BYkyl
KlBpUx+UIdETMMdF1tVgL1YRwjWbgFIceCi59q0341WzgHNKkLWafmxbMBkYblKoBOcF0ssIdpYI
0DIshwKv4aPWWxy7itScLS8WVtW8654MLoRCgdLxQ8qSTZ7icDqBRPGONjDPwAkwfEEYNP2LvWJm
Ll0EI8wOQu4qQ1di3tM8E5wQFriTgzfYSgdr5BpbKEDMKN6PzpT7c2OEA743D4art6CprqK1PsF3
zTrdj1U+0eavGPQOHydr8yYiosEKS5LuKfcuLyPOePNdQsqBboRz0iLohtW/acrKZ6vnSbFLD9K6
y3yYHpwQ0TsU2CTPhIZOPyquAKSZ0K3PaqdCv9zHR5fxKbWKfB99cVtaAIt42K51HRnnnKE0p4pd
7HNeHgIs4JpvNPTTFy9GjGO31bqlbxQcrEoxWD3ZmzAHbtJZCaahnigwlNb9GjfmBsadNCLk4ajR
gN/nbtv/g0NKuEueAp84iRL2B+0Mq3t8/fDa2iqL1UH+hLOL0Kl/YA6Zp5m3o0AIdjDapfry+gYB
QXHaEDOsoce+YNHmtfOVcgnpbO96CXY1cOR2Z1Q/7uwh5qPZAhoBxNY3WTE4/ZL3gcyAt/t7ykKj
pmERexWv/6zF1+KDpxsD3KxylpdssdF7467ctjTcA611efscB6A9Wlk0zG6qm30CYX/sWk3PFi3s
oAL1WALrr9K1yN0edx5dUxhATrcUTqg1eLP32B3xo8iFN7DEMzVKRjWnHNF+Xd5tUY5da6OZHXgG
1aRxnxxWidP/2M14dvonrYvXWXGPfl6FzLpwHAPTO9SO/zJ5bw12ok2T4sDdSIbnBZr5ztjengTO
l9hqQ161VzS2IChatUdxsD2dz8Ho34qysc86hBylN5OCUCwglGUuVrcJHtwF/9b7TifS92vHSTHz
jAArY0DCz8gLBhmxTSrmgT9LB54sYtJa0DqELZdBmIe5r1du5pnw+Iiu99BSfLWfYT+PXAcI3zDh
1oigFLdcKWQPaih+2GNXRrxyvEIH4Aj55gDKUQb30e0SrHKN0f/5ESJnl+lJt6Ol+xC5ubX7Tx3e
oS5aAXf+G2rOmjguH9idh75ffBG3FEUvI/1ZMF6Fw4N5hAmhZZx7HCec2CC7CnktSjJWkcbeoVkr
qJNuxJz13WROrYTwaRNtTVWYbg4+p4vGo6NtXpwyHCqB63sUFICJsf0kHWsuzBq95f025ojGzit8
h8Uksx8C/QEgsLSsMwAzyjWHewvmRy4w93vKC2XwGa0k5EMvSi8P7aWmtfSTCx8ZGBD169kvHzPC
1Z5mBWoVnpCOrpNmvMIc2EoJpzFE+hMDHWJv9LE5xOt+QfVxTpmjGku/VRIyLe0YfHpL7GwtKGTD
5OwquGKP2CwESIMAi/flfdE+/nKRAeuC2U4zc9dfEKvkZS+gLP2yiH+ANFjZIhXGsbiMztHGNVFw
Fp0LVTKmvYfk2Uh7pPWmWKvfk6RwLUPZtE8XaoI7meo2+xhfS8y2M5cCXNzxnlzK0XrIBnMf6f7m
h7B5PdbnjCB9lRF+Z1KYQsFsjUFhY81V3xh5kNxGzDUJyNLu5iy8vbHMh6z2U+dTZotVFQT47kOR
GIL7R1gwySVlhsQiwAfeqKjG8UciZuUpmBYj4DQjyhC4FwFgYZeNhiQlKY5ZfAw4j6uyJLzGZqOd
9nilSB10I3wSEUpH2FVHbJZNiBsTHA7vCrluXFeIGG9/RvyB71rlMg2ixzwLSLjC45UFF7wg+VAa
uIoA4WDQykTUu/BUNaDrAkGuhoUbU8xYCRE6fdgzM7nra9jFvUlQpvFtGYMdu3uOpcIwsWsQULgc
gRDO53UB9tr6/BAWQzhIwRCQVwZ2io5Vp7tJMmFX434Jtw0yCZlogYc/RHN8UjItXB24v0MrT0n8
RS7Ty9c+czydZCe0JZ7ogYXbdULr4QzKQSbOw5zy9Jx6CcLKjxikNx/WaCQV/aTWIqdgEzNJ5fue
GbpZWXEn6U2xJuy0PAQdLVArLCqSq4Y8hEqBrSSZC2x9cS4/RkvxbJE+ODk2DU0AoZ974F+ePegu
il6yHvGEjsH2l8G2v8kMzNsqFHLaS/jXata+JFmdZJO2UchVXHNG7Y360DmCc0w+uzkiRpRCLqEa
bHZSYQl096wyxeWhHlrlmpzAFvIJ2XP7HQCYNX1Oqn77+z7S36pTPuZoKDxCt/lTRvU++NizbQ8C
T90K7MoiCA6vvysbIyvkOt6+gUIDpc+2Ebn3lMXB4WULZNrldlYZWvN+eGFw5he5fuiyhVdfT8Ta
GsTy2dXwZktli1jKCpsJ8JIUHZ5qnri7x2l4mSYkduEnejD4xkK8J/RsyomMt6srqpfxziyn8jqf
dNnxqM88+qFcam8xkWCaahnAiETnGJ/Wt6QPguK6ktNPGXAGqfnO15tvNzvAE/8GaWIEF3cmIRGV
eLXz+1fCJ8gXxhUelMtP9E0bKorWPz7vqWLpd9anPIO3Cxd+8EN4B0nSWU0GONAyJNpZOOm5q5s3
oSPvuWA9kHTQRXbzdguPELk8eIUaff1fiD1HpBgymJXZhr/Og+OXMc6O+9L2v+CQDk4jDBVlrmMf
X1x9LeFnFh/hj9BNW27KlpBim1a2HvxV2iVZizYCCdfTmhF1NRwVvx/QU0Us9siYXb57uPQagfrO
mDLIa2TR3ulRsYVzMrtjydxDkd67Nu8XAgg3HEnHrV7EE4Ad1EIJYkAMSY9eX1lKeVN53xA/eBDy
kkVdsdzvMjztvi4mjLmUBno78HQQVmTpM8lNXvzX0qyMW4LNq5U+2Co3zQIgQF7J0tJARY7yzNNt
O+26nrJHFQO9y4P6MHAJEBJ584+UCV6SfPOPk8xCajDnB5keyyQyewzFlgt1dKtwIBx75AdAWEUX
g3dSZE7NCxa1tMQcPVfNpivP3s6m0V9A2JgncZ9oks4nnjz51puj1+LrgimRE+w8LZ9/JK8PlgDJ
xvHvU8CERVNqdzwh20j9a1BvJbNqAhs36PxDviAUysG5MqC9pMq6gUi9HnZ7OCQ72oguKR+j0XKI
tdXE6cj6Eswet7Si6wnZzJV4Bqq4j5bIGkJUHU4AVWIYZK7GiTtAlMqfFtLs8qtG8Tb5oyObUYEE
gaXVohlA8cH0ZcqJWJQwgnbA9KuwqL3eiNzDGhNZlRB+RRLV5ya9ICsLDF3FOUOrh56dzmI4c8OK
mU7VwfelF+9vCYBwu4+MosE0ld0paMAuCOW2nWsC8iSjoPYvBQzdTId1Oq5vbwZoi1gGNNUxnyJE
9/wEHX8737uzLp1uy9KNhalnYKTxNcp6BbpI7nQwHHkm1LhFyx+oPIG3utey9x3FBaP/O/CmYSXV
XmICvX6/Cbu/iVrYi+TdyEqjNDIgg4wq9w9t6r0gjEwRoQTEBpnadSYeYDeylDawa8bEBdixkR4q
heUHVwhuEtCaX8//mQRg/y6cFD7Fv03RiSuJa/s0tNj9urN51GMVgCMg8EF9qdFC3DIDZ5BQXvfO
zumaHdGZVL18hAM2dpFEhzdr8ijDzx99UO7GdK4nwV2r62Z0p6xhLooqfWZ5cJ7yNlI60MbeybLg
ZktrBe3BfxmF8raabNpf1lAcU1kPd48i5q/VT2aLvZse77oD0O7o4UQCz1QGBcG3AcOMoPTLmSkZ
l9+7xl8SN1AXGVhl3N4HSUMyYd7hxMfsAIFZT657VWIr5KV569NB3oGBuyY3X/krBq29FoAOXr9a
ws//t0ptKap+K2Ly1+BgaqtLnJEOj0KLgQs31dzugsXNa+S2EQtztO5grt0Vdrj3R5handbLNyE3
JnW8JaZf8EhH9ANvCm99NlLLqUftOIkJ0HKH4JGGnDPvlsL+N9NA1e9jg4w4mNhLP6pU3So1HziA
7xSaaEOTY8Wn7fRKCVKbr9cAV5oKHwL6NZPl1yI6/JNhZyEuVKdsA/ilLXTMzhL/IyWEvOd1qluY
JKUl/n+R2DGn5Ds50WjE0hYeO3fbN+Su95+8w11o/J26B1PN8dIcTjUTotyaI4YzRANF41oKMaaW
B4ADK+93YmrW52abXAsCxRKi/twqVtbh7BqOkly3EJ0yf9U7jX3blJf/kjQDwlna30aWdWSGR73K
LK81a7tfGUuZc0ZYvu8iktkEcAa1o1BM2mSFheT4eyTkol0BjnlfXKGT/NmkmgDk/SZXkkSwKScF
XmXYs5kWgyGksrF363EBM/JJCiKZpFcwhz5LDl3Zb9kzXb+3kmaIrhn9CzlVDIjfgJbGVZHSfk0O
CVeVvc7BTzTIrc6tsnYt93kPqiybnlvpqKVrEYzdeg8xO2G4/rHo6DPgaj8U4is2LzoYBIl6AuRf
6G8aqHubgKMvuOCNz7/SyOTzmx1vJeYzUn85EBDANf/el6rsM9z6v/F1l1R1xmE6Foz3dILUfsyD
GwTcNgJ95IYGULqgtbPsw/xqvdwIqyD7o40gvW7s6rgbGAwfWfMknk197WHJ70kGDJci0XSxUEv4
LfRi5RslKGkY2b7bkX2p7ENySutQRnckf85RLeupVR2xcmArih5TvjfRAbrOJ6xq8IfgR4rUOikE
ve7mjnYTtY/WUzLcWFXtDmP8vRs/zsIWiOqE4kRSBysuu91vy0kYDjiHukIVAEu5JNKSyfyvrRRI
TBSZWpdZQWkMKkQVV6pNRIvooYM9iCi+SduWoBPgC6fw4jFLOzKBBdA8+BEjxsRpKsvOcGeApV0F
DpAeKauXD4LD6R4Q0BZep4XflEHlr1wzYWru+RyFdQV9lqiN78xFLwca4XXmRMpxGgCge9W66LBF
dX6ABfc30A0AmN+Rk4IVF/LPlcSa1/JQPpII74O2TAm8WufxT30uOqZEZEG7nUR6Qt/7NQkfLpuR
7XwrGQC+9IMZMC98poUxlBB4Jsf8SdmS1TmZTgIRZj7KyrC/xuDAlD8KaxVMCMCFQ3VE1oC7sQRI
mYycmG4ep+hnXnsEVyO0YjXqvgxMbFzdnPhiqrY5xUkjGpmw9ghSmvswdTiG6hpwND9E4mJRiaxs
iaDDgGb4DI1RFpeOgm+f7QbMzv+nIjn4Tp6In9p59W9J0W2q+B7wtZJp/GPvOg5JQ3x3miEJp22/
7uTOWicFG9V2OU40KekvtuUnJ9SAmPL7h+zHkX5neO49o7l0Kd/CwTiOZNrEi86xmw0BUq7lzKfC
+L5zW2c6lzp7LXztmCVX/JQVeZwxMZ2lFC5NvrdmjKexMXD+ovTnjfIKUfcSu/Vp271EJtry9zbo
hZtzdkt5/Xv27G1WRTmng/qAMUa6RUhDzXTwyxyuVt2TGJX8CvzyPnfrP3ytVPwV2sJc8USeM/He
NxrTI/9jaxW1MQOpuIGyRS4JscN7RDXhQysQsNIrDO7sEOvRkZDZ/Y6I95NRYRMW09cI765rJOba
ihQ+AVlmeQAA3PcZOU8UilCe38Phw22eMXI1Txfgi3SQu3AXHX1y5TyW7kwAQ0jwCSd284eLCW4z
CMFaNlXHwSTW8quNSKPY5j1j4DyaAEZ0Cc3U1dmTHVKDLNumH+i3XwPse9Anp2wbO6UE6Xx7SiKW
etPs8RJdk00JsuLPcoyC3Lv+hk7NExtLALpAr8c4qfNga5rfxyfwGc1cK5ugg6KkXiMecZW3hsJ2
VWBE5ptRPfZlXtl8oFRV3oRHOiYbXzFSETwG+j3HPL7eD706rOHgnPu3JoKVeEIOmkp/D5y+4hCq
NcWiUx5MgLhA0EMcT5pE0cnrkzTNYFsvGj5fxezVU7NCYWwWHd/7yyJQq+JwW+E5CCSjVKt6ReA0
1HMR2HkzmCTsnLhdRZsq/Yexd9YSpEJpkJjAnboPweh+0mAtdyS2gtdxCgCn2r/EIL3jxxiaCQHA
6xOUPJyX7cJbA9W/aUv7V53XXY+2tgO3RQ2e3DeoBEIoirxCTiip0r9bcYD3+hyQoNbLufaSQqo8
4qayGudoAbHVpyyaHmzqJbOvPDxF0X7NW151ubi8xX27NujH3sPX0oGxpKJ2rMKwc3OY1gU1lPo2
Sbrthv7XCfO2APp2c98FQkxndgi8x6FPQOiuwmHhnMIhrkzkcn+T1tcjzZuCEUZRIlj9IQIZVnJe
KD3ftfFgo5hAl1e6eI0uGHgNJO3PcRH1fnSmywz/sO3sjIO1HYPq2Aa6iJKKEDlyhiFZA/Qp234p
4NM6w6k0hLKMlctYDfsTsFhBC/VTsuSwF9prW5A/AoOAOlucBgW55qndpQNTDbp/LSrQRu1TAnla
68/6Hohj3LZYELefZpSsXBCY2Thx5Jod/yvsN/MEbyM8lf7GORPGLlsKVHTfvroa/rxTqH/9icS0
PAAUSe63uS6c0n2wGJrO8ZnvBJRvJyjoEK7cxix6rRnxJQnBBXLxbaJujLHk4jxQ0lK0QVNnmX2g
alG15ZboVYDJxrpdYKa2fSceTLm98IZXj86XFTQsnm9IqPmgPyv4hWVyXNEVyplWOnTkU5PZ6AYW
HIT0h9N/tZlEiqmzk9KchGqLlCluthThAcuvuyEPG64xprsDfwdE/Ss9lUz13kbhyULGpotrlsff
CoKAGWpOD1c5PpKwTr5kcawat++1RxvpHurmTIU3FqggsT362ejR5j1Ubz+8I/oTJ28988ftc0xY
t/i6Xl28tsCBruRRS9iHnLV5Ifb1Sh84cm91eS6dWdV84Ro2fndeL+8bDvbIucLEs/ZcubdNOyH2
dfdnRqP6LeJevv4RjeF3G9FUP5HvoGfvjKXPa6Mkiny5iDW0xg0udelKx2bNaNM0u7xtq0MJc0/G
I/MncNA1hmf9TyceRdT0IsRxKgIzVEX2tvqsk4NSNNm4/km7ilLOcDvPEKh4nRFuRtpixran+qa+
qDdQ4FC96eW+D7eziKksCLdlcs7wzOQJRjKm5uNGJ+pyvqgM5FWF2aG0Pati7pFXcww/PDNb04Sw
tMl2ovu6UBVMUqAn34XsTNzKWJgmFRFr67M2rbXHJGnPvZvr/SZM880D0UaGeBKaaSZ16g0VhICj
6xgwdRFOFWNMg7WShOtDstFRaNP6hjKOQI9QYeHDHNYWemKXB6UIcoj+ofxgE6iMqs39e9+NFrWS
yvoIkZUqol/BkSpzw2BfbltZsH8MjbLJr/fe6Zq9F9XcoKPeV2etrUMQnKvnsEldOa7BlX0MkPn/
6yXXO4K+pkFbStCBtHRj8MZBT23Wrm8o7dcc9JQJwyT7DViKRmbuHguTlD6xGR0PMEYtbO4MvqD8
rFOspgo8XAQY66s/6tE3ywcTUpbIHJw79PhUf6PUsaTg1K+45LuivvGXYlE7Bqq9dvlZLHtoYw3k
KnRLUSOciezQeqP2qjL1gWfQNZNgbxE3ZWLyiz43sBMNMSNQtkZ2RyjBYd/hN56PE/w8H61g8WvW
LrUNFzTq+pBHvcu67VLTIbPRyKyYiV8PEKHtdqjscuxdvfcWldWmIe3JVbThpMJCTsYQaauLbng7
sV2oKClirKwHTDje01i0H3Rrxjczhdfc10CZXSKzU/mSntL5AsLA2849OU9V2uorNrgvjBvm/yz+
LIWSz/O+Uhiv54k9DkoFmTIjFIRKGcEaN1hxf03jVK9wmm20SjEJsidrr9VuP/unv/aFAwlci8QB
GKucswH8G2SDR1VBz5TX2a+QavrHZRIxd7vo5ZET2WanYUnwXVBD+SmYKby4DYpP4J0tEJodVbad
JCjCHAzPz+OtFc+XASsNR2Vth304rlklFt3iGdgit8Cq435Hm4TxrG7tw2yU34ErGTMkC4vt83DP
X1LWDZAKX6Cv1KIcwH2Bo1wGdEcA2ukvZSh5Sj4WlvzV9bYcEhtCPp/NVkfkJHhyHV1eDexQcGBB
kop8+yaYCsVZu8CIV3bteyErjZL1Xn7+rFtLO+/e8d5GtfwBjQfAASJ7WR4ULUh/MSlNUr39Xe2C
fYhf3K9VWSlUXx466oc6Tayete2921QwQyDODdIHG1eSfxYeTUX2aVB/Yo40QGlXMwcRdnS1PYm8
IDuIcy/jMMAZBcqVv2Ekdw4vl4pF0DinO/vONjjHkLBuCiGqMPsAgNO/r8IdFYTCy3TpXVNVVl6k
YQSo4/1oxdKyJh/6b6T/XTKvx1ydZKtK6uE5EPcPX0S4+fHSAwKgRZHy8mBxH/NKL6XRmdYuQay1
2DUi/h9dH7ZO93i1V6tANXwKJHXR2u2gZx0NfbbaEndYhOJu+/OB6yDo4HhFWFJde3ls/6TX+h3l
iL8MnR1gP4pnWlTFD/lsKiLte4hJ/IXpdtjGgxd7yvHfNg8ICL5RGqrOGjwb2LE+XnZ6y1fiKWSH
CMF9QMv1bLm/oyTJUN8dbCWQYwofFqvkYImNey34NBf06Zke2k9/vzmsjo9cn/evI+DrLOr0hVrw
m/zol6eWKl9Wh6ZeOBLaUrOOO1T7HLtLlLBHTSW/aUohR/ia2qP+C45e1BFNNP/9tRqKSfeSRBzp
oB2L5a9GsCLRV+YsOnitYXvCxzUN4dt1MrL2KnQpvoHPAZhh5WlgxIrKpY9x+nNb+rQ6pJJoFpH7
g4r96FxWYqQwbWNdafrvLooa/EP8DTvobJI2kUKLUN5RdG5jS0OGEiWrw1+l3i/hSz7DAgxHXiLU
axLHJJqz/Hea4s2t1lQ9O/ZMYxid3yj2ZIC7HvpwXnjnxkoFjVhXvjwd56dhPsRASBeovEyjJ76n
A6RRfPGcqH/MnYjdlbRHO17V0KV9drBf9W+OhSwXpSdd6hobn/+4ynoDrwyJgZcUOqkm2Uoe9qFQ
gx/11FYsjmGpbK3IH6PRbmgMQeNbxtlmlc0f+7/g5HBCCWllylwDswt5ZZVk62MMplhOi6OYnoTv
JDjARHdDE5XqO3di3nb0iBuxc+8wFodw6GckyCLihqLokiPsJE1albxFxPWu9zVK5oRkxVkm/JtU
bYWHn6AIHHhd4xRVp8beqEl1m09SaEPnmsGvRpP08gCZD2KAU/VaXeCeg3UiMBI43Vord6JnQDRa
nLAC6nau/5AskKWeeEfGn1TmFrPHD+EDiqM6XqLYAZWdcLj0u5W12tflFQhjn+5LusaqkVLZq9m6
R0ZHwbe5iyHIfiIyvABttRrTf+Fs2X26Os4GL6zzK5lNsOqR97ehBZ8Z4pq7el1+zstH9hACjbpz
vpSRXUWKUs5YdEpfGzRfSRSwKPiJdZtx9yHf6GFH04gNExqSxjbIMqjwEdDKib5HixC8whgTsTeR
eA4hAEnysq0Jzm+fd1CDxIMYiEnKPaWIOkOMotMme1eE1lMReNz93g+qzI5vNPPNqC4iIZM+GAbw
j4xk1powtILzghE31JNhUy015rT0aUM22HOtOgfD6x2QSU+jzHVEc9UClGyoIWwcLMqPA6/6wUlO
LcnV6HxnNLTCqNy124O2BJFRK7g0JnmKkMIoPsJLBUn/7neU2OFGBRG4L8ngtWdrcV3djYEjbtbE
AJR2rvQYq9IyfeA7YXKC+EHaCSpdoiluvvH82ukcWDOyN/J20xEwIBxXuei8iUNH0zxOu66MB3xZ
Hn4tNsDVtilxLwFABCicOe+FbYEeovyApwpXlJ3MXGUjX9kFylByUxUpGQyle6hcIyo+rwif96te
Ql48xywr7N95kukxBcTAOvmjgDSh15O/BYCT+0eW81URXDUU5TyY1H2QVm+6dcTPbV4gvwrGMSAV
m93zZNzTQqGZ8DFjss4W71UXB+CGnwaFVk9W7mGXi2BVokge+gdFmwhau3TjK9JQ8qfLM0FW33Ax
amFbQVwtHfUEe6VIs6+MJS0MH6MQ7IZpW3/eR0fZ8NF3xhEGihaJxNewgTSa1FtsYOnbGATl5v3b
OPu7+L6pbx9IzTuQWGaXQCpxKU5TBRGzS3lMLreTnPrn75lxdFdwO90bBOx8rBvNA+48i6T16rN4
BKHjflea0oqu9tI7/7AnahcIpYjT8+JLEAxJRRFUUtc0m5nOu7M78ndtryDdhec0/1qEnh8IjajG
cCyAtAKLsNBbfBJgXtMbthMSht0HS2btvvAmVbltfjNEgFECKsHakd9bUIED02NGnQQs9+JCUpyB
BvVGsBUwjUGXbeAkDGDSe7iHe7/u6kq2HMuSvmVRsCqka8SGO7Cj/uhkY7dudmcdIplZzOmAuZmu
1FoRKAirwYakHVGTm8oz6bQFJHARNbDFDK6yoX3F79AaqIRIxsBK/DYOBRq9usj3FlIIrWvhXiso
NbvVC6mJ2lnOzeykfLEOKFKlaFYWGu1j89P4acF+Au2hMCzkWbNpj9YMAy0UNqBahirfiKlAA4zI
jX9CE8HDKFCG0+NMTx5re3AXsuo+VQhCv8LUb47/vyii6AN24pj+fgLHgvObeGLeL2vhT2+Ojj/b
GHZZ5teomkA9oVuqynCXxpwqfNn6pGsk/wyVezqU/z0n4pjwr/5cwttIMvsB7MyIALKQcFzvpz1v
wZv0Qch4m0gvrQiNLhmXyMRf7BQjiaQkPk8cfYYySCDqEROkTDb7UHpngmiXsuh/6QrLjE+Zyb+h
OLg67aU84ynEIl72xAISY8nYGRe+jlL9fMLPb236vX5VhvEPWyV2qkccex8VQdcZdZys/4BnyrNb
dLSmyTG2Qyw6A8Wfe9D4pJriAKoYtOq+eq+m6GRRyJNV/KQjloYPb02xybu7DMC4735eVQB6T/PY
bLfC9zDxNEJ753mUYcd8b7UCjA9vAW7fe9nh+CcrS4LSigsQyJ64QcfpM6rYBP5WdRwrkiKCpZUx
XfOJkoFzOZiJ9Kvpyu249l/MZmiSI/6gQlFfgPbVg08HfOPA23+z2+Ty92Zg1qXfWSVuZLwGzWjq
x1Y/CRAG+lc2NGeCyR2j9wDNkEx50I0QYbE6gCurEL4PpCqn+p+oj3WRD2MswpijSPCrpn8KQNkm
PaacxbeeLYLi+TEBqzZT1GFPkUSfkNSO+zXkeEw5o+vivYE3zV+2dK2gyN/14q7fN8ibhYmbMST3
Wuneh5f3qLkV6Fcig1LGt6BYFKKx8wr6nbqMBuVkTTIIa/scWhyFiq3TWu3Hd3IcKR1rhaC9PAYg
y0fhZgTkkgucQzOApN4an+q43E5wwuon9VHzUdCETFDL6+TVjaZiZHT9ZSSBAlfb2p6r5PSIUWM6
hnPI7l5hkaXW7wZYaPvFnSsoXCgVEW+5Uip9mSFIK3+CKBF2w50ZgOc/YQVW5P+n0ZjODqNo2/Y7
q+4d/bKO+IwK3bKL0byNYitibXmZtJ2e0vr1UBawAjHbk0SGEPkU0a/5smtfsjQYLhe5isZ9y8WH
DBzilJyI5TXx0eC2YA+2pxzG4uGI8DATNW9eK/FPYo1ZZU7V2dsX8TOVH85UooCby2nYMmaA5rTY
8aLoJhBONo8Ye25vK3avG40zYXhDS6N0tUCcmoPuBYxt0kWQX5qaZMSAw41B0fWEgdG6xx1B+QDc
Y6EYCti7DgR6d+RahawmKAStsNP7swj3Fdk07ch9zxlxpij5VsrNmoMoVEBunWDzTpONPfhX4iNo
6kdBv6/tF7CbI06/PkEBUG8ziZwS5e4Ds3KSBW1/7Opi462F8EZ4EvznExZdVZ8OP3HiLkJ91LmP
MSuhbuqXWbVzmCmszRlTI/1q8OS5VLhFSqzJ6nhzBEgwaCbsRsBru84kR91TDnBFDH2epsBI+cKY
cW8aMawSxUc8GDGeAjtC+9dbNxJAQqU1l71wP7rBC9OCWBDNlRmkTmrkgi9Saeocimlq4svGtXXy
bwYVriVNo2bHng1t3q6xXOuYLc6Y6oTEUsY0sgzT5AKnT82kXRZYyiXmRI1NMZZiCN1a3G0uXI6C
0ozxF3ulJgW5w4KqVL0hipFDCVyGYBmPso5wMgQVo+4Et88C5wT+gbAsdE4SDO/Ni6SRJIiftqy8
zLrsIJYM8qrSjOa4r7SGZ6dhRJX/RWuRjyKHFUcmxy0D4XkMxoC4WfDhe2r0edKJrMPpJchTtPza
4BzCcvtLd1e4oAi9h/J1/UGRGrBpmdRsG3MaGTYklB43eQPu3wY7su/IgNJLSG3gFAtwrydQmW0O
uRVLOM3+Fw0kWoINb7WuMPfg5u/h0Eoo6GDPgAV2wevtw+/R/jrHACxFJflEKdgao0IY9QUFoNSd
8U8msV/QKAM1/wH1T7aCKSDwye6M6Y2UaoR8quiwyEDEMej6182vq4+8emsMqE5YoyFXDSGdpkiH
IWSMqjBHiMVX8JUJ37LfVGVDY7AZqT51U+jlZFhmJngerxEMgwJsYgykYQYpjU3vGumIQGNPnOk8
Ou9uysxKKy/ebQVVBdsyGYVXLhKy8lkqEw0Ye84CRypr5vnVdcRH1ftnaqK6tfDXP7TgIaGiJh4b
qFy3xFOtaVUTW4tMPP30SnDnXbcUUFBpAGaN/c6boR+kfgL9OCTIzP4P0pS5AQHQCY+EnHst1jNz
55WBeVK9eudJzGSD2OpuCA4SMm8YFntUXnVB+v4ekbvllzFu1QWCjHXheo3ubfr9zIFUt/p6Q4PR
KTCqELl5UVE3Vd70bcNpmCJ5w0Flp1bVwo2fCrsbD28sVSJaJNyRW25MlGqz5nO/G8q3TbWpPmnJ
or4pKIBgqHGKcdXVnWLdJF0+tXILzJniatnYAdm+zNe/mR/9MdCNfoDfaKc4grPSf5rbCsh6mnwk
uj6twWG7QrcahNzNpFbR+jJPFxw9r0YYrud/viUlyfiggcygPCApXouKkbehByh9oUP2cEeYyLSb
rEi9jR0U8rNRb6a8RVldvoVzGGjGQQcrtBwtIa2EWfKv0UISrbSuCmk4LVB09VnWgOh87m6X5XGZ
auBUForBzDV4VqqZk0e5hr0nlDaua4P4YRK5c0BF5nryK/A1FbEn3bOaPOD3i6CdQ5vv4UtiCjU9
CQWUjLStQdkfubeMG2Utlyap9aI8o0vE2udLhdToVGHE6VVFKZMtnmXAboA0y4awmUSds2Zy8g8m
p3ND/aC+8tYAJ+KoQRgkOxY2HexRi3ZZCpA5ZqaZQ2cs7yP8z18IGhGUL9p31EuCrfXZzJ+8PIdk
SVAjNkFLa/Ux9b67qyKSxLl27CZUYG79thXYFDs67pJX9cQgH/Jl7ACQA468u+U1mNn1+srnHbrv
Zq8yB1dsWrpV2Fq+qsEczWWMoH7V5XuBkDr+/+XBqQrJDsUWMA1JU9OXajpjOtGPzD2QgulCRary
ucAMAn0yATuUUUcgXxwRflIm3Iyq+wG4R9SCVf9fZp9qrnGWP+5ifQI9KeoV1clueP/2xZbW7goe
mndp4UJwQ8ADFM3Q6ylPopvGE1hmSUi8kB+H0l2WuwEc+JFF29veB3MbxS6u87OUMOsQ0d0mtZUA
XEIc2mJiCP7h0dPDb9itFYBvMM6wpi+lU9P5U/zpCzB2rjcO9zVw+CA0c5WzNST+P5pzIqy74L9y
mFUi1mu1ULraJQ5rB7oROuju6P2QWsvlVzNUOBh5CDPFQF2xnff+xNry7XBnDfkDT08p5OxMf4bV
HwiWpAt3GGq8vLQGNcwNYLfBbNJ9hT0NGE6sGo6HZ8pT1opsvkD3jyo0AanVraOmn1RU3n5b+asg
E2aN6nfCL+rc5QrhfAjBx9oldnvhj2LKTSwCJWT2Rq/YcByNAlAv1Vtu5AWedYezc20ec+/UIkVq
JvZOOAeeEcwTJ5Z/bJPi4XkgiskCxr15vqxeoY0kSAFcEYFPYul3s1m770W/Mv/yMMKuShAnFFnt
xE8A8tPc+cZkEFsjZvZzhfSOT93Bd7WkZLLy/5z06770xDe5jIfDGrDphahxbyvSY+zjNZKjFrZv
y1b+V+dKumi7uJVgyqon21hCdfoOThF7dqVlE6sq6rLFOP20k9XPOM0jNa0u/3p7WemCG2vovrN+
3TnB0WYVRa5709dxiqQAjlbToqTEbFdxd+RANsSqs1zReoXq4DjUzGTvDwNjf9TD7/anWNbNU1bR
csn/daHt3a6VfGB/ENLHSsByEBmjZP1X4STaEFDf/0GIVACQo6MFCTzcY5bfQb1JdV3z/+mH+qP9
odVxvBMval+k6pxsnbRyGnWt0EK6LWyQQeugxQEcnvivsoK0ua+KTEC+Xfso+jXy3xg7J+Gm5vtG
CA5BnqIW/t1fNHSY9ivMUXQGAYtwLtSF/ZyD4X6knlzhEfVFmGIpown2QGyhDcr47oJQHGlGYdp6
Vdd//XIp5rSn0g1TUM3zXSWtHZ1Fhyq8WOUX7xyef2WulmRQH3bDB31fTSHZS7NrBrBnajSiaPPB
zBp7OTrhgi/8LlLTbCw5Dm1ZBl/zf+l86K4T21PGo+lDmRroZ/HQGoGX+h0UGYR5sJY7EWhLP9BH
3U4z/tdGdR8J3nm9WV38OASc5nzRdLst6JxpfGdO/vCFLCT3EQZhnyEz6v+Yh7RZQkSUpFuHO7f+
qEIAfLDOVMHSTTY5198T+69Ym8tyj+O6xNIuXQkwEhkmCqP8cyIPsEi3ZbM4A/BIm/HIht+MjyCD
zw5bg2t6KCMgqmDjYmQ79005mUfUGw8p8Qp5DPfMbhPTozGHM/EcWXlmq/yQnVLXp9mvRz4QZ4lu
SixPTMwmvir1uJ1M80o4Dhzo0BILLZV7vWBPLycYyRw103Ls9Z7YXjGhOOEiydQJgXYmCIRzaroL
vu+7eszOsHUB7M6bZLG+Op+P29XvnIN3AgyW4qqk3CKd7C9M5Prhc0yVfbLs+enLZJDFttQmCMol
t+0BJN9OcsOGBwwLf68sK9Zkd1hgm9PaVdznBf8hdkomhBiDK3GAXoNaFORPw4YwvbRVRAd+Z83B
XQlo8vvuePAFAhyKkH/kB2W/QhiKg0gfPFSPgdGsLY/LSBuu4izF+/frHsYJuP2mRNhR281MacFA
avjXzGF525/E4pW19UPUJT3GoZPHzZtasKipTY9nRpE7x09BxYYYZ9bhsoNPM63cAdF5tqiKUV0I
GFnp9M9k2/7SBvpcw7J6Gsc7f9aCgiQ43X1wsOCcl4pCgPPYMX15QtdxHJ21M+0NVqKXk2nCR651
OmbetZUPtVM5w7j/P9aour0klRSHNYvqWgukpB7FqpSkFYwfGsubqeemO/y2t6revZflUJuD+kwW
4KBNId2BmxN4hm2icYpmHbSlavrvY9kyJ28jA6Gk28pv9D4C4B7H78/TYVOwU5ZR1XSjWvzxR8rC
6uQs0LGRKlw9WseBF+oeIx5ksG1YcCM4kZfLFxnQqfDIJy5yxEQ5vKfwB0TaMC5yuJC1nVsV9Sw+
2J3izoeFyomu7mt5QVp2oxKt0lPgPmUttMu27uU9baPrW5FJK6KYoNmym7rIz/VhP3tokvYeXPn3
19sVT99I99QMMJGvqPjDV7GFcWKz4/AHg7IgY5VseALQIzl/KVyglWR0WmIAxVaIQW7cSXPbNP3e
6gSQ6po+IlaNDUvfhBCRQkicudMZENzzlAOgmqbvZUOmBHhhn3NtzZFvJtebs7Y4+Z5zWKfZVMw5
thRPkZRZlM6nBF1M1uSoMVnMAoub6ycAcrhT8jBuDWMUCSVlBF8naQev6ApWTEyFoVVc7olNrNLB
TalcXCC3koa2SetU1wiCDi4ayVFv8AftCB7OsabC7S4fF4RliDE9zCkLvdvZANMMwH3G7EkLtQSN
FmF17wycpENztIReg4DuCZy2ptueLCeFqqf+r/I+pECELXjSbYkX14+e4piHHp8plOfTjqj+i0oT
bqR2dGAJhUpCgxg8leS+HrHgyRroHnOlGt/LT1SZzfi3WfE1vM47TlJGF/AUiWgp7Of5D2rGMGGX
6v/HN62cparckm2Dosd8hHKpdjPcj/JpWKvvzh4tLP5WHKlzZZnJRfv6uKfCXZqOHCb6GiGtPkeM
WwJDTg8Z7dxg15eaBbb5eJe2oVBCF8DnBI4xLJ+AKUoob9qgTPI6KGyRrE9e58p/UYkSU/Pl9wSi
i3y+JwRuXYXhYLX+YwXgXwmaHtjUkqFqXFLL3VIVXyJQf5IcDtjL6FsFhG0uOFUJ6bpIZZw65QWy
EbovdwHxXMOakZL3bxeHq19qe5ATLMjcBDYV6GJXNPrbIC8XiHVD6Osf0Kvcou5p9UrApE7B8lmL
MpAtuhG6NOziANqIj4mRq49FIyUH5cSadv7xOoRjEEErJq1F+idUAYBWba1Km3Wr7uCaEmYS1+Vg
HOuLgB7mVQnjonUfmsk00yo85+lHkvC5WadKAMvZsTbjt6S/clwc9AHAqHr0cB6x6xKZG8wYEtZz
u5VAiNT5VsClQFL/if4APjp7fQz0mZsFSIMF/PTMAV0ydkHfJeipK+9uqjB5m4taNnrYFCSA9Am/
rrXqI5sNWAo9vdeB11wrrDP2AuraicEraTDIkJx8GB2nsksp16SkOVZUagKhCQ6937pW61s0xTHf
9FCV2Kh+uaWQFz/iY2jS8JzW4fHwij+0m0HcjRcjASrpvH6NmhbCJuJzQ92/1uLqnNGTbI9nzUxD
r8XAusjK7cRInESYiL8zSrcabg/uHyzdxZPQz68RtE8Ovj8vauk4UogISTggRlDZYv1+QpwJdsKJ
kT+FFFjq/a+MzUBJJNCU6T+jXsWYtiq1rLTgQej1PRP8GDUAV6jyrr8dKDMbLDiatJeE6kIn17FM
lLBlb1DO5G45Ju2DUvU47mGK4xXWeybyBMFbI+JoxQoRw65PJRkexq0D2gNCS+DVBu092rj7Etot
yAixViCGoP71vn7TSNUcdhMzxyh60OSY6WSitF0TvMt2DVagQxhUODZezkflZDZ9YI1pqGPYPWsb
wiIUFLC5LteSXrRgJZCfpa+IJgCz+s4Q/nwV7tmqMHSpk3lzobu7aT1XIAuzQ4dY9Ktqtc02KTHZ
gFI3Q3rJmAJHv8zmQG1eIKxQSNNZd1yCU4QMFE9c4QJKO+TnZrKL8u8L7k8ds/GqXwwm6XK1l0Eu
4Asb58gZ4Jrq/yWD/XvCap2wSaK/+5VfGqeX4pbVNFxhxHoKgIqPEaAUfPDOrwv8qkUc2Xk1BhSA
cYannMilr+Eg27jWK0hizR0vu1npnrcdzRebvB/5IAbtmTzwBxIkCPklHExERWT8kGwy81Ij/k1T
XIRie1NL+MjZccatBOM5ZUO+mUdE8yiprl2mIvy/5VSj9NlTK4d0iFJ79XZWPNmSfdEE0Bd6voRi
xxnx+++k/H0wKnHH1NS0rOIftQFmEHTjDSYVE/Rwv+mJd14JxAryYqxN7Ndz+hB07SCAj1rEBxRT
P9CVdRW0vD8Y2V8vst+fajg1lCAHE4Y6u6txZCopXomGRD0fUYzllVHQKC9xIJssDP0ZtjsEEbrV
u8h0lHAWZTeVsdvcNzBMVsL/fOc+S0eCeOm7VFuNoPu7HiMdUmEdURQz7CQNiYm05A4XJAHs1jc9
X0QegF6GN3WhRYTHP+EgeFAV80/TAxiWD+ATWhLtEUnl/O7Aq+djXpS0cF65eUI7qEk3H0SJaJN9
vN3Jc1PMVgK+chCWlZRKfZndeSL7jasxncgSXZvELSKr2lUfMBj57xVBpr38zVNDp+ZZoo0DbB/R
BkRBa21rlHzlX6VPv+ZsPMmVEEcWJKZdo6l1ROjCqSG/3Eye+QSWNGji033UMk1ppWXty8UiXdhM
PMj0OryQFoAUzxOA0WB8WmAUKbvVQkl6alRI1et5GH4kf3DqWd3mtnGB+L30UeBvQecaJ/2lvdT1
yioZ7JhxHt0ShRBxhJv+/6bkKWtgS+7rlxSOs6SAirYrm25OnJC66v6KoqF3Q61gCqQt54My0gV4
vSCW06aOlPFTa+3S64D7e7UUoNC4cR3BtEbDAbuAkM4iy4M1EY2RP2rnEWEBjj++76U03IJnhbY+
32k+nLgB5BhiK9ywN2gmVkIQOiFZnHUeXZkofMx94nr0XIkow2YN4crVThywodf6GEeU8SCuA01s
ESJ04EEXCE11turAb1Vo5Bj3raZ5OkXaUY0O2jWvhT2qEAbH9PUUTLxAnOR5o96mIW7aKvdBkkHr
FJ/vK3u2rIqYmo0jposy4+gyWMOq8j/AGtkzFOcL+klPI0iUBCEADuW07nastNxakghGJWgttV/G
nRj4jpL8JRcq16UoQkNaSe4OEmiJ36lYJMBSO2oXkVQ1ucOKhfHVOprMDhyEPOLm2If2vH72HMJn
tcx4LTXa4hSSypCxO051UFWmTFcLR8SOXs/6B8EM3OnN1vpGvV1LQDWTwvABfxPSFP6qpaeaAjvg
nOwgcgdJUfDrrRJbTuvufWCPRufC1wtdBU3rji5vxqSF11Lat74fTyl1BX1b0b5w8ZxcIps69w29
3E958gmmL3dsaQgbT4Dve8JM7wCrPUlzDuA7I9BBB4CVxBu8jms67nNsj7gnRe0DqU/mCXaC/jAS
a7ol38ShAaoThgYdXqa2Md/oaKQyvsxe1xCmCb51zI3BcQ9jRIVfgTAlrvb2ZEHYmbqc6LdOjv04
qg22wESer1Tl+9Wksxn65rxBqz0F/IqpmFIIY8UCM0/pYK9GEpEgdNg+QRhN9Tsn8x1CSw+IsCC7
8UeedKe3+Exdd2L8xklHxCJF1XSKK3ibGkLpp577FCZIY+IpDSxH5CukmLul8XycP2qLhEgWbuzB
v5zYB17kYpE4ULQFVrPVGwFKd0Zcm8NQBlMwd65Ec2j7OvA6qzlm3dRYY6+PTvqZORH6qFJUlVVS
uff080Gtq6v4gRiteqVRzKO1rGAFcf7F7o5smAMk0Qzn1ELczZKdTL00iDW2ins0E7d+bbvq6/RS
fmW9jF96evGlfPaxkVIsU05QQAciEERpXc5bRAnWhYqOACrExJa/gsOh2v0z/W4OvsOoSc/4lJce
QVh8kHywtjP7h5OMYKcD6+rcse6S2HFLzyoLP8YrX9onQsfSiJHTpNP3nzt+YZBVB92VFWOkK81K
HiPkTx8E+x9enuO651uiM51RX0BUiEgs3wztexHeLhgXrlRYTooXIQlVZfAAXDJBGipYp8+tVBVx
PLl4ujMlc5ufE56Jn0+B6LTjrDp9izCMvlVrx/H+tvwG1kwWVm4xsnq43UXV5agnN0cLkVEFUyWD
LCl7OjdLU5xLqwa5NAjQ8xjiziXz0DfXfUlSxMPBWlUNpo9Ru6KVtXxIkrR9hRjZ12jv+yfH2Yhs
TygWX8HKesreWfWEfyN87CN0xBBWp0cjywXLjdzRjOcws2cCnHFNZR6edxriT9duyOUkhZly9Fhe
tFVaNpZ9727/68P3T7JyEhnPQEC5SACXHzgmEtWKtpEFY9n2wVioPU4hipdx4iaPzI7pTLZzbR45
jJ3QrFI50nuX5Bpalb3BXaSxiqHbD88ULN0s+SjNVIhpANcVrj8DwqbkEa0tqIxYDVbA1fXQaPb8
0yZozE4ERf/SVKnJFpMymwn15vJNlT9yu8peBTOkOWoucY3lDNwulLoe+S+u01r4FcE8Hc/uVdDO
/pjTdJgUOc6ZyhqcSyII12dSGGgJrDevM+LPkO4o++vMMee7G7cw+G1XC1MbxmvQBuvT3WzyCe95
iOAe9lFwM89+rYKhbKxtedhem5RyFfUHWtcFP3AG1KLFT4TRxbdH/lk+9E077i0BQd5ASmcOuIkE
rbyMUXSVOg0f99MGZfenidULOL9jYCw8q1b9j8Y1PdOqrt7txLuRwO5tlRwY2AV6ZUM9hS+pZg5G
PaatJBVDsf1LKBodIoflYOYKowsCRj/t/+SjgYdacgB6xgFVPCzShI+G2vwYGjtXossqJyWq+ASO
vlJQ2X+3eY8tr9U/6E0XmTkdNrWVCA3DueKpXHdGHYWVswcOLFM4VqfxHJxYZ+7v0Lzj8cHwRk4p
qYVVe5kuKaVLpDNHhWFVNbuXXuUIPcLA6wrQ2t9WGKbnQnwVQsKMHzVqgF/a+vt+1kO2SdU2szne
hfAS6lx6yCZlWzJmdhgkUKgiX+4nBLMWoZPUwgIW0OtaDLevGEfSSmTincNybCBiRqIuF3Dcz8ix
H/m6iM86hK5vc9JkgiWOT3ZHVyuvPm5ZeQoErYSzDYXtEgDszfzM0tX9Q3iVNK8x7DJLfRWvLmj3
cMjCa6Byx2KJfMe51TZdD432WWHiIHduny8n+6Rd7+J4FiGBXeh0xbSiEPTMag0giX4i5FRa/DDY
ot7EO2oLOt2n2ki4pjJLcZDRzHR/COQJdzyPSQwjv2GQoDzxSU/uwTBF7qa0n4P4ZezXmneWUxnx
2Qgl/YQ55J6D+SQnNKoNzdcWjyecrtLFOiSpd55+3YX7tnmXI5J/BaNsTfehZUFaMSxfV8/tOPf/
qqqDjQpWh1v0JYJzOfr8X6vxn3sUm7p1dzd5YzpHproaL3GoCS6KmJWRG476oMRez1VIE9OBdU8n
hx9Wi6rjUzNuCsN5BVwsg8bZ9AFaZN8j6suVTigWcLLyq8TTeIY1LjDLsg3MOy/g34XMl0yubGoH
MuHVck3/zyPrQTvpTmkx8tSpO8VecWN3u1m3yxGDeysEZgmwjttIc2RDOdr/tezdoKHg0rKFEaD0
RwQCavAILg+hDEZHldzP96B18CILGPLhavOg2JDVjf0fCUcVjU3yIkE5ksoGeZSEyO0bQoMHxgS2
e+XWDm3hdezc8l8YyMasis2RNbgMC96OnHV6OAGJKL8KdTdDxdBdxis/b4ZLNNGNNtTQTuCdQVdf
0U+B8aR0yCeB6ge2JEIUHTOFRflMygRXZm3y1y/Ny0KWGlcLSt/JEdDsDZqtCfipNc02Nv3ua8fk
VNIEMSKCtx/r/PWamgi4zqrWB/GeI/6UgaOF0iuG9G8LL3A9ViP1Y8rviiOrxf1VVEdK8ZLLiqFx
jChscVS6mQP5A7USByk3vFVsSrEQ2rVgWPkzLIEH7zuoPv6IFVTcwFx4Q4Lm1X2Yz43vU0HA4BDf
M6BhxtKLa1kBlIG2CD/70a7fCsBa+6/hyx114apZsSvJxSwsNiVVNnaZHX/Wjn5NxwcVZ9lfnMpV
/+/cDU1RrZzeiLFxlrHFAq1Sdrk8JFzGOX5nfLoFw8vvmM4nv0rdOJn+VXBa6t4orzcUkSZIPIzK
EseVouVx5vQVfHvXS+2c4sMwMQd3G4BRY09V7MgtOscFbv4zjOYkMJRvCiaL1thvNY/f8fljXkhf
jfpeVkOubfUpzjI+I3vVjrg86b/8G0NtdAwOD+FgyZfu4TDZr8JUQejUtKpLFLHGQkxHUfNu/zZZ
s0WAzOW+oBk1nrgHY+IQroyOz+Cw3DWIUVH1N+3OVmTJRJwG2HPAyFCKk6Rv465cGRc/Yo+XxC/y
1LIa7yLSZgG+YOxfyNRpgsKgl1RUbQpzyurbGMEFKoD1/agPpzg11n4JJj/9CBK2Mth2qOGT5t7y
rC7Y3F5eeSDB+ZgHsloZtdy2NUJsNvmfX+pSP8td4KJHvH463sp8Li41fWyLJL/CrEHKhUrq8Nxm
pOzoa5FU8dXJt/Jo9+y/FTgGxbXJbzf8e/uBPxfV9mp5jnBoDBZcw+7verY9Umwej3ccdzWG2sIE
3YEneJ4hZXSywQl3cTjgVE3d7Okip1pL4GgSmkTuHpgANYUzgZWKOjjxB7rd9cenIeU+mOErNHze
rEPVwhwIgKkUKkWUYlDidWuNPQToCmRAstbJzp+MOY4UG32SuSa8eswmTPKg2Ha2s7u17IonRW5s
M50omeqmSdiGBqzVoSZTtD7sQPArd+aDNDkH3+jLRKmf5TgIrjgV8L+sZ8Rxip6Co15uXBQHnS1n
UUwGc81cWk9ePoqsjUjVNSbL3woGUnwKXfQ7S/Dw71taM8jHQuEiC+wJwO5wubiCaVFqRSTUgeBh
w/W5ccBGQTMvXIo5PSAJyan1QlC/g/TgnIAXtbQmyPqXOUSfJDe7x35RkNa2tr1ZwUTDsKTTE3Ye
S+7CEQTLVTZZSg/DQUFcJVxqHxsz8FKqgKBUMOnKyHUHY3k/xKyQJRfkb0b+AWJmwdPl4gvo8OpG
LTRJkxwEd+dIGte1z7ahPZDKMmizKDrLzIDcymRqAzi88+KY3A07Es5pkjWhQYA14tmIjgtPeqXc
t/5YOeLeyuNVsdUzKRmb18f2Sm6imRdg4hMImOCWm63hyvEMoxx+bpBCEk7vXMBT8yDjuaUc8TBK
pGtYTrH+hXE6nigNuYbzAsGO+FJWh5Wiu2F2Tn0PDRGVKcz6FZdV5R6zSx2zMKannYYoIY9PeN2C
lXSmjWksBHnGND/wfTVbi0au42TWpUc5dAAI7GVTl5eZoUFSJhuERMMZG0L+NX4qInrTOtZFC/Q7
OFXT38Eq22K5cN/510sWIuPX9W+f4mhjINdvoeDgDrMXE1dh0r70TesSmFqWzWvF0W4W+wcN84d8
QIoQQjakfGBzzn7BzfUaE2gDjW574Gzo8henaeiyRi3spFh2msP94t6peejNjOBz5mq9KslszjHK
4VyZZuevpHJe8Ho4vcQHssvVUcHQFrFgZrE2fA4agW+UwnixRGqm99kkO/gYg/z5EIeiM2cbiQgz
id/SNtqqGSzsBu4FnctrB6uzCtF9AqP9rWiR9+uwKHTo8MtvUj2f3FAn2SUm+nA3vNPBE7azhk5J
dJBJiAVZONiuX38ELQ3mhxm+yrLuv1q9Jntd/HM2mEFPyhYcvaxiAvVONfzBBVyi+g3+INO7raXQ
C45vqPxNrxl8c9bVAElJ4qiDvpJTTJiLaaDCY4q7cXPUXXq2h2W4tsuGF3gFoPGZfrfmoohpR+FT
AqOIN9tEMoarUjWtnWHnwnq3Q5AsOXSeKFjRqAR7+1hHNHqbtnsWiesB3JQ6b0oGz8yUMQP3Co/H
dlL8MIy+W5c9SWNGDDqFDMv14fJTO3IO7vNtwPPEjqI3vqu5AaLRe67mf41HZRmfHt5bT6DeXh0U
pjAGKgFZ15knBLB70udj50CmFkOA6dxCbjODdkJvYPnFGhP/rDbtikrXMkWarN9lqHv3ZQa6hpra
chhbRp0ewRbe6U84B9NNYG2w5W3etJkicpxtKDiu28D4gWXW6e5MMFdo1m1YrdktSqz+fZGSww9p
fgfyUsjNzTiOSGgBmLhrpTiFKrDg50zJCKXZ7+n6naLz0+JP3zvxB/PzFPf3FKZQ7Uut8WZeTGRL
WQ+bBtR3Vk7jKLjtAiMtXNWvnm1dyC5INlnGcaA+vi2FF39W4ep5T7i8BWUMnY1QTEUL+IboUdJ6
1kkBdr3igBXCMXYa5wpRrWnOpnmsWB2RlZ9e5ofxtNN28RMxiXYJfSo+ktuW2+12O8ArSkyQmkXB
t2cs/UfPhFLhOIlFHaMnwbA26dD0I7XpQa52CZDvGUbjCt4ept6MoWJ0aL2JzHomb8PO/4TpSdeH
kUDIihke3tdMrlMuxM+G5zkWAWEfWTx2LE72wHFypwdbstle/rNVF1Lc7yf6glmTONtbvwWVYQJh
BG9JDm1AolP6jrapAt2q7z0EKjIZRmc9VtDFbh1FhyZ3Shm5NzvvtA82bgt3kpCM4zQPxzRpLo3b
4VWEgVP/QeC4rC6jiBaeORDawEwGxGtvVY5dAgnW2RWTKG4iYJRC3gg3hceaLvb80sS3DNRbRhT0
DJz5LmEH5D3KEohRC6hn2TJa75llKOp1JiH0yBSlQBZsOW36jtc7xWivNNOz++QzZA1Lxly9k7z7
zDzajmRtH/x7vteTGA8EIuEApERy/zhvoMpwKWODqGGtFlP62xexzZ3iHzvyCBpaHln05/ZeCTaC
RMew/1RXMF0SxXGfgMc5GN7X0fxE9egERRrGJvla8diZwPAwqB0QubnGdUFv1NarV60f3V/+Kd31
/eWZZgPlLUMXSpLMNEAjAqGijsIKGRBNM2SqTJBYVPg5KdPjKti0cRB7uOg5yd5hA8PxfFJIpovV
FINriUVwlHg4fID9op0XacfM1lvzyHaWaSvMDsqDeXJn80d+itJRvowfHKQ2CD6fMlhKcA5F+ZdS
hCOO8zwmK3D6OP1EMarU9Eclx8OhO5la5xgVuPf2VHkZ3Y3F1eORenuWzIsAjxpzPKD6WiCHowUQ
Hz8N1gqwCEv3ezO+gg85HD40hqtVsdoR7oPkl/od2r30CwwJdNdFkKFoPZ6yn41mo8CKwrlbumBX
g1ggL7UNlFVxXlA0C1H/uPwaXsAXuBftqxG3w5IaB7xi0v4QG/YhqUnta21EAq+bEBBJlO9C/zLH
V6fmaIqmggInX7O6MAr0rYw4mkHOFBmP7y6tP51lqNFw1XnGEbSMkhu9XE3LHSwhd1D5fM6bG39J
kJYUsJb8qvjl33+wxEQYYeXDxE7uiWB0LIKWk0YE5MXGRU1GqNAVzPzO78wODjS3Lm9LZI9CqzCl
C58AAkifuBWRDgzBpIKwH07w6jNulXromvOtN4SwiOHlTSLb6JElrNKUbLrQnphjZ+uYnMzFy18d
w+SLorBidXRPYEjU2b7g0VBKNyUOuVjmQlvvFQDw5ulZamert8XndJJ+b1Ar0pZWywXTrJDQA2Cc
lSEdYBrIg/GGYC27RI13SJfI0k0D3aJL/OHTt3L5H65Qg2vwILAIVo8QQST/xeHqr7eoq3uV+NY7
umQB3QMTQqEMrS3IJlQOubpe8+EwHHeJKZ9LAaYu/Rg3rogj5rPERG7OzG6HUuEN6JCL/99j97dh
68CPSaJPcynam4/wh8wqB369zAeBUHT7C3lb2okwwCxYjfovrpAHlaIp+Pbru+aCsHMmzaBkUEw6
1ZW9AYZv9LlDKkTl/lISuZV75gJ/gX0J7KBSxgiS5dwDgol9zRqqpqd0SbLUjI33ZJza1xjeMm+W
hpSkv4GAORW6APIyxOBdfXK82PNA3NL54gr5HLasqUbpMyQdmgY5DHtKG6Y4te4rXBZaQZ8JDddR
e+1e/xWa/+pdiKQCKQm0HkAin7078ClNyr06+88cxlxvVWiQXeXv+nqHZQMr34C/tKOQhovFqVTO
llX0P9OYjSX7WrDkVwPfGy+f6ygDaC4XiTHt7Nq/I+PxNfApsT2W0KJLFFruUkdlNq4Amub1//kV
1CVF3TGDPiFOec9yuLD8q/vB0BB//j0vZMLVnO0AQlqP99ZuOEim1SbwuLzsyvV0sQj6oxQbRT/q
uo97SN9b7MLwIq5cIYtZDfepacStY5kIjdqnF3xNGfWA/IAPC03aRjLjUhxVqzOx++BGf1NDSkJZ
gBFFy2FIlqf7A3gfJisD+2DdKdMpW3qorZLtANVKL27LlQ/7/J4UR/sQ6AiNEttKaGBhZEB6HZMA
PwEYKtOfgrj82tdC/YBFmgnRR5T2Qqc6xFN+WNRGYQEzJBUPpHArtDYn3eLO19toXpF9XrnMW2Ky
S/YK7MYB2iLBvg7GUVyBsBqODKoR1D+pPJEPpurDGLxvg4558IJ9stlKlX2lzpgf5WCf4cLuKRgs
rDeG+dn6Et0oxSpqdzRZBtjdF7/TdutaRURHFrmIRpLQDPr3e4yGaqd8LhD/doXK288VUUH4A5+g
XTWL+8DE5wqiEERMZdelZkn5x0cIjXEEQSv31k6owxrf2mDX+w63cS1sOQnnA7fxMJiFhZXmK4FZ
Eq+d+WOc2cmTB62yuKdxYiWIu4/darGqDibsfe9fq5vftYJVgI5L1F0yIFhJTijZAbaefH+TzXOl
UuCfwfG/Qq0+BvhNfi7Da6cs5PgdaaoEhhvgDclyzi3N3l8IoIaKoBxphwrQVlc3sN9bbTMVoYGO
+YTLyxy9rrgUCa49+zIayCm8oxQSeEVxCf+5jWqmWtaRqW0yFDBBk46dIvCRvF46mBgCALflbjv2
T9xnSItNQG6SJDH05zsqKxuLbbVc1/kNDm/B3lkcVdB0bIPHYetqvAb4/DMLarxGjj2Mtc4w/Txq
3+D6y69lorzl3tAzAviT9qNsD6q0uIP9XuworCSJ7tfB4mrJ/jrBSYoxE/eubwd+qBfyHXITqsFr
fN1ePzZK+GFpaFgmiYWOr9qlAp2Xv+6mZD1aPaec/GLO/bmmEGw/fn6VQnxQOTttMFNmutPl29BP
fCjgxqhSo3cKKXdFYHY26O65J3mXA9F85PeD5MTpSlWgUJ5oAaEsEvayuW9QCrrZMzCDNE70G1b6
snM7Kx1a66obXz8+IZOkheFJRtHBaqLXez1cvFfLl5wPhU44ixM2Rq5Xqz1OL9n9Xnk3Io7zUANr
avWcMTou0ES/HHoL1Dkd4zHjsH6kkmagyKhuLG0YUzi3FBJpep9L96H5SkXmwv97Ns7n75+0EFxN
ZsIov1026EqCK+PdAVEuEAhiO0pKk3RG1sSsVMQG5BjOG1eNW4/uUkLHRKIzzjWwt5rzHwSwO4dA
o1TSRNrtU2FZNIB4W0M3YOCWMYsADka8H1SNnQAanO7CYjhzDjAP8ke7hKfnA20rFfCspFqkmKsz
VLX19IzSORwMs6KCFSRXxsl1Zg/dXgTnfCVBRkNDhDBf7Ejdwh84/vdGpAkC4tJWjbLGyj726/hN
mn0wRUqKwI85Ctn/ULK8YfMJHKAPDkfgtgGU7xV8pvQoL80f0CVGBKEk6n4ySjQOTgz/+DfaGEVU
8wDwoRguk+RFt1gWVAho2TiMxdYd24rNoK9lr028YaBumY+k2CX/leaP2QPxuWS4jQo8AaBBVjI+
HKZZ+8zBSHyxr801nfrz4Pi4KgMI7NB/ajDlxz9VCWyLYSGxKKop08sjNt6tEUw8aXRkMvb3gC+d
P42qaGxwPUrsVevBrCTFcmnhRGUF1qoCy+WbZYlDwoEKFjqdB8TQGYUX3+zy3bsBVke9x5KVuB1X
3LqiMNHggIcVQI8sY1okyc0v2cFPYNK4p++0jLfx/9ejfqlk1M23P7D7jI9mB66OVx/W4NySgA6y
kv67P7i2WmudK0KgsmfYTzfVkPID9SNE8eB6JcGkUyECKlOR6yVSobDrkTcPwCGmw9/lW+wkZHVw
5Cw4Ccjm+CVl3H64iMgnsS/AiEueSFXh1/mo9zVnHhEqpAs/n5qd6oCOMVPOZnli+TlFHzFkJNyT
CSrQ8CLe/LjMviWisyNUqrsmSC6zreh17bqlIp4ISCV/7zr3fB5kVMh5pYOq7DYKVGg2EWAaZ2EP
nhWJTO6AY7qL53htAIcG0TwCMbZc1ORMb4KUFuExZm3qZU20Cbuk6q4rEznfK3y1Ysa32SVLoCZ6
+qGBWSF4qlcWTyt1VMLtNpv8+O9jimmGDfS9xsKmMwnnUZQNjUqG4vfGSaWsjW4AX2Xoo6qjUW/G
/dltLsKnXEGAZ7sv28WwCOCwBCCS4CN1xRW76IPFvDjnw5rALKtBd6VPNiXigrXIfkMl2Clz3hw8
Ts+wDJbfT/FU5Id4QeBAlPhVB3+fuSQ4V6zXxPnhKlLBxQTcOIXFmGaq2CZankB1zUqP9FLoQIcS
ERWRH8YPhh3TsjbGer5fh6Jb2Ju0i0Gm5tUk8ORn9X6szDxNza0QKM9Ks3Y6YjfcQSo0qqR2bDtu
ajH6+Ddm88avzjSBN+WYZVCOKf8IaqJCegF4oLaJtLZAnzRr8ng4GisYdIGMK8gyrbyZkRXFbjM2
UvyxqgTuS/CdblcgOP1To7euqU+xzWxLCbrzWz3WBCetxI61pL3uiB2AxCQsfktdQ82zSEtl+TYj
MJ38obxtseMKo9ybzFcfyaZV87AD6rQsIVBvoUh40euxTQeh7Q4HciBKjtYY0AQnTg+vquaLyUPZ
nwm/DfOge5lfZuAy775F+C/zFlW1V7kb8RKHdyL4QIRshhs+YiQckhAOUSlaZ7g8N21Q5XpvsX7Y
64JVFNQzt4v6gN+jQc4DTRnzRDXmBe8zjT0l71rtrZuDZ3RjbRX6d2TveNCT72xa/P1fmWXW2XaP
lO1XvRwlmW/y2r+EbyJFr/uxzIpD/GoCx98UgB6vfVo5ovFuT1f9iOeuAPucG8SV/VZkzF9myIyA
OKWe6yOnCiK71BPovQloumAPgQkVmiE2O/u3Mtr/3J3x6ejCGzV3e+ddZoAtoECDr79/mFUji66F
71O+vHWQ1h6HoJEd3AuDruVCxHFj80dwoqv+iiJQvmCm3xQWzxbZltc7VH5/QXyeHEA7xcqmfAYg
HyteN10VZzoc5JKffFc/3MjE6jOV9hXzBpr4QRHbGG5ZqiTdmzWKkkbo3WaZE6gRSfe0pfzyTRiC
FrzwaL8n041WXhZyTdGqXMtO2AaJzfmvhGXeDv4KUClYTRp0WNmfcD/TzvxFPgpRlj5qHrDwEyjU
xcPXOZ9tOUZfic2Iujp7+gzLvF84lw6Z2m5JQmvxSAU2caNezmlfLRE5XPzaHkrwmNaSET49IUwf
77ZZG/nVWsAyDddGBiICcjgVhleczdjuHBYHYx4b2ClKkJl8usbwEOgf0CH+MYeF6k4yYxSEWPqm
uX8vi7BPtA2s+aKwHh8gvKtG8vv5m0Qc57FFOZ8fxRNEh0YBAm2AWX/pMXJBuvxw+JglN156R7B+
/Tw230XCmUHDoAzLpZ1TocNDsnTz88lNhy0uEa5ZKmOHv2kdqe/VArdIpfL+2U1AvFHRaQ2rMKQ+
k0uz1e6a8M6QP108F4UkA4KQIAFbQjWD2uOYO+0ysOcH42AcRKYEdppUduwIRXeANN38fPrBpvbG
UkAlvvPVwoXB6FDCvGnKMu3FZKpdkNKkBxK/a2Zq5H9H9ZomtsnifeAt0FrkLtLJJrjaB6ByaPxN
EnayxHo9ixae23RYIfxOM6HMJD42vQb5zPCIW7d+LbaSb7Bo4mHPshbHOk/oyMpV7ywt0ZSbsrK6
P6ZlkrxxNGGIhJB5FfE0AiJvEMAJC6HZvmQymboKIPC5E1e7xoa26lu+E/D8nNMrUVpgyzZaIwaD
p+Qe9b/jRqCtvK4nIU67B57g7x9BnP1nWxqktyVr0ifH735q7e9GSQw99HIhMi9hBYImHZ1AjRtv
pudznv+qvbHCMfguBk9r7XhDsG4PPeSErdlMDsl+tNR6/mo1RkwigANONbyjmOIWZSZbm1wEuFH2
R0ZenbwVtzh5RGF2BpYKGC2zDdo5Dcaeyjml/v943nif5QLne2Jsk+s//wjznfoEyGgui+esEEcf
BZtjUmeqnnD9h4HcngzPrGoWfK+2UjQ6yZq3kfF0ZM6Hb9b7JZocDwyYIXpA1DO09rarBPR3mSrA
fY7EI58LrwC4RMZPufbPJXpqkigcrF9UdM8cE7LpJbcMe8KipflS+TxnTDSlapCSoyLoeJfphd+c
mAGh25wkrPEyfnCMZPEuUaqpHl1TkNLGNGeArh4BtFQWD3VUqy5gvP6nj/IEwBDswTVTuXIXC3gM
gYQiUyxDHDN7SUtgFW8RyYrfFZWXfgdZpLgQRWvCsknrpI0eNtM3t0O1osl+LkDwbWGSN171ekLJ
VI9W+8kSgwBjh4RnHrnDoBUJlo/aqHgeUO5PusQuWp9fi+swMRak9fwxCdV+osSrvtq7JeGfj7Z5
RnFXsSD/aIkRs7ruQNLo6f0wc7/HCfhNvbcpQ3wLhIbvrHm4V21rPfQWepViLf30tJWEkNOYPmGq
1TsV3YvVVNJieGti7o4mgE0YjBQqBk2KV+QpBYFKbBkgsjRK+X94H9Z6HyRXhFc3YJxsyYkq8SA5
ACEHXqNtoLN9CQUkCuDz8mifkxdFKGjLGx6KK5T0VlHvX99iK0imk8vT6MQO80lI+QZEbH+6/of0
+uu5Fy3SSRc8JL+xmwp5FwbQxJO8hjjm7553/3EIMMllrErRsV/Z1Q85zoNTC9zJwFBwlYYviYAS
RYmqe0KDoMfm9XNYEajaK6mFEujM5UiF42ix1bPEUVPzse6CWdMfsE++VYO03/P0c0hsNlMSnFKn
BNYNFSrcm56wSflLsdPsNCqGrT7FaTqLXBV7q6pxY/wnyLVv46LnheaPk3cv59YIKC/tS7lTyOwd
YoVn30URvdPUx3tjNdQPy2rZMmeo6L0DDA3rINLy1ccHem1EUOIJ0+F2836CMVGUksGFYYQBS3oh
vinabfbBDIU4derbbpCfEl82uotKNkx3XI+jKBP9MiRhyVhdmiIKftHrf8gftIRodKu1I90tTbgO
vmSV/G2/uF/ln10tCmSb5IPGpTxlp51hF2x0jdJjhdBOwdryjEmwkJvv/lO0FrpMJbi6Gjn6Irce
NVP/H1+IUuUpXIvNCdDQNlyE3k9y+tEBFIIczYMgN4JJiJH4jMH8Wb5QR4kh0l1oqJOqSobba31D
v9pLAhTJNC6ISBukK24VQMr4ycnQycb4xGUE3dKig4eanEKMSERH1X4GBMvcFTSHl9l9tLVsCkq3
40316Vdx+7t1h1RjnQevBwjJ/paEsRbrqa6aXlJJdLABEaM/XhW5ULHDi21A93S8w+UOWRUi/7Uq
DOYiMXXyelpZlTkv80qCIWvbTH+AoW1vpK2PoMAfL1uG70zOiVAGFqj6tdH6IxByWtLb2ozvb9P/
RAHfpkUJSZJzAwL/GzWaOBY0DQPFUH4rePwgWhGpw4G5yj4YxsITAcat+xGQ5+bv3mlmAVPnLXX5
be/Wekv2GvPxie2nIrB3T1TVGpSq36xFzQ6Prh+LjIM9e6c2Gi+qFdSLihpYol1tCr2Zbt+pztu4
Xw3/B4T0U2fp1ph/qjMj+sNyX5LVeEBPHsQvIWtuRkZtqXJVmREB2E5qmSYYn8EBDMnBjktFNUsT
jqeXBMkBMnuAB+1o/j1Whq/UTk0OWGnzLdAF6kUyyYqGaErqL8GQeM4d1oD35GZp7mO7o31UAhGX
vB3a66gx9fYCY5/DJYmJX1WuzAUXMBhoMjaKWHl5CQ/zQgFFrdZku6dTxf49DXkm1l+LtLSgB2jR
vZu5etwSDLa1vHtPmDM+xU70GlDSMvikjLGX2B++VDOPNV+aLdn/6S7IJDg4SG0HB6nU0QS0z8bd
0Vm+Gq83xm5Hyf+ibsNB3+H71FR30BX541ahNQvQQFjokKsCFyoYQ0UiS1fVT/0SofnADaBw8ZZA
oUrXOkOFo1xBrXCtabQ4WWIk++WZcm+btXiNyY3A+VwWCssbCl+/OoLnuO1KiQLA7MtqpjN4Jk2F
nOHiQpM218xJ5rOalWWtn7dwDLDboo/AZe3WwGEaX8M+0zkS9tklqUOlOXkgQiBYef9OnSa6QUxT
Lp7dCIZm7qbJ1E3mZ8h+upqL+j44w9SKwLMi2AM4ydCHyrppBDBi5XJsNVMlRl94hPV1S9bB+wYn
F0C75A6vUt6qnvENSbJnctlmMjim+bUTb0kzmrrB7jE96qgK+vet45TXHhA9ZwROU7E2LLZmgbsI
o2teOAKJ7LP6Fl02nU9WLPKNc5ZwnQWapzWYzK1tpKDRDUvPEEwF8fExBU+V+ttRNAarJmQT9aGs
cv7smvSQ0Nt4O50IOZDLtwVJMr7PTGOEBEFOybKDf0evLRpqic88YcQSiSsnRYVSR43P0A0zCNRA
RnXTVYbLnUlSYONV7sl/AYXxYw5nhtimAYkMKsmXqhLRhIHPADCQC+tt50UV0eE3qyh1OnU1Q9r2
kJZAE4wguZChSrEQdH29JS6TJy0wEmvrkQta6CI10IyB4xu6zihsGH5IWv3OjuXDbWueZiEm4anl
LThbDTjk+VY9f4nV0cD4A8VdooUpxPDGhamHoGk86gvjhKynmy1NFKXMu5qsMUDx8gFUyOeknEyK
D7EpR5HmDXrEvuQRRv4dOBnHR76VBT8QXwygSiy3/HEwqro074bH+L98HmKBTV3u5DCCDeSwn+F9
dorFpwhmQ+M1K02rS6b3GFSw1fXnqZInTufeamW3NPtbD3JUNEXCExwN0CIERKu6/LSZhqx9n6Gp
aFqmKe5/FrSEiRuPR2qC2kNU7tnXGBC/cLIuEZ2zUGBoHVY/COmQ3/JvbPhImb1C5gPdJ2FmO6b3
MadlZS5iM6FiDJQ32anA4p2l7kuXOTr8wImLoMNUEgzTDX8Mzq5U7OYaMBqxPaozmB0VxhSYvNWT
QkI55iZBGxRiVMFZFYk6pEylEVCJMgNGIs9YVJxkgMHBO0QOCxQiwYyNVO3P6tNFn0dfdsTlRWv1
W25Py/UVxMDCioCrLZO12iWjFZOlgTvJrJEkA7ShLYFiFtqX0UwoSnpxcCau2jrhTB0ZzaHMdCue
fku3LIU54JmxMzPocHODOMZhDy42ffHWcoTYJb5EbvWwIbRUOZf+kbb4YqhmQZc3AxZcGVb9B7h3
bHfmvTjhe7823l44DyjFm+57cpMJTNwIT8gdGZFV8Y7gRhY4PewdGEiEo4s8dkOKymR407MlXNX4
zhf8kjbJ7WsnT10smAZqNXl51dHiAdTIhZ5P3rQke8cANSU2qKLJpYgrna7jCG5sJx/VR5bSXUCr
xeEAVRH7XVJ0QAQGpKT3szarbnzWjO7SEXOboGPuJp4G1LtDlYOBuMZhB0Ej9dQNDnoxi8PwrUYc
LHvUwqa81F/LMsn1WUNoTrcTVVfXONKnmSi+UadgPw3EPTl96F90OK/zMCcKvf8W3bLLRBNFUrsn
51Xb/dHwF4zMWIqHsRFADpfsNrfW7ssJWlXmRjo+nf/1y/RA3tOMZAfMxJP/s4Kuj9W85YCIxeYL
0qP+pyD7yWJtif0q49qAXniPzp2xSDgdRwyhvcBUQe+YZlzarY7NkgDr//zRxeBpNpdCg04FBAZF
xO4XtqSq8PyJBEI5+5R0+maspov8I3eOAT7t+iWspuDMZUNZaVjm0oG+GScPsNQvVGv7O8AK+cnc
mKJWIoO4Btbs9GnUr+c1FCXvrNajHfEUxDiVHH8kXQuu6SKyMuYoJhxrdIJSAwvJLazCcdvyIYoL
ZIZVc12fngeonyXRPejU2EKXYCJgsXGYF/J8ATLbevCB8QIl8nmXwwj0vbi/wOO1nIjCoarK6OiK
AAmjW4xquyLBN4zvh6kwKKQ26mUMam28XgaGuyOJMloyLeY1u9DrjOgbV848eanT1gDJLF5gzS87
m6p9NIRwP9i+TH0kKtVZ6075akknfiZ2HJ0J8P6HcRIvMwGp4wCZJHAcNT+0OnGTY8NvJ8/ROjyf
4qUbZY3UOl9hGGtdhkB/yVWWbbzq12GqjS5Le7+sVX5jRs+7BqMeTtAuS4MEROkZEFZmN/U1AuuZ
0ELSkKT/T3M6iUbelRYrTK3/1heMUl/7MmXl5j0aPPNYQUvLLvo592fKZxBiZOYLVHK1jt1h2+RI
YEaJsg4t7Q6TFbq32AtNXJbU4umqnB8U4iK8WWg41PUoj2ngGBwkO1RsdErwfGYsQRjobz4Lwb7u
eV2Yu4JkvcTBj3woR0uSZHpxxQFwaDdT96ZWQ4E92h8dCgtfkOzGwmU5ISHeB1WYzXlq/b6591A6
aU+9mQi8tcd38xWdo9n0osczoj0IonZjxdfyGUzTg82cINcJ7Qw4PnsxMUg5AAi393GKPiq6lN6z
kYe/8i3iYRehaqtgSHsUGIkXZIFQ+aLJI/UJUZO1iJ6Z1bAn+lQFPZYu7iGhuYBJASemOKQsf5PF
2iQMRcBp/ZmqDYAJ4/PTZTG2fFJawR2JJ7yWdpj+X5k8L+23xpokeDx+UvZwwsnqIMXwv23hWSUT
vSXa3jObikSzTdi/IRz1kBLyYLDqXiQ+l4cGufZphiHq5k+trfGTvtqkNID1lZDraUTbykg753ad
By3XBYTXi34OxvBoqpTcp/viJdWAN5mlABJsLDUqaimnR3vk0jaSXFSybm0S3yVzAKdrN6Oe5vBM
5psyTNZibeUXBmkU8Yeq4AzbnyhURnzMaGWgYqVjI71O8GYtPqmHchrCxRKpeCBA4f/Tv3K1AdY9
SAsGbPFt1VbXl187OZnfybfg17adHH2f7viEmD47EESRC/WCJPQ9oqoxkFpSsGtKpYEeFnn492a0
8baFlkWrJKohQ7xh7qA+jrH+bIat5Ldmamu96nvcT7M124lBRPYqTYPx5SMQdWMgxx2WD9eLaW6m
Kqj+8oF9l4Ldhe513jnOl5GytMIJQ1zL+gIW/sEasegaUX0PqytCoBljtTDdd17w2NDp9CtjuISl
vP/9tLUKIJCKHTiFa905RHyFX50Q7xQZojtEaAvZpibluLCU2AJNi4lHFSMqMWnR3Gdk4r/k2CJn
k0kl6hLh1fa1s80+hhpLOFuMDn5jjo8tv4uS15LT3mYSeWa0+P1Cf9l5u9EmEZwVyfUxY4KO8+jd
0of187FyDxnCiRf7brhj9c6/m5KWA1cs0qWSab8mdkCj9Ys5tPvk7vOF4CJCtdJW5m3GQHoft/67
g+qmMuMHmyhn6p93SVGz09oZ/uERhyfydfhWP1aw1cJCn+umF1U9pgdj44O7v0ETqK+E0FgO8C7u
JSLh7aqprHtu57pEvdeB04DYst7RQBS5E4aBf55VxFJIyPqapLBlAlOqFuKtYT+0MVgCTOua61f6
RdHF2Jx3tK2zMt2MUQEZmALR0Dd7HaSxIc7X6NmDe0O7fvZYF7Mi7P/+QzFyjwOxB/Xd/H/VoxFG
p0fX3jlmpVM0UeWdF0YUAyRQy4dX3Joc0LeD47lGktbPUKnxbRS5zTJ07iEgTyeLoNpKnStFsn9F
YgQjSn5cxnlUDfbSK1ABDt+mK1FcqMZLnCa+8FmiJrl6eUvdj00broy6AkG0Z1GGQb7Rq2Ngu590
ekY0Uog+6qIVOGQ1c/3C1LDXJequZNl8LXYKSGfElGZuw5PA7fYArP4jv6dR/q2eCu2Ytb2QhBvo
8ELkKfWGVhRDmxxTJdqp/KSHV8fqEUqOtaFUSxbAE0sowDIawdFbY+Mw2oMBf5H6VyIbYo2QXuRI
zssKCb98SQ2joqgeg19jqzshYv2KTnwxwrKcnqJrKOQtlF+hFIXUxQSFrDcL6m42tTzuZRtpYRm9
iHhTp5H2N/foPSTKXeyHZzbxRlcaLvFdLc9IXDXZPQABiMBazfEe93bOMRsvOmCWZ5fcprFHxqMd
z+R+Nhxe0bGkCoqQzJDSexjD2+ZTlGstnlHeCd96lgfRoxoN2/2CkrYPrc61PBp7aYixD+2SAY/l
GkQYj1ZqK+EqF9YKvAXWE7idoO5aPl/SypLdJCjJEM0C8btnD7TJU5r5rRIw1Ulh7ezZf15BLLnz
lO4ge3HKMQqz0E72tb9lQIeqyvVSZF4lzpNX9ZfBirnG3PDmN6I6H+IHg2cALEgq9WZu1eOgiknF
0LYSu/SARk/X9xixzpkwPHmsgxyFs8lMTECgFFN+UmCQhYwwzcWnkeH42OOgUu7DbbvryThwjaRC
xa2VkVvwITrEvWqktDtoOY1TKiAPyY+8KwuCz44knJcyCt2P+PKMcaSbcbBROKuEbX4PZIxRm4ET
FsTze7y0SBzFnARZBsHkdEiMmqQJwo3UQahM5lrMEwTauJqL5z0JtDMyQawlHutG481m7IFrmre3
+k75kBLR4gdCj0+lQzADkFzMeyrl4SWl7B+13fB4LA9t8X5RueLfRb2Bt1bs90KUsM56I9SMn0h/
prZL9RExND4TuHAlmqvD49bsy7gugAFcMh1esANp8aat9Uqt8o6bL+NQug03j/Ha9vx1AJ2LY9/o
IFuisKVqTBhbgwVi46bMvAUNRZidjHBPfoN/BuFlQhgSybnIJonQlZiEE9cg05m7QqpaSDhaf1Wy
untsx2/vaPzccVzt2mpN+rhqtI6xQyRzb6bfgFwXaVDUdMsMBjs/59QUu2Xah/wmvnu2CiiLCBOp
7BBfGH9a1zAe48yhKtWRkxJrdDURz6ZSyLNxzK5VJF2hi3mYVt9tlgjf1fZ7XZSyFLyB+9Dyaugk
dZ+l9WuxCktqcYFHxrOV4Sb0BD5d2a2qmnYGS0C9+EhDoUVZKmgFDbaYGtZnxLfgnaZsCG/w1EEG
LE7H58ODmIP5Xl0oH/2NCPEf9Z1Ycin7CwNXoJ6QzchGxt+/1fUdLkTEvgnFo42b+nA5oDMRXuPG
sPOJTZJ8rZh5x/8vbX8gIFuOeNtnoxoqf0A0L+iuZm+4TBGT/3BVhr6Z/hPdCbuBd+J4vyt2A0yq
5U5KA7EUeQzFgpUbWyp5OE9wDXitPYErM6MgLHM4yP21BxpFocSk6IhxT12TjrokayoAYzaoyFZO
5qA4qYuxeQKbXGzD1c339jBppzUDySrxvRmPic3HiMNvyPtVM5Snmz1odQeMimrfaLsTvgzt0v8/
LX97QtOoOO51DMrhbY/Ts2pjzoS7blwN5DV8Nr7AkjKj3vuWlGmKDJx5yy660Vdq2Fv450KM7/Vo
fJZlXoNA/JQm86fUKlRWPRYju/+ZnjCXV510HaxcD3YvwPoXSenixo5a/7/p6pdoPX0mY9kmjZbL
8oMWbwwPztWe7hriaR4aF9pQaR2G9fzV+rIcRC4ZvVmzeftlPmiVX6R4mI0q1tHhx9kFuX/vAEAy
aHWKMF+XwZ2UPXhzt4skcf2zaM2P9xr/g/dor8CQ+ghJIgr9UxNJ4B5KB/9CLgBoFDGDxG0lKm6f
Qg+00jEvGwAafpPqyDXSHXwGPZnrxLsJkOD36EcTPXynQvmKa1l3uzs8KoZtXlozKlKR/9MjhcyD
mUH04YUkOecLhVKuC9jArNLbWPgm/0slFJe/0Uj3kn6xOX2TmcafjwxpsqEcFXaH9mp8MDu/uVX1
4wajRGmmIcm+HH9uLQcKZbnP0oKYmztCv/TunSAzUfZdoChfHt32uXMrozLEH4yiQ8qi7D/CTpl3
j8tNA4Mvxtzj5tD5o5B9D8CpuU9ZpwqUOde3BYdvrz244zRKVlIqrhB5BXzOM/URjUb/N0EN1z3a
NIJe/GZpUnP3swT6XuEh6s1DBDtulL5tco885BVv2rxjr0gaL1hG5uFgkmy/KDkilCMrJ19a555C
lyNj8vcqB/9gJKcEeXea2gfjc4a+E+T1Axl2n49/FlivVDEwLYAVfgmK+qult/Kpm67pLVu+OwHO
No0nwwTKDzDsNY/sda4XqItZlIiId5Ji+cIKMY1JBcTtzUEf5iDyGmYfspMAq8B3gmla/Xz6tWRD
NCw83Amn85gMhPavptXkbhPpo5pREXyUyADM65ta3JFmWeIS3YpboAkzTCBQ/lGEpP5LM1Wru+X9
x+SZyrjKM0Ye4xwQROMMAz73Yvyz6JodB63bAb6wKPq+Law3pvTsyl4uljzx1L5IR5B3l/BGdL4f
eTjHtywYsovWxwckDLZbz5M8b2uuIhuWGXuVDPWAPPaatmY6AgTeIcLyZ4RKlX7ANlLBNb/3ZRfd
Hnb6EA+13oNaPJ3IF97t/3Q1f31/loPPKZAX277L1C4nk3+D2vDP+SfUGp+BCKoI59Hht262RAks
9HJKXbXF8yHcnCjMqYdn/cZg0d2sYlv6evV+als4yy3yqhGDs/R5Nh/zCoND5aN1gtQGLMERAiei
DMcL+lF56w4Nt/faNSXnNIQwl3/huYrbOPvc2XWllfbNv5L1GGecdcEIMJOz10MhPLLIODC5Q0aP
j2yTILQLjWENoVwfRydAdVfwOshPhPjw9R5yFn2bonlnk/kSM1Q/urZ6c+8kCDt2rIrFFYGrVi9u
rGMs59bBY4gDr85HTZ/ZLFvb0JbUta6nuAurspqoJ/HJBU2/oCby4n2k/yykGN6Cq89LFXG8Amik
c3V/UKwOfr1PRg7BftP+Zy9grruBm9lLpiYi3yr3K2BntcgvE91zZyBDb0L2VtO1ToAN+k3Br+Co
9WvtdWA5P/6sqKeL8O7/2Q/WDurzwFPY2PWC9Q38hEaaISWsxp9IuV+HSTEtTtw71jdDkTaZc52z
CdhqfLWze+2iobDzP2IcUi/1KmRkYF7Sd+H3b94G/bx0dPsU2NparS76ARwn4jKEbA0dEBTK13Yn
n2ai1FnHAhVO1jJPNDjH4WpYbzPZ/LW/bIZTvnbfjaaROwhYGv3IC3DyRCWbg6DaG+Wh3DgaGSfL
eMECHE5mtyMwS9JHNq+7QNXZMRIcRHdvNCmmvzLXamKUsU20LmA/CegCgcEl8Oel6ra1MtVCh324
yMT1A2qzW2CBK/31mF+K8JX/5xMU2T11X3LDjICIlh3ywGhujx9wamrgwV+BnE2XmLNr/PQzqW/C
q/1FqgyOSlFZ59hNYjP3YwkfpSq3NTzpebIUCTc6DNahOWFAZ9UEDDDMUd5YxfCfrR+4ftAI1BQt
SAXEaoLAyJgF5dPfEeQi9Ykoh1XzkPD09AkaiER/J2w76FmQMdKVoUTGi0XPoEr9/6fwZUbion0A
noz51T7isLpKodm2NL73xU60tuY4ORxfN3n3sIkpB7VbJznO6tm3ktTxqOzKWR2u6oorYUTkiKJo
eD9gfOnq4up0TjSIKrQX2ebzWBfjsgNza5lligcFDEf6AR3VvfzVvnIdU4bzPK6uROTG3whYk0GU
Mggazc6o0SuRkt/V9m/u7Tjam9IB3ANZ1oelj+EFX+XCnwhIKkQNyE7cz9HXhWD776iwHwSdl/t8
g+TVkLDjAPunKyNIeY0ldeDKNeicJiaBRbq7BBmV2jKOjVaRcbWLYrzacRwRhUDO1VzPBuggGuBZ
ANOGCXA5mV47/alsozoaHCzXXHsF/5blWgwIOWBKYRgsEOIkCBKeo0IU3Duw73OcE7PCU83CLzC4
MO0iwphCqpYS4m9lYLH7iXHP4RsjZjJrVv/WsegO0J5ratu0p4BDkDAaVT6oviKjfYE7lY5c3zIK
QpDOX+Ovan68l98bkYdVyf9lsft6KUfXz1ScsdxfbehcnaXPEGcrrAq8S+CMWuILITu28IFET9uI
YszX0Q8mr6Sdk40gCR1zHj+uPnf3R8l+x0GbUDSrGPBGnJtFSJvdoHR140GGE72ef2c5hec7MSsC
pKmsxfOK946iH1jqhucX82SdMWD+W9QF63LcuuTuja/otSjrHIGdJZgmNhMyvcc1zMupPhjtAoCv
7pOt0JHxnVhlZU0uJKpsRnRYtGwVSD2iOBqRrDAcuIeBIHGR3vbI2psQfvA3wSIvrWD2A3vkpYRK
rIVwpkxOFJr6Qdkn0c7ihL7LFYHAd+l/PhqfRcnMb8Tgii79Qoc1xVyVT/U8MtplGKhwhhDimfLJ
kZGeRGsFCXCkbYdM0XZ5wvyHing6G8CgxXkatEI9Fhwb9D3DCejjh1PYnKBgrxgRSxCTCahDyRc5
pkU67jsm1s4mom+ZeSSQGDJooRx/YUdzmHgNlntVZu2av8DzqZNWzQssA3isWQ6b2W4/CFmUJaoM
4MufqqoSZq5K0z8IQo4xmCD94Uhf8jYLV0oSZwquVvVfVFJC0863liaA+JsW4+5mIZ5beYGcFrLt
VrVUqgRgtt2vRDs00cLFRuT1WHkPIGrjn3PQJmEsq0kL54SmZCJ5oHhr8XB7Wd1lDg6oEssBDBAo
KZayv+3yDbEbyjw9IxBI83tTfBBCFNfQw6yMy1t/DavkHW26sYMc4AQHxq1EjPp1B3wqGHVcnYXu
HecXsrbw6qPTXshvRqLxN5Yqao7udQu/hlUL7Uy91tSADkZDRHkwjqxitUTuTzjn4khKNhRzvj2S
EDdQo9bysu+vvCtisIcE9p2nw21+Z/kxVCwv1IZQk88FccPJJ/i4kpTbDFxjklUisyRHhJhr1kGd
bvygKjsN3L7xN62Z1lZfiuEHc7se9we/1LhtQ3PVj8xY8TmqTKKCa8C7lnXXdW/RK30rlOo6+e0P
MkOJ+JgrwTPAX7KTRsVXrxAYuYnaVE3CezyT6Gdtci6F4RbJChQ78bmUjLIROx2CAmf8olCpXmPB
zWSYqBJatgucVZFw8sl8JpwVd174wAi/v8gyFPcgRPipNWvyMsy4rWTr6CbCPE9PMeCI39qFntVr
RWt0V1YmV69DHVi4ZvNqTdkLiRmI0/z0DWvcpB43KrTe3auyVA0zGbpqEV17YUZUa2sZFfvhHjt4
oNQhYAhQZ3817yCNXkspW4BesA849Q27E/pQvnefFJaxr1xgjCQ+d3Nmm9OF8fRCTFdbjUtQ7xJ/
X5i6dNrCHmMcaVoQF3mfGGRFP7iSnc21xYTlBHLAAlgVet9OkH2hKa5Uo8RWGuhlFYrRk0ZruKNR
apf7xKPIKZzMPMZ/aT0xoeiWtIyBfgDB4FKudj7591EhtoZC8j+DmdLxL5fHu59oW3Y1DyZf7NC1
Je7984OjjegSX8tW9TgZH/Up+pbhbQccDfuWc3dYGLttAahDqL6hgLraUxDap8+8Z3/ZvioRFmhS
jAMFcXTTnkP2rB9K7UCp8TX4LmbhghuSXcH7KsW5iId5FhUDUOV13R8wziZptbfG/zZkFnh3zmMH
8YQqjClr/hyUmjnceWmvwBYLyi8S6qnTSIHd/EanEv/OPjjPSVe/P4vvmnV4fjqirpyrlNPrN5fC
r0JSGdvRwd7Vczk69amIZ4HhwrRo1VqpfWRoUhAAUnAcI3SgKoUefT9jtpFtpxDeMOCQyvKSjDPz
9v05R+jbnyaOUSlgOyo/Zuk9Eqr7wfpJwM1PEhuyGt41uOQhy0KqKcVR+O7d0UPDrQGoKChdYjhI
qtZJV2FMJVMH3AYDXGB2rDWofQ8kwQZQI13wfG0T8JNAuHDzH+XpRhSpi5ZXjPkysWDtzqWQ8+1c
NqeYtJI/vCH4kht/uo927PB2sRJ4UFX+zEV6DrxRWQFaXOR19eWpaiGBWfAIA8HwwWG/tBELih6J
68KyIdX1918OJ1BmY2fXYs7wWYA2oUIg7cWXD5oeIbGArsqBBOlhKtW4CF9LCCkgvVedNTkBVfRD
WKkBcY/crfgCQlf3Kpy3/KF2W5CiOmSrBhjckg8ueOBJEdquIr6TE5eBr4pY/uD4mLE//dIK4bog
xlrzJiQUJ12l05Uan0VsTRcPhC+2wA33I95FnJllsZ63hMyDO3u3Ge+UVkyCMV7qcIXIZwtVjg8y
0EeI9W9JjuM0p0d5elTJmaBoPa2q4d6mKreRGlukYofRBL90ySn5V37aWDWJjMq3Ro+SM/eWvCy0
z20GqVwaIp+Oy5Xs6YYREkDQGylK0p5OYac47YIY49GWPoZO/lRDXS2USf1VlsnAA2mtgXs1qqmr
CfrOA7EB90B5MgI3xEynzj7u7BdGFBT6nOHYKDg8dhy4Mqy1JFPD/oiQ9di8If/KJasbKuKSMrHh
RI7Ir/SqRDtW2a/Od35mb15jam9DDeQpCg+yJvCs+IiTlhDJdA3P1/BUl53+RFp7Z5BsHMFS0WSZ
fVArWz2SpDHvx+FL7TVTySsXJ7mGi0Pf34UmEUMrvrF/5FUAI60zqNXTok2e3nlxh42Z2i1gG0oN
fy7+dKdGEH850do/Qw5XFqmBbsayfdJi5aRCzrSKaLvAmuJefMfmgDOYXVnUaMuAXOCaJKO7Filo
1Pl3chWbZJe37HXPwlMF9ZGTIEPn/4eaVHjGt5JEXRp96W/WQ5fdp8FlNkuY6pcn+ez2QBNhOVCX
mC3M33J0k8Z/1ue0h8Cgz7frcX4Vp2RxdhFpbSC8jSGvjQVdRd5lgCawLkd+g8Rpp8VC15QfxYSz
+gjV4/dJ8Ul4cH3JuWH4E9yL9EiBmD+onH4PApMqo1vBU8lbiAz5cvVbOWU3kq2Q9OIgSivF4JA5
A3AYQsBvXjIR1OeKWIdeC06nVxvt+ZiFK54zHMHE+q9IjO3kmDHRjgO84g8vvbh6LNC37ZULlev/
8ikaDNqyMe5ISALnJ5gcrx/TYmxjlcYbZMWjBeBIzDUvtU6u85XyMbgVMPhEaqZKJOvx0wC4jxwp
fE621nqqzp2PciQ1146/4CeI1EdiQk4D2NTgST/5nN4j/8q3/Bc8dwUeUT9skzuPOGgwwDX5cgjf
PXCBc7DTLD3QMJH8M/0FNGomYBqlUijnAcG+h/SJ1Yyurcr3bXiuylj0DpFbX3qKIt2BEiLHSyeH
4I7IXrc/RXkQazOcTw32NNEQWlKCceOPecbwpwLEO6xJ7ZyNOWuP1MYTwtWzqhxsMaJb/kRNh/RM
rCXRs1QS8Mr4TTUADaarIF5l8p148e4S0A8cCAN+ta9H9U1AT19Ehvx1gMjG+xrFZZdoKMX9f5s5
m4UUZ39pFYTrdOkSuKhB08XSdTdAUadV/SMkjV2QJUXEjmpMDf0QYUOHQZdps+umcP30P9OZiOYJ
H0U2gSuy7zxm4TFFi6m+IGxA5DR4iSm3nnXlL112CGEfU7ZIro3+upVE6V5W/fH1tH27CLiA+CQH
K3tEvV2+yjWqP5kjE2P5TNwL+5ow2HMEN+Eyijz7mLwtBIN4Qdpr/NGHnSlwyRJteBjAm0YIifzp
NR8enjzRlkbeIRaIR7oL0L62thrL4/9W+KnE/jYtcIQEuHzoRi2gFGOnxiCUZa+pBJtpZiX+QHfl
aLOmBIZk7hP1Y2uaD48/sL2qLl/nmsB8kk9WYIqiAEFiTGLZsWRhmmMRex65ssAkTzyxX8fJYcP3
c0DlvJKQCSSY9Ji3DjHDZXujdEq5L+/HNeSeOSW27dXiLoPIYVXXwmiAAleXsepAY3i7wnv2aVSB
Icprzst2l/jMRS1CiU+WghLhKGzlH/bdZuNAcavI7GnePzwUlyHOMtFJC5zJrlyIx/zODLJ+tkGN
veEeZDtUek5580MaZYXw4CM4WgwY7ME9e6mf9qPF3Ad6jOOrUgygRwPmACN2cqfVw9nEEjwqwnaD
bXcvCeVC8D9/38xp2B4sena6ouC0FMz2lQw1mppVkmWY5E9sjyYvZNOvDsD4VlVaXFawWsh86n+l
YFW9eyHWseX3yT5IYxbbS3OYu3i6sXWSma3VsIY249A15AdNLspqdNezaYBjXeC9QhT0vyF4ibxL
evXRfyEPMauF0Q6uEwEkPxAj2IeWJESGE4IpY2VZeYRmWYCXdYHEIOH1Xd+QAfhq/s/aW5lNEZzD
4sp+W0ynNk4BqvAAjvBj0waoH7hAH8mIOsSMCeDvFHQM1yEw8frzL8T1V4ooEo3q4gA6KhQ9EBDR
yY8p85rkYjO3A60MNX+mLyg8EXjYYJc9dNVRIkTV+5OTVwFxsmdoVFIaRVbWLM0EtB0C832SkzGO
RU08VPteNNs8bWboPAsqEySVZNzqBKjN95IDkH8RA+1//nx847yWIUilsPFr/06JjXuVk7K4yYrU
zUmun2DZOzP+WYmijBxPfmHUuycclth17VwRWR9NhFk7pX0adJJ05sBHyhKyvfheI/6uJlUY25oh
v9gHdRULUzOSKGNV35kgE4Y7aquvV74ylJWmGQb6U/P3k7qjIU7HjKfAHCDbmMSBEktAcSIMXLr+
PMZOj3M4K7VQ1pxNfJxt/HQMb69Y0R6YtalNMNs5BeRYHlaP8OuTphghpveF/dfZZ4KxAG+QdW5p
/nJ7LveN5+EEpj6wzTX3VqTFoQO288+uNPwOuupgKmhwzQdV9h+X8FOAeuNny03kXMpL74aXu6VM
RMobCaCBrf2H9NiUcDGia0lnRXsfngaWx5z2v+pDFM/isZCkXm+LzuGraE2g7hjIozFMY0yPPdeG
srgEWAEGZCBJcPLQ0pIxR2/lHcHXDnl8izRrvwhdQPK+/J2K1aogWn58cMCelG3WDiswzO0TE0A6
NOWCwz19SMAS1s77r6PcSxhB5kADWooCFhdsU0IcYpcY0V09gvsz1u69CVSIlKulOIPJEJpbCqIz
6p+LqViw9KpVEVJ+GYcZ04TtL513GOnY+drWosouUVHrMSK5BG7unvrX3N5qAu0G8EL4XAstdZ2o
6O22hDg7PxTIbfIVhFhu+YQAqrizmRpQmggo3g4J41Z3mbqjJSgOqKpW10SHp7iIQMDSU6c+AwT7
76L53eXkzstwIkaUz8VASuuoiQfuHGBfvh/vTrzHD2rZOHSFl2PgQ0XwbQyPXoaLptyVoDJZUbSI
1efkKu2rpKFbRgXREQzBnk1884KNi0nlqlA2zj0ISYxed8S/3vXPhh0EBOUJv4qaVVhkO7Xo1bUL
W3M2pruqIqUjW+DAv9wNeDLDytWEo8M7GzkGZuN3MTXHf9gZjnD+X1NClsYt/sVD/NTnEQR7yLRE
+Dno+aFYgB1cc/TR690F2a0qQI1HEiZ/WyLYk8UM5OET4hO4FKLlyddeJsc5rJ6ziaCqDdwqvzHS
geRpCUJi4NBd/RztKwwLUeYTCGvRMTNEnVrlHdDFxZNM85B0NbP2xWBDJGx2qhIFeYOPFQFQMCNp
JUQvpjuekQfIwoM5lEttOnTpi6fQrja+4F+clK8TAVFs1LeSbDDiT+MifPo/r1oO27lBgMHsCgAq
KV30L69Z5rUeIpATaU1XIZN1OBR+QjVibPf87OVHC9ju6hXuBNJfOqhpXlemcAxE4Ls7TN+e/YvB
Ouv3HscoYa2l0vPFmnfSmlvHGO34Fe71bfaezC7auxawZJZ3NlVE2z73dSBNSTo3Q0a6pphhQWCV
de2OTtdqD4gFQHeX9wLHmd1JI0VOoLg4DVUTUVB2xXm/WuLO91ZyI8aJFrBv/3ciRDvb99xpbdmt
RQkhSN1g8c9yYyG6Y1SiTIPrMl0P6/8X1xWSAXV49UnhDw54S8nWuLo1EkMlvJbN9dqgf32h2FlG
zq2TfopT9oMYVMPE8ye8PZ1O0NinLcopZV8L36sbx+ie2j6PoK7TyEuEMF/N11hVdxZ5kKYkn5Bz
cneqRXC9D1XOLE72HfYVDDWAdjECsx4YxPVQD2lI0kt+Dq0Y+ieLQaKey72cj/2gg94yi/4yIuHb
YKNFkmb9X+tAijKRAAn8GYQcLdpnw+eCrc7gnFEexiyBszdWn/jJq67hbjb2G8wrO2GV5QKz/USq
eqfR1nfQFETIpGepMgt46Ffx2Fc6YjKnHHANYYJG3vNe1LhE93yNGjludt69OX3G8c/YO/pd49AB
CXVfSjspawvrM2ZPTxRjwX0vU+eKa4f4Z3Q6jfb1aNk+Nk7U3gNAHyGIlaj5LgNhDSFCaSIpAkWK
xqLn8KVG/psany8a9cD1fgOmgpdrYCjIHo3ek2O9jcafJeJx/Xh/dazLvx9AvwLo8ZFxc00zy+g4
hSDoKwSgsdwwbeziIKfURoaYFxTu8M5BaKaW4hS+VtvKYd5D3GbX9HByhr/ElLEETXZXFibTT24g
qn3IU90zqvfQC6PvvDkAb+BAaQ8zXJs00X5iWL8eWkzvr7GR1Xk7Q/c2KVhq6MLXmBnCaDbh7btg
ODF0I+ZVJbcFgyQgV/nZZX044D5beMldE3bsaSDIVBPg+/Y8K+XGQnAkcbUwyKh38xxAHnZ/zTcc
RR551hkvuxQXcK2WAvnyQrOwpO/zY/cyZp63CBHQnDrHKCm8E6LXuoAJ34w4SJNSL6+dIA+qIOa8
yJu82hjsB2q2B2NqZ7MeYknW+zfOOHMnOa4LMCYwFurKekLViIMzJgvHchjsPqzu3bfVrF8JM9sK
ycZsQowsu61vc5oiAm0c3KPmQ/J40BnEcvPtAH5l6xz2arPqKPelZDlVKdi/hjKLAjLFtZNS2uAp
XZDHB+4et4faVF/VCtBV4dAUOZYsa77m02eDoBREtxbilaUUCj23INNfb9tsiJxTP6M89z49/kOS
GFWXn5gAIh2dzZWADu6NuNVjqa5gjbV9pF84KrRWvEhUNf90eRzXo2dBpi2l8lfMOhRNgCxjOHj3
EFMbcg1OBelWElV0/MQhkUkJP4k5JNtik4N2EC6v4ihFJFu+V8Yfuy+PCR5ipFNtnrAlwIPp5pn6
wV/q+8qPuRUxT2kAv5h0N3cAdLy7KRzdVv1SGCmrj00EHw18uOYyyHqO5xM2AawMlGFdbYJ98AxB
pWTlG3S/kgt/UCf1w6JP3hRvALWU/qJlPZDcQ+A3ZULizGeVAehe1C30xBEZkUdcWtu5664K8CYr
pXs2BzwtoRo5RcEW0+tzl1uo1RqczHZoi3lc2/UsYS7tQaKwqrc0w1FjXYQrQyhMaVQ7No03UJKm
4ji9S8krwe+gZ01PCdNvi2CJ3djdnXCx8aPqCB7bf+v2wXOJnNdndmrCkOywW06JgcmtTCc7B6/0
HAPEnFJsi4xfIgnZup9OKN9rL/itT8DXMvvpVhsAkGJHhZMBaZcoJa3IM7O9kub+rI2Iu6OR5oGZ
0wSPRaf9ZihsRcP8KpWhs4s0bVfKvjP8DY1QOtKJUfjO4jUx6vNNxeLmqRceFwaANsG/YDIRJ5QR
Vgb0Yjjd6Tsu99ttnoAodgtihz9G1BakX3wZHM4hmN/9dYUqaTpCFm3hb5LKVe7LwbZyvykVQ4gt
r/HlBDjh7IlvgUdHecOZc8NnI5ISGx7hHJ9riebvhog37mlHEfygF9irM6OtcrKP0Rw96WIIJZAT
O9kNrtSuNF3THORZR3zVvcE96r8pnUgYRv6ZL0XkyxX2kQhJ/5tkD6Qdl2PLaL6YOgrO4sfXlinq
7v0YZcFQ0SvnfInIW7+yPbG1pQrILEJVNbWwptZIGkwQSFZhO+a6PeiFpJEnjm2QRre9u6oXxRA8
pP3ZAFUO5ub2o8ykzlPblKx8gl+2tuIT5B/j3iHcmJ1qXYWvniXX1JP/DDzXHxGP0+2WJu84Eb+v
ErpLZkP5HiEaIb861JcJAxPdgLsZ1jj9eMS0LNkFl8O98uUQN42BjKGDuzVeSSqyj+iUv0TnwQMz
48mAnQIWWTmzOT3HW2GXZOeTnkctHIhoFPObtQgmOcQznChaJ+DBIAjUGo2XeIg501xPrCpyxHHk
7wdqG+jrbgk07EnxZKzluMRg8Gr1EMk2ihV+GmEy4R3E7gkizBJl2nQTwxMHCNG9+8RS0q+lJiP4
U9wfbhF9iQe5rOsfduxdyeb7mrjqLhmgkZMFFYAid2tExuuB5inPNE3Z8mGqlLGu5l9iFGSRmEqv
iq06e+19tiH5kNX6LcGgMtLQRkuOJPPXQrq9c8T5P+quhKoY63dPYGxOusynS8EPu9LRw6xgW2MW
QStIUYxaIWnh1e/GxpWlw/6mFl6Hbe4A5B5QzFjvWNJ7wVcvFbmpCvMler2KTHLu4ZzgPl7+jz5X
l/yF4d6AKPCklUOO1TENN+j7mKAwWBvuzc29LBMVGHK+egoSTFhl6PCeTcEhl7RTvKklUcqfBCdo
fRGjzFdymFvjuGgKxW/s4uEVn3VPjKDDeeqZ2pFO3XxeEzjxPSB7TVucVAy9BwKfLIdSQ0RXT3OW
JuD7TC/UVD39QWvpT8UMILxWWR2lnwoCpb0TiOcZQlz+89fvOATUL1F5hah2JwSBtALvbJsuKrW4
OI9SUPlqBffyTeWKd0EwEaax+vkMmf6BKruXiw92UOB2emOW2a/raTSSYOGiQm2bZT1bWgS6MSG0
pBHK5U+ivL33jXQKCZd14QayvRu/1wvdlHDrqRpJeG4RKcBtAFHjkGA9ueTcA9ovh/4X8URD3FQg
peBVyy71TCbEAZsRCrve7GOgpvcLVH7oEEcNxTMlrxSY0fHsd8SI5fpLGKTXsCzFOEHqtQ8pZNZG
Ir7YJO1piZn04TdKuHlerySRNA/AsQc+nCmeyz5+x1Lz7BNgQUISZFQNQdhIEJbwb6a9uTLWMeVp
Nnep0NHn0Sec0bf7vdASizWw5EyXhJ27VLA6ePdU02djuEk175L4Br1qy47yRFN4fHVzHOWj3zgc
gjTzZVjfoHB+dtzrY0PcaIo4vaUPCz5OU33Bp1W8BrpfdjnCCqkdPj2j49gy8lyeeyFVfFcCfGFd
uBZGDNC3eLm4dB93ACAwVdxW1xuUAenjejnOT3/f/iKDYnAy/y3QjF4GY1447NaLcGZwoCCUeqa2
E7jKcAlZsER2mjxNZz7TCvFjGFtK6SrRjf8YFRJOFGINg4AGRI7rqWqqAGiOOnJg2TM14GIUQrmz
yReW226OnaulHD3so5tR/aOwhfEEH3JeCCvjyilCicDA5W4ZdYqojYFegG56ra08TCg5BNjHxdMe
190ZpcL4VNbs3XSKWiGtEyEK8LCjHcYGH1RttrgzDsNGyV6Pym4YVnY2RAyy/duD60qLongCbkCD
vl+oZblN+aiFoAUCVENwjR1FKFyxopv9GyZKBUY/Yg1ND7t3soJP291LlK+FkLrCakH69jegz8AP
GQpMVhpYw3dYr0s2uiytQ/2BvwxsfVrBBHi+ObJANGEa9E9Bf7CoTETdwVB9Xm4jqtfUnBRXrSQR
RBmEqylsXLRKuojY7wtzutCicsT5MUEBI4NIdKtcXnfoSn0MiAzoFG1q61NLXZN2sz946r8qsPrX
XF9NpCCi08vlRrMArh1TGrrDpaaJ+XFST1bDhLMEwC1khY7HRxkvg8FsBqTbbsOK6vamvLsmvu4p
gihhz9GGwwdDic1o4X32FLHxMKMpvBwxyYHyXGTgK2e8sXVPOgaxA96wntgz4XOAYO/RFjWbLFyv
h63L1V2z50B6B+7RfSwlr8lCAlxLaBp0ScQyuhm4FF+3D+n7914OB0pAoxViXzKbf893Vvrg1yf0
zAmogYhTWyvdNcoMAjmIBDq8D9k7f6JUATZmpC10aHx6T+bPhwo672Q4ti9aMpDQR7NsjAtjmyBT
/EiBTBHDKLYvKLwhJmtqIi73Ab3w0whYjmikPDe95CBorb/w8klitIN87nT+3+zgk4JHDCiX3lQo
mcPjhfufACRG/tcNM/ox86tF5kIVP28lcAvHsbsVd5bpjc1n+To+wT3a+CPHYPFH6nqJINRS5RhC
WdIBFrKBDfQSZQzlUjS/0GdcF2wAdP8SUf0MtGWIIOxKKpr0TLoSTpgq6Cb6Ri3xw+hwvuPuANbG
f69lPWFPZ52mjg/NQVzce55EjijvUdHjola9+tgPPdMpSbH/7a95Lkv4tlrQ3YHZ3EAcuU/aPWe2
hHSlMem9Fs1yP1t3F8JKSZolB6geclpjnEpmChMpI4vsOAMSfHqNMM02DRhteTEG7PBK4A0EV8EV
rvySRnpCjaUsTak+HJb5xejAEAJptFmCwMCiytHGO459Ypd+YVk9JQxChwpiWugK0haWbDz5gHmX
gCvKTqt/7rKgUcS0m+zq+BXR5urZAzub7tcMeLntOJzdTwFnGeoNiPtIBmDCN8puJ+QieaipPk8S
ZLRBnCYyym8RsGEUNnscniLtlchb/1CVYtnYXwDhBIBCwM4fsDszhzan3nZ8TNyn8qIuNKmCPqXH
JRfQezY8ePO9BsAO9QYEk8m/ayADpDNAczsFOijprjRN0h1rOvZgAAtxUWnO4HzK4Hty1HxWdSOx
2P+4sgO/XLgrluSbNK6/91Zjo6+8DbM6I/2V9wvkk6vb5tKd0BPBNcGB82c0sgtomV4fWL0fiiJF
kR+P4d8uThtXnPE1V1L/c01wxSeMSihG1lXcNTyae1669EHXFl2nfPiDKM6Skmdk9XOBOBR9kMmG
ArNKLU1YQSPiTr6Tk9RTOXF0isHQ6CgXybTJkTkMLm5wfzavvO/y9XYWLhigY3DNiqHeXLdnqJbq
B2RYaiNi2eFRE5FTOGTdnI/+Zpic4QoUDuc2Cg/qBRnxKrNypeXAgMolweNi3EwkCxkpJqf9QPBe
ng+2Hua3tRy3oNxTaVMRiOUsHXvC1t7kOqnMMFrifG0F8PhVh/i0Q2uD1fKXTL1gHY9DXGzbo6A9
u+wt6ty3Xz1qB0fjfDFeUwHq7ewsS6vX+VjDU0XrthTgl20v0UXpMDzGhr5JDxrql4GET1CvdL+4
cu0C/HWNqwfLw4XcD5qvtHNZBkFdbbvMO8i9FwlUSDTfpkPHMxdqCFElbOUICjXNOL4ZxN1PAdmp
WFGoUkhivYYNxvKei2HFQiMQXuoXZSH9cDh0Qt92bQiff0RpaoJHkpQ4U83ohzeb9YPNwgocCS/g
TtHfGdXdif2VJ6RXrtqBdMe6U/4R6w2kkJjqE9EK6pM75yMQqyZrt1CnUPCGeQ5R75Cr7hj4h1TU
YM6ZkBguZFRNAK7wmNlxJz/9CyWHeYTEflX7VpHPEBCoyi8zWOKVnivENAGk+X/benEfMNtw6XKx
mhwCA1/qSM16Few/XfdQPl8Vq4sTqw+mw3uaAUwv2F63R/CfWgEerKB5DACFRCwk2msSRZNJIGmz
53rVlAn9xRFQbBHreO9ZspPzwy7sIIzPWmqqgIEYr6Vt4pZNrXrZobZuq+5ZrtAQKc1fOYy1vAK3
F8k58g4uE2ql2erwU9zduDUY/1xFCmxkr3NtmuR+byemx3GnnpavY9ltXHxN4WlUkXSwio5GudMI
5XS2oB3BGkYsYfeKiZbtttJDEDFDWgwADBnjVpZlBrr4J7lKYq5mvZ9er6jw3+tYW3Xw7Jl3l3rV
lJnnh3TzeYdvim2tV8ae2WkbFnsg7OBFYRpRS5tW+Oe9saUBVIP+zR3TIuVH43C2jNG7N9Xe3TNZ
ITP0EX52Q8DtJGtomEeec+rKlNFDxm15q3drFMhZ4atyGjtHm95HpbeDpL0XMSMUHmVdagFUyyF0
gGCHLLeUYe6wK0ycpNfTGGFABWbbo+1gqjZpURsiUjvJ4+cK5rUk3OjzN64u8e/UnnKCSRZpFFKc
4h7lsYMZjVGRaBp+sdHX0JrGNNd+9RibEBAQN/DyMR6x22bhv956R20XDHVgg7jHARRy9NExMiM9
2+FNgH47wOi1ZAbaO40TMtaTs0MsKdIkMfYcKNRj9xaqxnE1Qn1z7jmRuFReUMlcMpacIofnKy1f
FpgjCjkCuMxNEgiC1lWoIkTvUty6t+H02tS0SRSip4xyXX2ll5ljgbl5w96EVZYpnMO5P1EFBQG5
YSPKImp0aDCjK54MiMtJOoyY4rhoPHigMzWasOotJxs1WdG/DwcVT4bZ2MHz1fa8ABtbcKYX6c2n
VekvYFzhOZkcUp5BBxafYMvC6UAtyHj6lWDpMBRPHb7sGXpF41QSbKOBu6Btl1kVYPmChWQNHFV0
2UpUYnbBnCv5j5WZHwEi7X3tC+kx6WmiftUS7KhGJTDI8p0Hh8ZMJcYMTJg/h8w+M7x+5K49nWBb
sS3GEzvg8NekIHxFVULRzVx1Sb/E4j+eQGjNG29STbkZtHgahXwTNN1lQE3GonMXsVVnfwzcs4bM
hojJ5wzCpcYyVSPstUxfGhFlXsnqGsGLH44/OV4H67JOFvj/WPjRAzRsrvDiMP4pqLl9vX31eiLB
i/nYCqjSP5tewp5eENvwb1ePb/g6lG9htRgkm7y1b6gT1NeiU/1k+FUf3yfSc+HsOXwCnmWjsjDa
MWDXZTb2T+wfYpWC0GeyLDjQQPMfjWTjvsVX6sR1+kkI1kmsIddgMJZ0aTd0DH0JUZAH2dspWPrF
D7QC7CfAatkELd0xsRUhgqe/W4AUDAV/3J+V8JUJSsTuusuEGx9ianuV3LFSaAsPQGzSpn1QPLE9
Im1OURk/h0lfR74pbg2KaoZQiOyAhSfyyQrjxnYIqQJyOKaqfC3vLavxixwNiqauTkhj8EIAwrVH
dza5COgm69o0agmmXIliaru/pgFIKHSGMByu7vj9jnC0H7UaLKJlAPU1Y6ELkmoVCdFLy5cZyTbQ
BYXX17CrxUqyXx518R2pffWsslVgX7+kkrGldspXdq7+671nWtMLdRMhzwv3/SEIcmRdup2OBCWI
R709xin/girFveOl0Z0I7uAjseY+pnni2AO87xhVkXOup052vUUHMmLs1hsU+rL4o8CUbAIshMc7
Cf2oCu+QmxhXDpTP6HwwpjvbDWauksJ7eDd1svcYM23ogoQtUGoK4CQof4AY3NtEzkY1DaR9PH7X
1B223lGTSIigHaSsnCZuZuSt+QkfzxQuI/sxng+kS6BwE4UGae1AD4xJyvvhNxR9oBgV8D+wzC3V
+RhECzzdDndKEl093s0uwM15pRTZr65irdSiLAtKvW4cDVn5BiWmwA4aOSDevSI5aOofvzqZFAfa
mLizk0Mn6WAKMOO774sqo0SgwziPJLrdi30GOKtZOyBWItd6o6hRmsKpsxvUrtFqDiXrIHc6aL8N
sQ6OnNTkPc0HkDdx6CcocLtCvZAr3sPIhtfNG4JTd3+y9MbKPpkKXl/taNffZ3yUbAL1J4BW56/J
YxO5rgipc2sCGHUim0KiHGQy70JuD2cPJZRZhzxI3VWu+kgrGRKwreABKkTfpi7yJsvVaHeM4p1y
Hf5M/Wlu2E4ca0B5grrvMUHlXo/tRm+GvgzzFOkU5LXnmYSEGKNQdeUFCzyr159CWwEmQ5Cf4wCy
lQSyhkMttvzYCsWynqAyH59S2jXdW5VvhmNRDwwzA2IQhui4k6sLeIXANc2TTIh5MYjn8ZYxv9uz
DHzDka5UZFh3ELn4cvT3wILyhmd3Tdh5dR8bkw7hAx2XIY6vptpebc9B+wvpzrGZQAehenDK1U+w
xGJiY+t0Am9nD2y9GGLCq/aZuOvFF0m2RcyWQFKIrQcjeFzqEBDtYyq1PbTSlUdn50qNcSLdAD6d
SVWgRy4ZjC/Kxhj8zjZ6FvnUO0qa9YTOsCPm28OrhalZd5Tn64H31xqQfxN7wpDiYMkpj3fOpxU4
+HruDn98jLgj6b49D5og+OiJ29/OTLVhTI7lp6zvRtA3cMiE3v15zHOQ86giadbbksDOhRusOeKD
iD3qlaAtfnLesr0agmpbjZYtm1hIIXrW9+/1gEWBYNIxxiTYVJhg+7yUSJX77gdje8EpwtG/42s9
ndVn7vm3/q00e0fNDc2/8olHU+sLX2LgFzWzGFWN1I7YjBExqC/IOTbY4KWx2LEH4rUHuW4tuY4Z
518wQRYp8TuRehLrmVps4NZh7rnip50D86vQLxyDq7UHHhNkHS4odrIbvLSVk7QD+S1Mmi1Ixo4y
z3xrd+YyKnC1hxlnH2/MKRnNeTf/JgHYhplSDtk5kccodljftv1LLKTCjzDHvg25tJvx6zbXTEfn
cPB26wvnIXgjEFikqPmZDISRoStMbXTa35RjR3rPxcNNa9HervuKokUfkRMBGMhJfHprTl7opq1I
QFrQ1+MDNRGiVwh1bVmCN9TrGVqg/n5tcmFvp8o7YPdbnHLXOFHbel/AsFV/3M39oJ7avWXtINsr
x+pQ+KOo7afBi2v/txduxV8tcohRhXzy2qghQIOFqIOwqSVaDy4nUKRz9e2wUVQbZtyZ6yKQGsAA
8SdxI5bU4krjPFcbGe2qruZEXGBKdbqZqRqIfMuRekLvEiVaxF1QhccQaTUtsntIK4v4i23bANZu
QPgmnNZKBrwiWg6smIcgzaUC534nevKLOBUAcgNsNHMgD0t4jgh+SyE0Q0Bf84KRoyLWkhoPCYOP
aaa1DYYn0yR74RKfGo8DHgAYRCLRccwbWdlhleeGiIrRq08WA+qcaO0XZYif3EJ68M+pFNrtymhg
6cuxYOORhWQhTb2NZsX+UZXP9G0+kb96SHqumGDmGwIlEBJm94psNtS5vP7En2YXqTOpvFlAMiVH
D1nbbRE7F9OIohVTlICTHNq6bUZc/p4EyB+pT1FjI0SIFjV+Jhw9irl3UQOholWX2TanCBudkzxQ
Z9Xl+fevehNKqP4JkoKHbkXDb7AKsgkCajhvJn/hBQkYWcuBMtEZba8rlbVBY7580zrxZp9IGTa8
tFTNtWBRLDSBPK5H5GXFuHfFozcTebCJnDpifm5Ek/Wsou5DvlEEcTbi2830KO1+8gnt93vMDZQU
UXkCMsIESlVcf8FAAgvAvEbk3qss7S2BkFiY7tyBG6eTWoXaRq/j3lUrHbdNVrF3Ykh7g6My/US2
5AkK/7r8AOZupuXsPhFDcRz+wfkqv4dgzI0bR065XD00g6nAoZFesFD+06EC0Uf4Nj0NGMFOfuuO
um6r6OFXns2os0xXwXSILYXHAkaIy+N0ptJnFWTkNaPPaeWNbgXk1QJwP4aK+5dPjEa8W9eX20uW
IVvtZr+5DwhEFdStWoZXb7yleuEnwneQiC3BPbwAsNAQhy/bt5m/aAkIGinyNM3rQFOMmsxE8srQ
dYdf0qqrfrWFKQ+jnvaqkk8NxQoCOtywRZT5Xrjo3RAc0xFYF6fKvZ/i4XajJKwgoG/ukYiR3cex
1A7OLX3c6mGvpeYTf5SyOQHQU97olVCQejkHVuPrfcplxAK21S4e2Y+uqLTDYeRB+QOTOekVIlkC
gSKI5p9KNzcViUnq4sSf5kHTLE6iwhL+M0d/8mskgB/TeRF1ARBIUvvywLanYoEIvtCLxVyGLxqh
PzxpnT9coJTu5w2ATIXxXQkByTwb7udbZrpDIo1hisOL1s5sv9PEVZFIypXN+HLmzKDRxSpAXKjM
2H/FuAVj5E+8IztYMSi52iL8NgNOqsqziNle7+9cHwvRVUyiGwpbzSgVgl+xwXnRTxSS7/Bqd+0x
V33YsAjigDAFmW6WHpI2u+l+gTgWrFRylVlasy2p3eqaakpn33Rp0HbWDm532dZJwqEOjJbGwgD4
2V1xvLxsHcfQsA56mt+QxeZ4Xw3wQHfegziJ4juMzF1HMMqFgrYLHONzpbcyjU+/1fYP7XZu5kJS
mhjiEDXO6LybL4ZchsdohiGZLFVFRDf7qCN8zT2iQDpZWUI5XnfabH0obxWgHj3ZFkVcufS7kOtB
+lcK6nPRLlu65pJJBlEJDs4pK7ClC715fHb+IyBR8WMYz5QgFvOt3uHH7JTTo0WCP2VRP3nriXFm
G91vIYSjdmBoHaCkF8NscxL3iEQdTylHzTLvHL3qIuymluIA3kMJi9ovZhG+iSWx3xa6dFc0XKZR
YsoI5AG6BxM4xcC4UxWgicqX18mNWdRA/2C+q1ZxnzaJzyuip4LaQwgBDW5grLDIAZM7DkKdppqz
ip4flazRsv0Kpv9FJaTfPKGJ72wvfYW/hyiFVb4v8ujM3hNHkhI26hP8YvAH2bemzrika/q3kPsb
VldTJUmZ3jas7okhJ1Kkm0CRLdEmWG3WqxKUc9ha5PJMTZhjAItknmQjJ9S+9qjyKCcaP9DiFLll
EKZYzEQDvoCNfrHRPoe0YK7DT3LcDfccjfopOJsLySzSYg61tAsb7METHf+UME1HT7tsTSb/yDJ0
z0DoOsZGX1NN3zBCkgW3fkfYrbmRMCnH1uc3WeafJEhKTUuy1yDvSFSC9S8avoPjwy+qjCPh4oeE
ugttAnTt+05j8oVtHIFMd+TZcdbLX7C1K3BujmWGxpExTIoChIWDlFXsshYSylEYtSdjRBTEux8A
llboQxkCP18FKDM5ooAf9GMdr6GebELFdq8PrqHqooie3qTkUG6AJJy0k0X1LINBHJRZA1NlbtMm
OcwzEvEY0BiFOGSqRObBFG1zED1igTjsogs6Zylue9b5Rqx6zPdMk2W54ViNp16hx5BChcu8lXvh
tBk9aV1xW90dM6WgF9N5N961+3Fxf52Q5SGqQW0KlhrBAEN2TrwpZ3WIo8Y7qbsbg6f13UZAOcJW
+NaO0TJh68/VHJlOUfi2EeacANRNoaL/0GY99QQLjqTOOMixUiAQR/zxZkxCStp4zD5FKJOyqZBe
4Y0qnNq8eCYdQk9YcAk9yTBTZYD5Fz4yE1pk+nJFdGO2buJOfhGYG9Wc7pUSkQxYPZ/Ak3i8IyB9
UT2N8iTOcTmSGVX9wFMCMTnXzHgTjcbBMCDOSRFsIVI+gj3lqaKqDIJHcsX5ZRiaJ9cdOoW+nceY
z7ZPa5fiI9+CaEkfbL8z5SoDBY0AnFoi+GRRUE+lgH5bpl9WszIheFWjFcUNmTdmoUms51xLwSDx
0CKOjl6za6U07CAlJRa0uiFR5ZR4QrNxoJDDZU3d7B/oEl3fX3gCG9tBTSrRcPizI8LpB/MDXJK/
TZbQyHSpse6YHmLdOleZHUirGJ6kPF6UBpiQCyFY9f28LmSnHaRUY2fssfC+iX3S1vwDw5RIKYK1
+vdJzv5s2J0ALcS2kEIGEPjTC6sDrtNclb6lji1rHRDAN9wC2CQrygPHgLNvJ/bJyPLB6KVsyiNB
/pLfCdVCjLfiFlL63cIJvnE4x3wlx2U6REgc2PqkhsgfGitKt6xvrjGlLGGmotsiiag7YrLNmg8g
FzYnQ6cPrMxRqnU1c2o4wnYmQ9iklHixAf9LhG3Jh+Sh/A3E01xt3X3ZN5kRXRcEabqhos/KGfNs
e9ktlXES3FTG3z6pnxOuO6+yC4w0iJKPYn0wXPaAFLM5ocAdy7zvAOFQcsX755p+XQTz9zARi3Wo
jziyV01LHMT4AQ86W3Cs/qxZgmUwjJgh9I4naxbA/5wIdJdQY//jwwLgzX7iea2Msbps4UT2boRc
dOimdxgMfcXPZA/m2eVHlGThd574WQtlgX7bQV38kSzhR+mbv6GCtARX8mqznIfoAoXVHlvhDIQr
yhHkZTrYp0A+FpHq3zKyL5+3Bj3JC7Qkl8/SGytx6Gx07SmEMDqTg+Y3IwMhxHwgQ9GHBzBIVKeh
7e7fMRr55qDubaOfHtu5vUrkv0uMcD0jAaOwRye278KuD5A2IBpAL4CybqHB/hv/gtwEYme1jrbO
TRvc035NMcLj9lk0cDjsQT+WIc4qmPuMG8kmSWTIvpAIzR9vSu6iWTmiGeqrh/rjpZGmsbIckh+l
EDPa16h5mKKniKS13X33lViunoduEaFz6FEG7YOh/s2OoCs5PO3NJsFK+bxM4w2y9tBY9W23JzFR
mUKenUWlTH8AewJgnv5QWLJ9o7mzh6MVbCBwc7J8eQLMpC+gZtus/Tsn1kOUi33LNoryyRQlpcjn
P9bcoLVKdPUqvinHbHIRHwyR7uDWfBBDMLiZL3TjC8fkTPrmfgH8fXPZG9vQ7nX3cV4SyYGEfNL7
5Nr35hRduGQwVNY1wIL4TRzq660un/7j1lifv/I4DuQTjgofiqW2oh+7GjxRZnmnwKcDwWtT6AcG
jVVEC1pB+3+j8hxzQ+J6Tpi8sEXWmeooskCjtoTpe7t0bna1RjOVFX0s0bO/K0ev5nPDnsT7B0yL
gbJUlh3DJ3k7VVX70raRJ+B8DosB7gdYZD/gugAenpQu4SnT8SemVIdOIeOjxoFpM8ofaQLy+jR9
W53H7eLzLx+Ody6UpSchL6SzrnlblKeJlWceqIjvIFkp8/QRezoeAANsI+RPb1iSjewLCdkCXdO2
6K2n+UIyOa+5/AJjLENQwbKbWwhXm69sJlnZr4dRofbwydAV1AZ4+Igq52WALknm6v45n1ZHXw89
fLtM8JLvt/fi2fCktcRQMhbBJYUaeo2WDFUaCGyukLcw90YB5Y1l/u/gYt6Tlsk/jf0AEl6yd2JU
XCaSPoVHBkDhyKxD2dXINbu+UaDITiazQvGYDFJzMvr4SfHu/t1TaH9VgHfYRsCCKt6F8nvlyI1m
NDubmM499T0EHNwA63BVnaetjGpPKhGBNHZNMW67g7Ho249DnY1acU9jhOTeS7H4R161pPoJTt/c
JuGdKEjrerpDk0/LelPERofZv5gd3hnZt9T2aRobzBRiZ97kY0K6E6GJisIdFAp1rgx1tfLr24ai
tRGXSGMlccN5F23Gyevn70niq2aDfNzjEGSrVs2ZkiM94I54V7dNkh+1Te2jZoERAZcdx3j7RocG
LMZtluS0fOMT1KUtmWT5QHBJ8ilOEQB2Rk78XHFZ4xLAuWTG9NaLaRK4uGULW6O7MHOpX1n/PORT
2Y5+513U740mUqa1AsZ02Dt5X6GED6E2VEBjnJIaUNlbzryYu/xWSQjGn5K3WyGtIBkdoMgT2T1G
Z9zFz4uR0KmwYF2ENz4uqy0WB3mzTRuiQ+ivfBnSBtBk/yeQGxRhhZyPB4ZnzuZC6WZTWSpeBaC3
hFxJv/mkVVC0GGAUKZ9RhbocLZbVA59awkW6oLnj9jQwZUscgbdnq/jR4rPa/y3ehp7uL6B4AU6v
iE8PHuNdfiiJveUS8PEFo6skXfUcUaQ6ilW+hxCTidpOU7yW5nyZXGmbQM7sbHrb5bRYBBWGEdMe
NZeMZlJ0Olase5kPs4ekgSy433IoeBmyJFg6Kpxr+2v4AuGDkncSYMJUjLo9ID5HKnGD5lqhh/Sf
/dtkehHcdIHLiIPlfGC4mObtuuFy5aOQTqPHAKuvinl2Y4vzTgurpqGL198ZXm+QjOoHIuNqZOS0
uPh4yE/3/2wSdjZaOx3RAIm1N2RJw5Zsqqc2BWrLKCZwEegvmDVx+xVcPVeAkgJmXT5i07WgLTgO
E1Xpl6e4awRlmuP1XWDBh22h7E1EyIRHsSkvcVrCX6nvlC3YRSUJfaC619vcmZ2yDnvdnI14llyF
ExRv1SouzM7Ti84UoC1sPU11VGLfy9V+1JyOMhorg2s/YD5o67lQ8VNn1FY19g0Yk3cSNwfCFn7o
nIHBKB1XrMJkvnJ8493rnRVWbCmG8ltQyxxk0Iak3ON9QPS7DBAVP3CQNYqcWpceOYFHDUHC1Xln
TdLNAKwMgmhdk/bUiS+3U+Vs6aMB+qmCLQxcEeFLn2liWQC9yrS2nMowy7hByuo19C+42WcFp4+P
HY+0lMCN7f1TF32NaD/zzJSiQwttkGYTy2Cda+uS55Bn6FQE2BWDV45D6OfQpb1Gq9ZumVRtwy0k
jMdYDqMMUwepnnUNtZc+A8+7O03gVUaRO6KVRI7XQVOTDHhhh1qltV194fJj4Fxlxs47uEbYlUJ9
ggK8UbsHxLpJCxBAXZYv6nuoWe+l2W1IZjtQ1ubxCwqN1Z9bYHWJztPJDZ+Z4mLm3JQVEokwewxB
L8hsf8K1KZQJa/tfqJN4ZHJb9ntXBSViE0Lzd/QWdQ0q6ZBy2P1DwUGp419XmzDQF+hzu6E4hlt4
7nELyh7y+t1Bcp3pNbugKG8F57WHNvkauX0/usZUbNhbUwh4V0HXIt2iLITR6oHtVE1dwfAPwLCp
4ROqYalPLCzk8w6GIpoh+WhFd0e0VDW9GevbAhGIwGjXhmPBDTZZVmZx5RgNfZW++NPIgZlSCFBD
fGPXDdq54SQhqgrTbUAlj2zRSsqVzr/jG1WLQ0xriU58wMytJZXQNyidsDaycxLETsSt7p+xbNS2
cCmr6cwKB5ojfMxnwULDZ8P37JcAY59E55mwdK00FsTZZkPtkDsveSJMeu61+D/TI/uABe0RAv5H
QvdqozbDVLiOkjaSnLdYSswfTpxz8BPiJTvWt+MQj9QhVMJm94l5uOwp65AF1Y2ixZMuFqTDg0MD
BZ1OHQ2kT23uS3ISof76zgMfmKTg4FcHxoeKVCwY6Ny+k0/6DiefgSJZrEEXV2igVsp+n2lUnFt8
mgx0Xvc2wHYSpezXCXFP0WXIulIlTXmZPc5xQK+tV7ujLEcHk6D75Vhnswz/gRebA24u0BHeVR5k
fWsA5xwrGjC828rxMmowcDHgTlWTBYfG4bRq+gajabij3EVSjY54YXQDaaLIqsSmgXI73bpEOsmQ
eUW5XwSAEMfuigutAXVEJwIE8dpgWMwc2x/OLTivyvVKut1KQXXs/NW6CWYa+Yrh+qSzMamtAvR0
k6pl6bnJW1ub1SkkNvOnTs0uyrjHo8sCSZVYVALXxFG30Tb9vRnZr3LueHJMZeBt6IWxqPip32lc
85FiZqrgoDw2QOYRyep9f7rfzxUGLNRsRCa7E9luyTk0jRkhlhNJ3JW+3wXxA2zBZEqdN+rf7LMc
cqjfitS/Bd5weeSIDe1oOOWiX/FoF54olyzaQh2i3S3gDV237AUXd16dw/WbS6eu9snjHmd05ol7
K+vIPlNJr8mYx8I7AtH8+uSm9aAiyqX9z3yOfsdx5Gjh5wPmGA49GxPmU2nm340udzskOKKSPRw2
v+PDkAew7/fBZPOJ5iXRaFKe9resFUQqhZjP8GzIjCN+KQSliF8PtrvneaN/wdZ2gtGCVkjuLSE1
QVjIem2hYTCSogShrYOMvdsKlFhf+DzR6jnbqZiiixJqbhp14mAEF9FaRMb3nhiE0ZQGTKb1NT5L
UXuEspLKcOeONSQDnufYZew5FcQoS9lOLhP5r8t/L0KDlZh4FG01lPOqTJtRPf5wnG8mSUf1EqaP
SFJ5ISClKfoYMegRpfw8MzOzmFacx8juPkk+rab5MRMagt1jvAnF0bAhqkoLW7vqN5OsNglvNSwS
LFKoWqCUI6X8KsGwE8yS0baaOLvj4BEvy6ySEETVLkhiQFuilB8Ifjo5YXmQNICJNAi2SJDpveiI
kz1lIzVAtrzct4RqrH5agwuAzNeQyV+aLD35rNwpLqvfk61iw3qf9CXoDH1z5i8Sd4zD35DGtSvN
3XkP6X3KX+rvzgHCd16BqS4CDYo+6dR/A2IP3chi2kPlC9GS3qUR4rgd0bilksI6cK9cPN1dIaZC
pe1w0gSfnCWs+R62fiR/tNmwzmp40k2IgmkYA1be+Y5dGwczynH9TiGc3EdzT1z2MnST/yFTCZhr
CyQ48WPwVqnFxo2Ne+HfKi88jgaCh49UtRqKF4/x5dqHbnAsWO3C18zGpLRoxdkH5+WKTdBQByx5
SS+OOGbuCTTZJrWK8PX2u2jfcghZsYytRbzSrLKqxQenHCNxX3XyiMI6ysxg/bzb++p31MkErphO
5f5Vf9XeNzSiFukzXQ8B2Fvus9xxS1xLGCLifCD/tBYMWpa7SNt2U+F4EOYxRIh2nt9Tdynf8chL
WsWB3F5dn2XgkSEl8c89ekpBFuUtyj+83v68pXtsBvZMbtrtVG39asBodNIPBXw3APaQ19TcsrU2
DcHJQwuXP42/gjYOzh40m6fBxkqKs4CsrDXuTmY746CgKr7ZqcLqAKmGsO9iZyGi22jZd/rES/sZ
Lfh9W21FUcJdIncVHzgMG8mhiC6/UcDKSkQx1bbuW6Rzfze+XBEURSrk0qZQU9ZsFMs6kSWF/Hx2
JyJ++FOQL3lATq8LXrVFkuJC7x8K2vUSlTuKBaXZ6WtsasYAqXXf9KxtpNH8fIS2W8GLKTGFXK6g
4pUz6C9Q1IkEMiOC98sSeXkjpT/nRIz8OJil/OupejMR0axPlqByvfiUZt2X1D77MOv9SlKrVW+g
/fU7iJpLKI53cgDBuAkrdLvUrN5qYP6kWvHalHrRcwf3MTXJzNBtHEq5y8kdmqtQRCIxvkz3XntA
dym18pSzKrXcWxv4wZ1p8YYhOvqzAvZVmyFGVtxT+N0I06pBBVsdnAO9DE8G9OXgR9WjSpX5/wdx
/k0QOkgDkCbMHVKqRqE4kcOXO7BzStTbie56dFnIZmH4l5C17Cb77XhmpvJzn3FRhqfMBZfT9VyR
gHNfKLogELY8q/DKThTGc4OlsxoYyX+6yzHpl/P7ELjC9Bl5m97a5v2MKLNOFSva+LcWAIPqKtSJ
i3cUoEK2BEbu94DQ22X5KG28PEfHpPFucEVv6CGTP5rHQuDOAtTjegycwjeTPC906Bb4GkMt1BYK
ECMNw8XCzEKi4usd8RGYz7/fSoyUqk4u+yYhRKeNXpK67WE+b05mt52xmT7819YXLgVSvSZf1Umy
s5f+u9RIiSRdFt/qYfAUud2xmkbG+MQeagSADqWP0C72TDuyZLh5OI0Jq1y/vc5XO18LF0QDueMo
7xXxawj/32ZA0wtXXMynpzL24Nnrd2FVbC0TboIK3nm1m3XCHfyuyO75JnKB3WvanvhJxbB8QlJo
u3vGAU597jVcT+HqIjDC762OdxFmJTw5qIDISWdpya4j0O6S8/dst/Djl3YzbM08MLFiz/bArykn
ai9ZkwDw2aS3twwEModyEviKeTLDxCWiNkldQDRNTxmrLNIcxug1KLKAmwvejjidIZhQ/3H6n5AA
LnyqY4zGoaYivdfgn9DQQhtw3Boohopdizr+1UkOiz+KeAv7q/QWVEZ3MjLtDQ3UNhZLM1INE2KD
mUDDPBG9Nuu0SW6AwJz4+Ist/bxNCIT7z/fJFophtqDPjwLSI1brsns+8OR2ebq8hEKlfIT5ZfCq
49x3qNNFZdFODKgEMbECaATbyIuhWq14mgqTp19ZG+vQvcifhbW1yk5TFATct5VeK16obeb4+j91
GhxJ9GO5Fi6gNYK5HZLbNdvCTL8oCwP+qWryedbcnrb9BE5B5VEpN43lfbz5YgB2dmwsrBixY4nA
CAzQ0EmC3dCWn/4QjglXZdmfho/tkg6POJPteUZjqIowpNdbum4U7YIOr/GWhL9QvpcRQ5+EZx2f
nPE7WeCdo4k24Y6UJphLd0MTKhgPmK9oRyijAOJV6ka/nRw6tqisMxDKOGiRakzKLWxuHtnPfXGN
sZ3eHyt1aHxsa7VVtVm3944+f7ZTxyVZEQC4FOAIVLEI9XGyUQAqNMr+gZERWofkC9vjKVR6u+o0
iC/rT8fN+RXszmqa2XoZkiF3H50hzLX6xFHan18RjfryfiJOA4cE64TzSBuai27N8PmYyN2j44QL
7hgY1/25nAGf25qgw2VhSGq8mOuhBqQIiw4xOMJWUGDRpTlbYSFx/6rMFgMqFFrh9uSq6iTA2ogV
umEPzNHaNYzVBABYFebPfqk30wgfXpit8bxJDZFNIrjf4pYbS1ypyxLLcrCit0fu/t8RpzKeh1nE
sHy8lMafUAF3T+jKUzQ2lHBw9f2KDm/FeZj6wjVth+3xKCAlfOKbjNd8ynqOgnUZPLRi2dcjDUyN
NLr/A/CiZSwk/jd1zVigJxTdv4DQPkLVQAEfZGQv/8+tGd1FP6ecPUdN/sC4tPeDzOdP4J/8Scnl
fp95K+qZL7uNfBr+QS1rNThYJRZrU7tuPqnmIs6sj+ebwbeiCkz0A56c3eyqw37RH2dFgLXvpzjj
9SbhZS5EETFZBxqzlFYV3k+VpmiAf21QK+zmwmTYpjCFxGI/2MXMM2JWptgH4BvVbzbqgATQ0Wbg
OZaao73D7rY+6nt1KDSePe6xjY2fqbzVlSajYiB+vf50hTF2//g/VZmb9h0kzrl5L5MYmpqj86PT
AsDjRXSxOElpRoOl24y+l7VJ1Z0MJYCz+EFBMmUelYt0ARq/ItVO/wb31aSH4CSowMrosoSdPSHS
TMdyptw9caDRKbKqREn7gnLw31HYzG0m5aSY/HLsiY4R42j0V9W4yqPMlqgH1+h8REkCAJYRfoVi
LBGJzFWqzlelLibUj/Jj2V94oUdA0HpyQV4eZbOwRB6APM54c4to3qW5IyV9qskaigS9vk41ebG1
7P5P382DX16q8Kga9T8efEhNcswZ+tq+ng8g+0d4l0lnThKb+7lkzbX0hHaStAFi9XBl5YrOW8Qe
SrQ58FIENFt85lUNDredcULfeIhprZ3jbtuZ9mOtNj4wgLoQ8TLjPocV2mL3FfrMplNVtz9bbA3J
PU+7YCFN0/91y7+nBsQz41Jv9eYef9IC1puoIRWc3DKWwKxLOiQ4cjN7R6sBZFjshun/XdZmzkqe
AcL9efxlWzeUHiUU6JWQ8hUL9RLxsEyOHWNjseu5BeJ69VawHUD/s40u0zEyHN7xWM4s5ZiuW5Zl
TGvVtndjcPnEPA37iEHVJicZUouKUMKK4cCB8Zu92GiVtyIianBNM9uElquWnoCyWEVKccUhN9Tq
+MJzV7Tvl3HHsOvEDME41uoiDaBpo+z30gd3F5fBm6QHl2vfzUaFuRBQTGosO6cw6Oswyutg/1vc
HeE2y5RWmZaRBl5iSCC7oKG4hScaPZ5ila+RruP/8YtUuQdALa/mCytT7k37UahUo7lPMZomdnoK
Cbou43O+yQf2dIB19jbEjnUgefCATh3FGjY58B1kdcPmsrWjAtN/WFsXGCvSPMnvjDpxuZ7y/FB6
SoQyugKkK6w+TJqI8nQV4YpH1Dgblv1zaUz0EhfOxqKaBdlpDsKX6nxTreQmCatrw2BqU1rytfpX
llhl/PIKcxpmqusCSzCPZkPxFGJUVX+Lv2SHVQJAzYQFR9IPaCdgB4qkmvDqwG1FMrpjsrQmmoLu
ydKwnMjY5xrjekLz9q5uIfkUyjrYCQDPNphuNuLrsfAqtnEulc8skVgnFQw6ohaNVuhP0RIgnQP2
wz1XhRI+FJJVJAq3wAJL1PaR7HO8vIzOU9vrbDpU3oLTB1MtTd3iX3EkoqadpdzalVvBurSPVE1Q
p11+it6g1HwjG/lyPPrfZKxs0DlwiINti81q9giQiesrTIID9shKiOMEkcSeAN9JmCCz0vFrzhbf
Y9P4Mc85pw/PRNsv6TgeuHjUEFceiO4rzhsOCa2q3E0BNrO4lScwVDZVvHojELMdHKrWXpVByAes
1w9TbuR+1WLQ+5PmD8c2fDqT4HaGbB6LsceTK4HrsGRINiuk1FZsJXtoWj0Y8gOPLSIl9Crlq9qM
jsUKBH2OfCAWUptIxuVIKKVE+msOODVRFhJi3SIs/EoSBdJ2kCyUfFLlUkYe2z7s6IX4irUnV1D/
DKeHGS4kNWPOhncPQu6mv9HUUOt8GEZ6kaq6EldsYk/hfXATCw95fu5d9IS+/iW2xBj0teQrFW+D
HuwQew8X0CbVwBgL/CZWrLQ0/e40Wzu0iEFal7LUwRNX78t703O+8uJTocckLVljcRqfkA1LSLh/
CgbUXQZyDiOnZC3ZuYrKieQIIPVXNwpW0KyTNkn80BiuM+ZIOW/NF+3wnXOEL9g+bbdWtJujUZuW
IWWuJ5C5aBhQnzj1V1i5UpdS2Pfc1X/MwqGnnaevj13Q0YphDk0ygGoKU+ZskLtVo7LeJnaHrhhg
kP7C6bxe0WgJey1susPZH+SBWH18oF5VIindS6r9cHrg2ABCSo2QMiXuAVw62WsJcs7toUseBgm1
hWYJOI+jrBSwVZJ2pbcoN6UorTch3nmKLfT62o4E/1jdYndSic/kIYIGuUOYYh3otqC5TqkPCR4O
F6qaCid6v1lMaAonV1PxlOlF/B3pzJ42vyNx6HZnAMD+m4cfLnQaWKnkmEM4vgYS7r1ovFOPY379
ZvNCq1gotGJrVDYoSucEbNG8fWkkxz+3+V6SFYhVpGLM0TdWbLBbd643sZ0E3pOBOie4y9K4Ym0I
2Oai34ZTPVVHPRz4Fk+Rqyv/wapRrJjwSX4nXlKNQ4OIsFCft/OMaowis5MqcowWE63zuKhH1YJ+
N6xY9j5/uU6/d4lxw6qm7xxin5iBzIacD5T+kIJYYYqZpVIpmHqiD+ajh0OR5SNo+TFYyC79ZEC1
VhTDIr69m8Y01bTAUzmrqokQmmSWpLn6ihXKriDTRfWoHIxHSpbVIhnJHgJKxcEWf2dDtNw8ayZz
/um/47DGyQnHd8BifjlJbNHlsYQF/L8dif7Sa88fn34Onk50AR3DLvHU50+qA3n/xQDVY+G3MLog
4gyOlBkLFKjISanLCnDuuaNoyeFl0FHtrP2KNl6qffwGIhRTNgwhK+5Jju0E3ITuUkSob074xD/Q
too2TdkE4ggDjPtVurIgCvJhMJYxc0ZNm/HePgUrPyvJUew1FeIxKUbokKZ0/GNtcp8OJdwJM0hn
Jd0iDf/84gyMIjYGWPbpcMTPxBpuNTBzAcOHooliPIWFB6prel5/+bmyiknmTPPbfROjsNaF4SLz
4wBsIIJxhGdawgH8lhQ707vwHliSsMuuHoYNurzKl51XSwMdhCMOOmQzQNMrcX2jv3jk+wUbX6/1
2hi4tBDJKUOC7tcoxvRjvdu4JjIPICQENDHs4qRFo4HgCIzRuz1udohwHjdby9zWQp8mG4dsvdvx
o+MOH3g/fRrBLd4YhbNk1ykL19aDfAHHvMp9iA2XaETpvdyLlu/Y1b3RJklf/UpJGkHhhSrBcgXO
piHiBLUf1c0EMrfyFwBvT+2bHK9oheK6m8YiqCQ1gQVIgl8vUn9XERr5Pb8PvhBKS9Chdkwev3PN
0ixnf5EyxZqOV+Rl+yGFWrB6wmqssdOYuex2krrGKGRpC0B5Zr2pK68KlXKFjC0Xd+AImWI1mxCo
ztE5k7kd/q/VtCJAjcKi1Yfv3zwsRz2MHWUE4wAyaFIYQErxPlvNUe/ic5pb1zhDhhax5nNuLenm
xCG7NneA7S3uiclaEB6xbGCKElwLE7IUMbO9nq2jPmy/WWEBHg8vQDnRsVa48FyEV21Koga+Lyg0
j36bbM2vA6xz/E6YlDdkwswFBCuWVLUutjvHHofzlRb6KSpAvLgF/J7IG085EQXG75B501qjwpVH
UKwAYMGWRmt6uP2jAMKLeOIlgqLGzCDn2YLvKetYXMZiea2N0WdY/tAIgf1WvqgGtRk14O16f20X
Dw694bIRzM6u0mkQ/gGGKyqxGWnKQBvxuJIyYTENPDA4rKZpDTgFZh8eZHFNba+GgtD1NtzTSpO5
PcCncLfcgNAtKorTMqIOn84PJ8IqLxSDC5a8yFFwoGxr1CUNJi7o+veYTC5hDqCa1q5VVRUHhrPS
zMiXnxG+IaI1jRCPL9+6/a+HbdwmNX8731u9neJn9+ZTfRZXlMcNZNX1Fcvjrvogpfp4heuA3rSm
4Bn7fmIi5gNMbsCO/yEZHLzJ8Dm58/hi0XxUdv9Z9JQiC7koIIH2uuBCdvHJ+7E8FwDTQPdAil2p
aw/YUzcRGo99UO0pKYZF6dzcEXqIV1Qa8YVyF/E7SWfwPhc3NR3FA9iHcxVp7Ob/e590p0fT1234
8DQ+n/YKJUtC/fWiMKwTpehumywFXkuvIsMlIpPxAXblzqGpbp2j3SRsZ3+t+8Hs+Rwm4ejE3eig
xh80Lg/rCM3lK3z/tf5MKTCBQAAZ5Y6ozTpi9aHtINxr1X3RgMax7tc5JAHStvzR6JDG2pFqq19L
qvdF8/bhNoqczMFdnhgBNskAkfYofUUepvbXbaeLC0m2SWl1w+uRoTMgB2vpZRdgfCDDrIMH9RcM
PbjckUCF9XKmDRT8X/MoU//Y269I7iDwnJo300e68LQ6ijCPWGKewO3aTXDor4r/J9GQbWAt0pZt
ZymWcZ2UBomENqp6qmnvJFvKjEdTwyMJhBCSfZn9s3YtwfwrpVEuLYfr1aC/h/XvK4CnmcDwfZ4P
1e6VS/nv9ntVQc66mZjbu7qr9i+Kt78d/aE8mf+raxNAg24s4oXQn5G/gRs3gr1atgJSVw6WjLQ2
36vB8iydEAl5hbPPJN5V1GBvdlDVamuKYdGtbtFPdSJK04zX/Juy4HhAbOQcvRwWaVgh+T4AScyv
b8MFCAAX+O1N+0fAwronbgdPew2Rhb8N8I/PpC/ub3LqK7ahy3LmW62HaXrh6qn0mcCnML9ObpDH
3iJX22VfdfiGRqZ85Wa1igTeeqMiu2Ur2D7tMdi7caWVVhEvaeOYeFSFUSK5PCgZyCNDVthH8gDt
xl4CWPb3qt9AQ818OmCCB0XSaCsj/XtcLkWVERcIPoEKycHgMNfHlj7BL2M130cJpzl4ezADlYs6
LE1PlDo1iGLCkHC8OydeZtMbBc/HvAWQiqfGwFmmFyZKYHjsvkl+o2TWjcQoBHoHMzkrlC4yMJL1
0HBv3HMkmKBw1cq62WLE3GeVzPxcS/BT7gUHiavr+9oMub1hbLr5yL2vAKRCL3wQUuRDjrCnHR8P
AwRwwNDt2CCCONLaoh6CSPRoyx6pQ4W3YdCvd0gMT6tmdkIipsFde0H4R8+f5SY1bhhYyaN3Ln5Z
Xu0z+q3dnT4o96cHvfzHT+n77k/XkGTcas4+yuz/6asZbEC+JL3xRNY9ymnXV4CCBH8oBcWv7UiO
V2MzxJ2LX7cjj7+HpIcxSSqd1h1khPf69fx25UA5/IdZaVvnw2Xcfpu0tBWPRpiQ8/t7Qt2Ib/r+
qVX7Pc5lPTtJcwdQ6fF193ul1AHNXCKOXKS1Fm5/6snWfMNycgwYzlE89gwQFsreScy/WX10Y7kx
BsfJ0+N1HxNEx56n1V7ixPVbZ1FdAerSBtCZTG/oHIcCIuuYI8IGImEII7n3aiTpgNxUQBUqHlRl
uf9xRTRpakMFMhJzwAqPJDpmYrZGMCyj38AT9PeZB5PRltmZxP7oG+Z8ASc6uDMlDGjCqSDnpAYt
nUepz95OA41GkEmHdIrDFiWrxQUrpCZ3Ot8cHp4KBp7/iATrc09+Sw3phgLAdwkpLgIrvNalQ7l9
R64k+l9W9ZiwtEoeGxNcAfjUOilNAn8aRSN+GQ3ED8fQCipmQFnt7Ep1JEDdw/ljjOwCdHz78/+j
c+NsM5bjL1+r8kd15OCBP0ac5FotQ4x5U+qqjXa0qRSEn2daXay4Mc+neJOrS+2u58aJyQl0/lMe
nNqF9W5k3DE31+bQcLaKVSXudwzS3hcHPtDoYZ1OiacqJxa8g4YRGxEoj5wpMYQAKmcuYfaFtMVX
fcv6iugQQc5wjfJmqB4xvzsen7v4IH5/Bg25zFPjeRfaMsOb+ZIL1FTDYS0ImNrKoj29+Nzl44nM
R0mKluYQHR+UbUnCm/lZepSmF60rngsvNIgykHoT3n2qia3FMTalehiT+9t5cGW0DbmfcnBQUcFx
HeOm2GD15H52tJxcoKeiQXJNpwZf+iZFIAacX8t+IBjylUQc4MT7y/S1HpLw0HwvmIzIywIeD/ma
2fiXhjdLE4ln5gj01DvfO1l48syz6TzFRHlXc5mTVwQhfY5HDbDdkGnh9px8DHW2rUAPBbGTyILZ
bSJUjh4LSP/y32Vb8ejqt+fqFg+z5IPnnK1BJqgjDh1S77firdDjniU29Gy5RcCiTtvf6VOFLii6
p1K8IwjlKndGVjoyToYUY0MlDzx+L+Ewj5XJ7beJMQj/bxW+Mj5qLFOSoFh4dGZynjq56LAbt7nP
/0XESmpriOklQenywWZdIlbf4qQF1gwJ7ETuilqhLsq43roZA2bVb1DUbuw7A0RFLMpGAmj8B9CM
t3wSyiBxETxo8SYgrk532gfjUTlYzzqAOH1OKxYTwQYwSlw1m4TktLHczRU1o0WcMi6tULx6efgb
A4pgkRyVcdhWBlWXobqdyYiFMGknhGzNKHVaBnIdqamsjvLYrUmJjLOrBirQ3uc4W2CcoOQ+jlaA
9O6oQibom8Bq6+DF0D5+ZYnvgXPrgeQMtqsJJRfY0D999dnqsVpFBlfphWRZbj0pfallFYUVzMc4
Rxk/0yW+3+7TfBTTlXYOi/g5KxqeLTDXVW+nTeNEhF8hbhMGMoM2Oski4Trzpe50DP0qhgp0ofyz
Moi7L7rUb009UlXIilVmvZiSWYregEreUEMQZz9xxgc53Ryxg4uzORh/jgG7u0PIHgcSiYERxhHP
Ys1U8b4nFjmdGZ8RSPyF3D1F8kd3GYVFSwZiZ+4kjUsRp4zoojBfiydLWWcK7iGXVgwpzszidejI
/lzAOToIDBuDpNez0FT7SUBu+3gE0x+ZFt3iuz8MXz7jtmTSpBJKXIW9RbWMd87fQrzQ3hKBcVlE
AfYJA3HN8HDZBZJWBIIydLKi2udhc0JN1eIiX+7zsy6ceke1r+PO/yXONFSnnXeN8Ph3qKLnrx8F
/UkbFmL5EP/Hr6phIqtg6IyaVLAwkUwo36WPLGMakRmH4XOZkiFtIut8djd2Av7ZPGebAcjZEScC
dtHxc1NonesPiJnPCrLDFN5U6CV6B87aoorcwLG3FwpB6ncRZqMl7v+ZHBYpPwwaagwL1IxxuwUn
HYDt7q1kYx6glLP77etCtBDNoAUqzsA2Pd2rWFSXD4mAj7DQFd4KhOB+35Xuj4pB6sqfqZzv/KxK
dJlm+Fq054OProwYB6Ulae7a1N6oi1UwQVJQfyv/CkNrTgJrvP51CuI+Feq2iW1YujI6QINJ+GZ3
iIAJbnDtBIF4o7A8GgYkrkO0ocmeYxU0bF5zbKRDvLihaCrf4WFsiVvTpEmpAC/++doYCznPQ8zf
5a3///hu8ONoirALWaqrO07fBUY4MxGFYGTJpZ+o/b5P8TTLGgyICgX7Iqhn31z931WcB5TkDdbi
htVTHIh1Hu7YOXijj/t0z2/c7SxDrn5S8g8GhUxmeDm5As8RXgddEBeVhnQfI+efymorcqJyLY8x
Eyx3UuVB9BSqMGblA6hL3MQbJmGlenqzmQH4w9OkcTdB8kY5D2dnAVZkTbYny2zeUDRLHORYYNq7
Mm4m39EOGG/8sYCqzuJDOgTVCKGikF4ayg2sYJmPqyfj6dvt314H9uOfcOYvA13QGeEwwAw0AEX5
bUN+Z1cNiR6+OIK17/pCZS19IrHvx2M1EbpRYZ//O5tgODdrIVb6BbJ5PEtGR4L/K7iw5d83ljF6
Ieo0J3NrUVJ1hOLQixMIlJ95SN/+5+5Gl8PWU7zDHWSNUwifXZJnau80uz7NX9hmkjTReZquQuwt
41kB5+8wWCQRuHVtK3owFQ4W+XQK0DW4kr0ahMIk1/0/BHV6cckvZ2Qt8eznnVrMGfvYcXR5yse+
Cx5VZPtYUdruGJXLXebt/vTttL6/zbYPOwriM5bU9Jv5U/TjtsuTD8QRp/NUaUafyWfKbw1TKKSp
9ho73gVDV5d5I6jmM+tjppulGqEPSXIilW5B8qnz5VEuM6U5dXHwPf2m7EY/A3obvrbk0h8ol1jr
TmSs1VHTdZLxTYkmuhESsLBJbkVffYFJiLqBgk+FOTOt5nxoXyg7X4ywg8F155WnI6pK/nYeXnAf
O4bEna7k4TVp0uLuPLN2IpWPTlgS5LQTv8nkW74OPH419pBUAm5EF5k7J2EaRnjyX+LfoS4wWaw6
TIXq44ENyw6vW0K/ySx/gdyZQo4xAZtpM5/VDBVq+n7jycIsd1Svxqxok2DimRflt8qxW4rzQZKA
F6fxBAXYFMTLN48SvQqlxXUvXEPSh4+x8LvhAs3zmPk0eMzI1tQ057kYQDeXFH29o0KltqXydOGZ
STE15s28Eng1km/5W5hAgcovfJNZhPK32w4UB9zUfLakN3XERSQEIiHMj127921OW8E4eFF5xcxo
yDqQ5Ar+fMg1GfKnmdFfOrFl09nB6zKfesO60VPFmMiGbYzCH+pp7EuvzwbFUECmbWWmmva3JGad
ehNtcKPIAs2hSb2KEqOYbYz/igCaaKCua9tOjv6Iw/5ajtfYCvW6TlmqzGLyV4v0TEkCD3Y/2uyT
54xOYELD90FM60iFGl6mCRV/J0Bc611HjoQqoKj67Fdi7NycIG84Z1lM95TTTE2kvZVrbISFy3EZ
jgj4UuCtoDWUseCcxTqVdgoVzzREPqQ5I/6vv9aIhcMfRCcidMnyoU1e+uZORlJXcccUBme31bTh
zCP28XB93Cu1YJLMe4DHNCSH7yQZIUAADGigIpB5xaILxp4vk/Xv8pRXnpY0MoPrTHlJoYtws07X
JFDWTAfvHztJ4gfoQu/L5SQHbtk8qka7HkESUytMGVbuglwo2ijBO1cwBmz3+1qaY0xy40D/bagM
Qo+jXz9FQS0Bzefo8OnRFWiTJqj0xfVrmyoHIWCi/QvOarM0tiaKb1zSeBNwLVPNY8mqbSgoLI0q
nO8/y86D74YPQ5G9U1TX5p7M6XaZiOK4xf3aFeZMH4cOK6eJx4j7czZobKfQCzE4JXmsNKJXnWa5
WzHyjFIv2csrWRiShkTg2TX4mafT++9zbOfEecsijhQuIo6OsHt+Hzkp27SYVmld9znmVYIhDul4
UYAMx29K6HI+8i+KCz8tiB3mI2J0VsdwvKgFP9a6rbhYBX2NM7T2iHPQoSyexqcSaJjvCQqYoVIW
qgHY3nRqN15yUngkIf0mEqiJJ9J42kpz6uGFSSUXmSKs0dgE9d4nqg3HNuyMMU4MVsAGYfQ2Ff5c
OCituBnMmxJQdyMyvuOf0VdKE4QwZy2+iiAB+w1HuwZJCPew/jNd7fAvlHckKbzjj3NQWSATVMk2
+mU5FDUqCQ82iWTthIogkawsBLU+naSxlMXc22kv52/ZIa8XiKKXRFRDSCDw8iA9dX7i1lCVyW9Y
ge3EMiL+zuscd44aKZVcOxnwRnSvZXLJTNEIGf2lzdyRHFcrGe5YB1JXKO9AtfN8Ynm7pyTg5Pdx
FEgtECfkoFDDVWZ6pQFYox97Aq2zZL0ErZhco/0CX7qr91oWFzKV9eSQ4WkkB7S5K5xq7FFWNq/i
OBJb7cUQaoRttbNum1l90bd82fL0dRMBRVvkrbJr6e8F28JqwbP1/Hi0wodfTOK1TTXrxny8zMGa
9OXaHtxtcnN87ObTea0YWYEjfvWAm57JRvimPc9HM6G+527XBZ2tnhWXxzIRfCuB+7C67UxUDIK2
gC9OQEtXXWQfVGuWKXiZWOzGvOlWIF4b/n0J9nvnnDh61/nofdpq/pT9myaI/TJ4sTaIb4nc5Qo7
RrOO+2CTrCscGN9FRsWXepxfvwQofa4kjP+E6xuog/EqQ9TjDbroLUwshZQswqR4/BZmuESVonQY
CPFNSOsQWioa6x6feNhI0EJovEOwA1gnJTJ5a2eWiGHyzhhy7onPTyeM0ByjEnjG1uk01jYpP5ke
bo2TL/D8/yqnOYBggrfv1DPMFnMXIQ1ezQQgvV016sJn6a7wafP01MowmN3496FN/IYRrKhtmqOi
K5M9sL7AIX7tYZWFtHoEcMNHO18IKZzk/pV2PQHkkZlfXDoIE793U5kHSBhJpMgS9VYK8XzuKKRM
chWTHq896Z/OInCcvrt1uS1hHeyxJxwqqoFhrymNHn3c/l3fA7Pfuap6uBFBeku5JJc+kY6L/srs
30DQHtBaW6zj8OJhjRofsCcbP5cpGX0sPLwPFA5Twm06xF32/3JwZyHIrtO930RackZjmf7DsLA5
1N00GgMbo9j1fo+w+Y3mNNQkmXu8Rrr0+g5wr2fsD45huazuIq5jAbpPjczlJT5hb/sv8WGaLoiT
V4Hxoigr6kUQB7ga/KZn9pItQ2riFlgxerORrVzLHnr2naVOeAwFcf22lIW3Nz4GUAdFyP9j7AEG
xAVIB2hkXKQ13AQ965D9B6yzrdlpifNnrmodKuK91H7XjskgoC9nBR/b4WAIthM0d7xCTBS2K4IX
0ZANy+hy8ZbkPyAjRtqouAyxPizU+oY2XJYV0xQ8k5Zkpsk009N2J8IsNp+3vuxe/K3Gtn8fDDWU
hDUcwbn7SVYpaGQBs1eHZtSSzCu4ma56m3nggM+4HZ3erD3J+atKBg3xk7ioKlZlX8kXh7Rki9OK
6ffJb8ysncrHI5QWLeDbOa2BDaow/XpoaKZhImLtHdiPsJ0xoBAPaHrsn1pt3H86ZAlg8Rz1JD18
1jroroylsEcWS8Xwshs4fa0WZcWGBjLTC7UoaNpNl6077dTV/U481qxtja4co+s7rxtbAyEDu3yd
bNKA5xJjKsddVxOUf15kCSGUVgzBJZxnFiEky4hygEiq6ImJ7rYpAfx4gesWewywa2iZ+QeBJDnh
RDRfJnuyJ0Hm3/QGq+5o9/R1v2pUX3jD/W6BZef8ZEoXGDPZDJbHlhH3bh2EV0s2e/Jm1tWiUhP9
MTLeUQx72IodkYyqPwhK5Pp+sgLGioqUXYmUcS8sGuoC8cIG6ck8wWbHnPJVpR39msd68QyjUSad
ESUofIcUxvTHqMIWJ4UnP+bGutXoD5rsHA4A7j6bPsutUj7LcCWgqQ99zClkk/W72kczvKS8w97O
2UTyhKIVnaP0+RNjIpa47zMlt3NIjAMKBCPTt/HJRLLY/95rzLsw3QUPfg3IzT8AdLs+oj5LcKIo
owAPXMB88WSgJm7kXMX/nx9Uj2BOe7rc6LcDtnmyzRke6keMtRdqeUAVKZdtk67+XV+z7ic9MTyn
Ol+Cv3yNelxR2OQ+glaD6BibMkNOU1ur5DGDx2fu/VOT9id7yMyISzi17NC2KTwXKeUzUepyUcL1
fY2pcjcRaXqKfM1JyUi2VqAfiUkkeL3kZqEQvmXaQUHGi4NDdoISp9gqN+AM4Cnc4eGvg6j6/qtk
mKR5q5YPzn70nUuW+47JatUxB2sz1Dcvfl8MQYTtcrjlwEOar+7suhdUDbtN2SkdE3ECsZqj0SRv
Jw+WGeoxi2hjri7eDIWicwh/ljziekj7XJ7r1KmfoBSmjOHEZfFd71igi4GIpJYEwW+nPRJvDRdw
7jdeS7OPOKqbIafuIfiMwUEclIVjl80UQHAyWDw3w3J5YGM/OhzXDIcRiOj/lJEr4Qqfl8NVzlmW
tMv3fQshkfRo7q6fSg94sBQUj+YceAqx1fILjdEr1CvhSMshkCFF+Qa18j2rxyZE4YCh56MBnU9S
TmkC95AiGdp/v+h1c40ku7UDW3ssOlytcpCAoSGtFkmFI0E4lswDHmEuEqg5IPpffg3Kp7jq4gZD
K+luH8J5AAM4UXZXnfF6qynI0ytVuC4X7fzO8uKF9NbX71Kq10zBnVjb45feqsvSNOxzA8/OLxR3
VhyXjRyhPpYVaMfBAwVE26bZtRMmcnuUw2KIHsW2kRz33v8vA90pJ+2jFy26mdGDlm6epOyf7y7m
E5ndoJMHc2tsz/a11aOO6Y4+GbzxAQjPppRzbXtO4JahrTupr8LDXR/F3AjQo3DiUjk3pbv7894u
4EPM+R+PQd1xqPTRphLFK6RpBA+EG7Cdlcb38XVJe1clFAe3tX7L0mWjYm+dOtyby0kc6Rjg2upJ
aTq+fFe7GJcoHtu3/FZRIAopjp5JVKeDqkKvgxFj2oxGuYKnyzMFSbko86G7dWfWRNuq3JueRE1J
ylb3CzKZof4p8cs0XewBotMTJBnz/+l1mRGmmXJ60oRB7HsjKlgiRvISqqD5aR4OTuOSpxle7wPM
nfDuMKbCWhw8tfkYCNmGST5bMvXdL5Evhh9juuLB2yrqQLGciKJsLa9v3+PiFa5oDNb9P2zN00Ei
n03LbVLEpzSIUIk/GqP3+6a3nSGeqCB99lo8jiJByQcJLkKZDSC2Me0S8VYgmtKxSVyo9Y0Dsm/6
VxVD8ESTBcHWntWzOPKBy3LOe14ZXTacvCLQeE+VVu0M87vJPHeQICmzlDV0g6MDJVV6mp/ahoCY
R0gJjON4oZjjbZA1BxQUOYlV/xHPMmKk7kf5iARtz3saEojmxVbOCS3Zd4LktwlOcODH/ODIMVl4
PuZlqB6GHxJAcgTITTwkWlGdt1vqwGcOI6dMN37CsW0yIaUqJrWdIYY1YuUUafhRxLJ7jewF8fXW
5dnaxMkRQn6e3c/OcEzRkD7GG9fI3pKro9Jy7CWd5kmv3Bc3jplG2AuPm8RNBiXuo+Bk0TxXk9Ia
djHfoEGEFqqf38euG8alr0qTDdw6rSbe2bWdqAY75j187aXrDm5aOykURMyOgY9R/2HTDnGSE4XE
ypSEdNrolN58jew6xgqRhumml17we0+uUzl8N12zWhdvaKnoC7VZY1sBf2HUkYp2ua4dsMVH9ORh
y7gq2cU5HNhVwu2nbGQPxSORzLQcZ0Q/VZw4X7wKNrGE5ajehjZFFWkDd4TDMvNlBnJ4cNNxUeQT
GpXOAzlPgy3N9ppynJj9ya91kD+cM1OZTWCXuiNAgbdYWhkpXCQJrGDPM4eSoeBrZHuICM/lJh11
CWt+QZgxuQZJC8KT/SIXTxey9T6OTXZKmgtRIGmOpEHMbQ4P+kV+vUh/pUPj1kNp1ffGxSre4Vly
xA6JAYutw9mIzK2qjvS5bTzAKnxT6KS/+mH6q10nJz0JxOk3uKezE6mviyMMPtkxs/UIh7NHxROw
k4a84g7SjH8LxRF1GQlrskBtUWYCNnyKNcOC90KX0u4khgfamfcgSP2OkUhe3w9s8I2sCYPnz7dI
TN+l/vpqwamXLL1dFVSjJO+GKrmUOKfiwqW2MGmCyACphMvHv4TacjkjN4jx5uObeUV2/j5RzMIG
SCJLc6A88nKzndD8hNZC3nfR+ZtrNcC305EY3r1Pptt3HseYCh909Sm9KGAZoK86yV1K0beffCad
wQtZObyMz6xqpO1u8zoyJPBRbKsWcvPG3l8NS9wqGfCQCQG/LE0ns1y+BsTILadryazF8lpgdydS
IPoDi1nfvxvrySGl5EzNP3H4knhN5mG0jXeeDINybtcL3yO/ENu1lJQlsh84DsasnKY6WPI74wcs
fRLZsCBkWweCEJoAACi/l0w0VioF7PiDE39Jy0Wu753Z9SkpiN5d8pQ4ZPI7LEaTdHgaO0wahPW+
PjwuLWvp0PULsaXDK2nRvvB80F5IgkT67NpAI+k3Uqi8dqjXoN6Oxm7L2ODTf4tAxzV075OlIsHv
9rZDYqsaVV3MO+EOYVGKbfC6pMpONeNh3XnoatzdrwEIoCFvpNVpQjyMZloSoS1ruhWkX+gAVBLk
maqXtsjfhH455WSvqYTu5U7cPNOCRh7+39vaelf8Hbuj+jxmoHuQAJrA8sIgR3p1tvOJLz6lgOw3
BKDx133KiHVxeKcXKjz9izoOd6hnSNUVCI9oCnPpvqNRCwKkRS+MN6lPx5S/xuiYcdFfLPJBS4VV
g7UULsDp9udEAmZV6k04fzna0yzQcLnc6Ui74BXfJiGu1k2oRbWP3ODW7ewQ0XCOAMYy4BhcJs7G
h85SaSU0aRNFfTqJUakw6ALhWeHfyuEDWgj8i/+NTWYPMYJUj27sHKwrg1gwqMiHD8avktn98Y8G
9Gu+K5rOLiMd/I2MChke1Nem3wN29p8XyqsQbhUyPtW4I7yuuN00t+XfU4ExPp/l2eRiE6WNr8Gd
pPdvQhdIagCvvFad0v/WBwXcGw4RcEW3uR9SdknjjawkvDD3v/mbQ3k2PrJvJYiy4alD70ymRvGE
mmqhSWM9RYwfAPxQdoDoLL8HkrvAEZrWV+9TigocIOnRrcuo9WIyUH0TFgHGc5gvkpY/Wy/7BxS1
ow56/XJrSsAq1tNOqXIwm7pZ8KvOcK/PoTceYKf5vPKbI4HoS58BVZMbfkYHoL2DPr6DzXs6mgdX
Id+xFv1lFmDuyhuBhOMKVAGtWmeTOSIDdtuFBN8a0F3m5cfgU3kY5MpEA5x9ZW3NLvBNX7fK7Awt
UwKMs78x6Gb69drdhAARzKdACjys5o0cGRPxLNGdVGF1xXEYLZdnLwTOA1JtUg7kIkd1Lvn4QHt+
73Au2PdRbZQ/5KEdqtHJpaABbCYpFlBo1484x6avdDPehmmz3yb63x9ye6h6UacqwDPwqLTDkntV
0BP0tfVjiBpjGGS/3JxVkpEdOsbM97Tudy51aSLd5vT2D4zGHLzyjdpNiX0+3eFSeDke97ajHZ47
uRCZGb6kamA4JaW0AncPePixPAt6TQJRpDNB3TwOwUGObRji2mPy3DmNu7eDMKmHRAYb/I6LQChd
uFhF4xMNy9yVAJKsasVSx9bcHiKZwWJGxw+HYdFngVpWC7Df/8QQDHGGJI2kcdeNWPTUYaRYItxb
0dQrN8d8WC9txBtS+q04ieW8w0OIWBim4zEOpRc9qH5iEtUTVwP3xhB3sVIqV7JSRs1qjiOQ6b6i
mmwl7/F67GAQEdXTlsizbYNxeC1cab1paDQ522YkWwQNgTUmX3zR5kdjpf2Yuwjeoa4OgT1KDDS3
OlGyQVpuKdoQmp9rHtNEgy+3XWZ0aUJSwRcN1TFcX5QEJ3pnnt7xxZoSLTo9IUvkfZJ67wYRZjOm
7Mbnptixz9nAHFh029hGgBNkX2CQFtWYChrM8Kj/bA3biuKcW+O43TVudnQTJWq2XazCrTbYrG3R
bYsHTMoQPaFU+KJnixs0g+QdjIYvqaXI9je5fSw6bXcCnbf/QpPREC4oEnw3Vci+y1xb3fdZ8S8h
lQcO4kc/JczVez7EGvoXS+TkK4WQtLEzMwSO7zlxj0pJaRpqY+CsaHYteYZsEnCkSflIUkiAOi78
ZV4cQrqkXJ2tZH+FIepXgRcxrwxj45ZkwOORM/W7I0znCWQBCQ+ZAtgkN/sZTpAVb67u5knF1vUe
xQmJljUd92WL0fH/+AuFJHQLeVO6qTi0s4NbmYkQJy7pP88Cf9oHuJ/seEvoCDTcTkhlMLyQXBbz
aUZ5VqFbZJDGdUEaxjnnmx5VSPQdrMl6VwEL86jmv1LoWvUu50JF4/yv31dlWOvErFbG3tVjYhNx
Qd2VBjvJ0kGYHEqPDvrSVQY6BFtnebK4V057X0RxZKaGj9yfmguRcsR3ld4v76VLyy5WNH2hKmYH
/C+sU+S47ptRBU6QH3T5CvaznPvb7QfTs7zOkGOwkObCvgffEKmaP0yEaAiAJw3kcueZhbRlgffy
Y0XDkT7tEzSo8rLe93AIODcp/Zn/E/XlnTBm3Evcy8V8keego+GzHi7HPBdSEtu8kdB45pv1zBsq
XfStgi9lSrkKNpsufpBpiTfpfCB94PXZv003n1NfX42ARFP8p91mPH8rP9y9KHJwsv4Rdfg/WN1A
s4LHYmC5t8ZPZmNmSxbaXqMcpbKoSbYZtI8qXKsqXdRe9VksY38hWGW9RP/DkqCt/XiijplEvAj4
Im1qhZMRyxnZhNI+cfoMtma1ToPXf+yi4ZloQZrh18FQDSwG8NrW1JstCeBLFxLX3axA2tzgmtzy
SvJLE8K+DfpuoYkXgnh7V93J3ssmHRe0bY3m9GQtxKVivClFFCLsUeIMcUgiknQ1Df9ocxgNWTvG
e0SZbgFMk/9m8r67dbEdmQAtedVj6RwTjt8Iu/KQPGB58ysw4XwzUh9BSCUjONRMz7WGMaq1aHGx
MpYvNfLvEdk1wXnfNQ0K+FZzzVlFc8yOu/K4ljMFnrF3U38AsaoZXe+Ose5iwmSpQeersr/+NQlh
pyN4GjMhaVetTPM/LTUT2+jqww9y4SDOEksbQhh5COWuofjKwAfYaUtqK9/zC9CYyoxAI87ysbB5
zwYR+IX5iL0NqPss7v7zzp47gVSi5zppdlEmsoPdl+qMwubXg93fu8jW1/nyS0vA4R3/K70vBpl9
kl9hE2fOxVfYEk/vOL0ly3yc5TFnBn10rdYzeWY0/0cn1S+FpRAMK3gsBe2nzznAL3TayUy7RxOA
xzAM+Xob8n6X7kTfEycTf1O9XwUWGNOdn0Xb3Ml/M0aQcwau7Au305ruRtQbQkGI/he17GM1LM82
j1KAVoWs3HwL26qTLizFsRTPP17BFlMvgX6v5eV3HsR+xROwa6BUqW0RYhJo9NKXt+XGsBDRGwTA
tLmF6LOmM2cZDtQ3nBYVb83lnSVnc+C2DD1Y71Q4TVZU3HzOpnxzC8mHLJ2SO3mbEDdHFgwkVtsv
9mw64619IQ9oJSeG68YLf67Za/XhatspgZEYdgVUawtUOPpL2Xj3iUakiGftMQt2G6XWNst8ITSP
0oYsXrDeFv1OXAOSrrNr/GDAkLgUMCbQYZFvXJN/yY2IKS9jFmtySQV0FaBMwTpE2bKFlSAmJh5+
5EEsG0lVRp9TOjpR+kTDB3o7MeD5KGMXTYcpuThzKsMN0lJQmsQ82hv/uPyscUiDeIbxSgnmBFw+
YUxzk7apJlqDSGpyKRhWpyj+aAFaZtEL6KGvQONdZsuZ9W/JwezLhSZoe0ZrrceHJP9KbEjPNLYn
mzcKn2eJcqCSKzNOGakfyFyaFOzXYWvx3jxobxhAXKMVv8gdlXqj2lmzZaykFuCgal3nB01z7sIz
mhRf5OJI7ES7t1jpBKQK0bcht0+Q1Gw7K+3InEbYOgRMmbXuSi7TCWBDKzeEbCz5LlminFC8fXhE
ehr5f3OVEFBHOD8ulpONxkph5+80lEKx57NeAuC3h3iYQCPmYs0DCo2nQM8fJzQdYnFLS6/b/81v
HsU1wj8JjAXDie6KCqO1sZfPWPvg+y0qz5Q+948txGWicv5QtaclROBwBFUzn/L7p0uZ//e4Iy0V
EkSaur7ib6XyquNeCjZ5zDIIq8U3ndta3LUEHlt0NY38W0CmjwuSR9ojH7Ba7QNoA0q+OuM9OGYU
6oHsOdGv1HZrnoD5aYX2cj8YPkgzVTItmNEwbFBfCemUcZpDMs6YoeBSwK1wMScT4ZEH6WaqCLAF
7VxtYS86sZ5oJP7u2Td1lFenEPcyHLTIFAJPc+ijDtY2iDVErOXiOmsuxoaiJjuAQ1iKyDtX7rDe
lV/1z+PbXHNpocG/Ndk8wSux2xzcaesO3/QfXWkeOiSipUWvpdIJ/JPYo+RrB6ZnhEBXI6t/OVfl
Djiev0T+YkvJRkpmSXSXqrEjYBZHay1YYOKzUtD8UwFVE7iaqhPNZqK6OK5JPz1xO9TH35DGn7Qe
fCWzJEWBrdYLKX1139PuhdnT7p174iA4ZKKfHy6Zu3McYnmx6XRNbsnvXlWGrtIMVKc/FA/gK1WV
sLON8C/JVtaiA/J1/EXfj6+Byf3jjblzw+FFqWoL/DcaRxkTwqt2klOkvfkyeAt2P/9Bmg3ZVVIx
YAWxWlRUVGZdSjBBqBgzEGsGzZisuMFt/4u6cf4JTjL+PQLs6MF4ndh8aZ515ui6+sLKuQRIvLp9
Vfv1R0z1KNWxo80tj+EoEPHrTO8mVa5ix8h5d51TGok07Df7V7Ey/Peg+r5dceqN2Kys35jckiBP
uUOxIeNPgBq87Tac/y2BTxLa0ly6LfsrFYBAYG/MtPf2iYuTZZzhiDG35xrdPFC+H/T76L4IxDjR
a3rPvhvuHoeoHsPIeBGhBICrq9aAgjbGdkBF9dXcZp5sC46rzyx60A60UopGa7rHc6N/b/B2Q2WG
aRqeNtqKT6fGSjNbot/8n1BaHlsAe4eQ9sWplFQb6cWsnKhVVVE9GnAWGaq7ZtaQI8yibiHMRWwA
XqLAllERMoM7aOdvDQ0ykJn3iknkKvjPJJRJkgYda8Uij9N//on3EmUjO7hAEa0DQb2ntmmCf6a/
N84iYuT4rHH5ZAGbQhrUwTBKpyJMgwzBZPKq/MJkZQgN6u4Z8KFb/X/+Td93cSrFyGubqxiqHevF
o1H7yG65hwFb91DaG8z4OYNtIZlsaWgrRXjuor75AwWv5mNNFZvZpy12H82qpeQjWFC+GAtYYbvN
URUaqlIb86yibY/XRQR9WK4UXGM6pci29bGHMZ/fsY9vUauA90Do1aS6jSzjRQ99rrniEmkNcqo0
X+QKLqQJj29ArP+gbm3aim4/m3P6kO00UNPTqJFe+d4uuboClSjBhdRcYzrf42ssFfF4pZAfGOPp
vkxBNCQW636tD9sQeroplPCBwYX2DFlCAgzkjrsw9+4vdHFtN5gswHpGUgUsBh+gW/HLyetjsWxM
3vXzcmE1fKHGbObz9q66qLWp9pSfRq83aBSRMRHPlxhwK5GxES5DkR55BM0rACPUoE7buP9677WL
qo1+iWdzI/usF7xvgEGQmr4j9MHrzsa3WgANYblOsOK4cN6Myir9TwaU8mHEfs9Hnj/H/BfNakRR
maWw3/6geuTH6uJ4xa4qIGDI/rFHip19G/jZPscJ8ZwGp0H3g46SFjN4atUTQILod5ATVriPlHRZ
lBWJfIAvOuc41EIimCKoDwpG+arNttQaB+MDSzeWNvS0UBj910CefEi5otRppVjm769KAIYELUik
S1NnPtD01021UEIiGhGNJ++mprHI7j+C483dxJwryKGxsmGE1p0O6xLdpntFPwND4rv1uHczJsaC
UsphawpfZYVKfvVzD+8r6nfcyyJ570CmIaGzenkkCeIZCOgNn5uEs3fcwKIGdk6ma7uTnkXdClLj
NppktOyjK57tturzexbqnCIW3lXK9UqdGOB6RxnI+xjKK2aLwg5xJIqmC2F5yIqAMif1p/B39HgA
lL/25buB5KM3qEgz7EfdAEV9YWqwTEXSbExew7vggx64dKrCiB7JWyo8QKxg9TMEa2Z9iJeF/y+k
1li90PfwxqqQ5CkN6/dp/MuEvB6qXQXz90oJRGIESUAb6UoDa6Z8MuqojN+i24M0Bm7I5b09cia0
Jsq72E0rzV56L1O5DSf+9z7edByNT6Jk2RhVdx6TXD58gjsrg0ufwdlPXLkEdIhpJ4uP3KgSvO28
X8NUfSb7MU98ghMsy/IgoTvginCpoUuZsdpjSHbnIODYQIULEG2JFSuBkAFuHcKRDqF4m98Z2IIX
wJ6h7VvuLwquK3hKv3/izE0oA7ctXNJJqSU9yqIbkADfkAfuUD977yJZAxWnbKqeH6vPFyAjPfr/
2l4C/mf6ZxpYGjruyAXKuzgtCUJgO+2mbvl75Zj42m+frlkMskvD36J9BXsSgjllfVxfJlba6Oae
Z7N6KB/wMk7mMIXD8FILyRca5d+e1dDoIBgckoTH2Cs6GKpN5NPpjyOY90RUTcIbMHHjAFMMuPrJ
o2dkNPhdySEbG/p9ByvgH+PNPpwL5Gzlemh7j4jFKbFthjefjqyYcYDhSahbkr2r8eLaRPtUWVPI
imlhBiw+vrEGbCm/iaehdt31nfiM4e9DDQ16jrZ12E217jTFIbxxTKERWipFHYoHBp0H2HTb8L7m
oZa9k9Zntt6RnRWX/wYN4H2Cjp2C2W48uD4HJcLnrVlIDbwLbjKKJS32rdzoTkZLMEezxgTBVz8Q
Byqk2+SkgpXrvmER80MdBmI4WuNt04aMg5QKW9+KP0YVlRajpWWG0ZIyBNmIaNJFfdkLch1aV7ho
SKLbIbBzKPvLl5i2aoPF36Ac40xgTxbiDpUHzpuVTTRcLSMd3RPeHHT7XWs8gvlGNypsbSEFAQJm
uGf6lzLanOh85lLTQ69X6SDVCw3qrRoMyjH0LwUIuxBYY9CUWoc8SHvzxP69P2kZDK/k3FTl8Sqz
Bc2lySfsOlDcZ4/0MaD0C5SG0UpzgnNcADipWxH5C58UQcsqogkFfZLg+hC/chSYxIjS1eJPJpow
k+v8GmN7s/Yhk4YmBcly2wta3Msc0rt/+ucOEHiOWYt8GyYkp1ZhSDnZYhlTagtK5ai64opQvtF0
sbunsVNTcxfcDGYDo2XCgVj8hr42S34kBx9hm2WKQy/aezBS2yz9BC+d8lSxTcDUjjsHKRvTekf2
p/7ZgMa2XSNDeI+rp339QSBqeaVOchMCWYpgeWQP3YHTXDGpVYaQp3Tsmh+Yebh5DsXFCsHclaG1
w6Mt4nXdM584ML8b5YsjQygp3e2+YXDtCdatLvQjpNNccFSH8jMlyDFTi8GgSwGQ6TRYYaqEIxPA
8U1ngpKj5F5LAseOGLUdqmVy9SdM+mpNovCqOl385EdFFQtP08B5+Zf22AcpuD78Jq7dwaicTgj5
4RNeVkvCuXZFuDIl3k0IOOn3KpJSCRDlemxSr6oCvvfiGkzLIYI94Xv9HNocYR+bQsGrl6SCyg29
q2ONvwNWtfNd/lAo0h/jzZVJidxusDgiw7Y07igS7LKRd6I12z1jf/pQchoXD2o+SOG44cdGA8K6
wRV9AQ8NKvUWm77rAKtCCrncxhf6N9q/C3lGIAWCoLi3rnimT6+UlPz1RTFy6rAFgUzy8TgsI08/
52h+j/vwtKRqwz/J/sGogv/nigyRRCipaPyfR2jtoFVcAXkuQCUlJAoFx0pvJ3Cm32MjeHgigkTB
f0nRPMeRxTgmoEYPJU+Uyl1QPVVGujb4NcOsJwv6ZmUTEpu1Zwns8dna9G/9uvA4DkZwPh8wYEnR
1eowyaZWxQ8YgM0gX8OiNkONazfDSUw7C+ESBd1ILGXUhQFKsU3DRB/6xxM9ZNMG9zFxM70Bo6IN
u8Hbs/lYNwPybpB6cI+EO2TJPSVmO9o0gfqv77qkREzDUkO4Sz7qguLlfgvMezCiUegpQdFAR07L
4QxkCXBRpNruxFwxLF3yJj99H0lE4kbnAdjAayb2izy9spY2oe7eIEVWVQTbmwhVWsYnWDs3No0A
OtZn0KSsC25y24aUTofeLzpHmUoOPT1lfwl0l6KWZjRivByxmO48heotltoSelERJxB/WrefgvUX
dQfmrTZCTNycnTcqNGoyxKmoSliCyYt174CSX4l4IziFxNA6YKRIAviuFw4fy31I/yUWiMvAip76
q4YvrJtBWk5R0xsZrhN2CNZ8ZoCLt6ow8QNr5sU1O2obSDVgTHmQOjmSQaNnpC+R4HDs0k9iLW94
+pSJwwPKk+o0idLZet8P4gQ8G4o9bfWSMBR7Ck7xiwkcOqjKdg+qjq+4Gp5+p5BVDzD8+mi6/zzz
W07u9wLhsTgQ0f6NueMNpbyILcMLjPA8SZAFxMNPoUlA13NlPvRXIvVHoEr8ZpPJzDE1427urkPj
JPi181nVDyy8hSoDYFUV8dCzXh0AIRXdtmvuU14Zdj7j5Y3EHzv5F/+HC+HCvZcM9SkdFuyatC08
ARNU7M7zbvG0+0uzopxjWRQLod3BPbnx0hcchjk3GIfl3pIc4kvSBEJxBerQzCVIS3crSZnTeTY9
TytDXpNGDMxtmlzbTFQ/Gjl4FXkvOuFhJs22Lx4Ilv4V18qdjYZYVdVVcbVOkcSdzs3wqjAJkArM
A2UWYsZ9iLT+zRQFB+is1GcYgrac7TbHFLO5hdqhe12dQ0voImedwX5OzZTkMaZtOdDP81P3Cj2q
Th4NvyA0kMbvgqVVjms47kc1ah86gwBPB2XYtrzRVktqGPZFQkZklxWkTXylLUnIIVMWnl8uZO5I
klyTaq7LYlFPzfRb6GLnS7GmVAlDGvV1FPgANEcaizcjPiz53GyFJSzdPM9TtNwm3KRXMmZgl8BH
qkwWYj3K38QMAxPbT7Ax7+sy7ln5qiQgCgdaG/g2PMvm3CMOGN/uGXs83bWZ7uMuW6dc9RUdugbU
ut378zH1ftkKIuPyO2ep48qeDe6Ur2O8rYQr0S450FL3amHPalRCrgjozSsJ7sUdq9oAOQJxUAwx
1GrNS8vz03mlS1H0W+PnNSw561fKxW/6Udl7ED94zt3csPtjTxAwfB8ZuXEQdRe1SOZQxwuDXZ1v
vpm/o9uKuuj0HJSXsGKsceqwQvvTotPh6OH0GYetCNs3VuOx4+pckb23tuLuoyfJspYF36WXHwKH
iyJp9Fj5D2deOc/GcUQ/DSEe0ztxqFGaTKr+r51bhEuAoQP2oVBjcXuS179+NybB7s/uylsOeZ0w
dtkpu3IGSLH+l8Zfagi+o7jxEKXDmmV84Zn/gzzJZ9e2LMfnDu7owDHPdHRIKoWmUZADyWR5aEzh
+EjOOFWymo3Esrl5zfEjTpH0hYVKohxeNcRScq1kAAVLTxmzTGv9qKrnaz0TfbxsGbuBSbTbmtBo
9PHCgacEuKmaVhONsqANj6Mk1W/l0vQ+02/clwQLuUhD7lshgXNTE2DDbiZz4GXPezH+3+9gfIIo
YWkHdu9AalsKoN9QSIdzM/HyUF4ikJCJKM+6i98ov+EnHVHEABREIwEm+D+10Y9fg5TUxtnWJl1q
HDLqaRMueYYyDGtDOzbouadES/20OCYN0VO+JLjpNrdGrX7aUwJGZMdnajAEjq4cGIeTX+C33mNl
9gSkVMKtYakhP7vyfFeEtW4tEpTRyweBcpFeMtk05fXSjkV9YYUZPjsfXEDQZ9a026MoA2+qxbZ4
Pt6HBik+oxa0B5SDPQ0pT8TVv+qUTCeZHbRwt585SMUivtQsH1PxMOlGvedLQMOxnavks37CuaDx
s1nrD03hv2B/IE0Ax9HsHF6ZZHssT7bb53UYbsjAfn9Gp8rwgDDl8Vw/8unYIeXRRqA4YikYVU5a
xooMdIxywmuSYG8DBfhrUZ7bzvSb4Yk52va2ROxEtuBWSi3Bx6ODyQ1SX6nYCSa3t45p2zaYcHH6
6LVLqoNTT/RxUwZfo+6fnv9Hf+URqRekC4abbh8zwB7HP/OZ5huD+ImS3V0lyRyySJYZEm9Evuni
zUsUmbp7hVXE0jcmPUvjXbcR6K1flqjnmEUvNrmFvLQzXnrmlM0ypvfHALRo7Cz2F93ZLEXaYReK
o48z+DEuRqBf7InZVyAU0XGZwXwwBURGhcsFMQaDLbis/dWdq/3xrc0E3E/NFgkmzazyfx2qBD59
ZhRh06TmOJGJ2Z2kMRJPvnhivfmEKb1PEeDVOvIXwrm7+KTv0LRUOUlHfSGKNgqSaXthl+I9s1ym
DL5kFtOZKfrCrQknAnXxgSxfVPw1mK9Y9FRyL3Kb9EskqbPwmXgGzkQsEXVSt9AJRwhC5ZIuljm2
7VA6GMJIfqDHKAsFf0eo9t+E6XDeo3vrg/72gx8ADKLKfQvGjqZGQt8PJqCpSBto8PAM8nCJDFR/
TgFDQQ699joGpq2+jEuONPbs6EnnsoFWBygwROv5QetQ6udLWkbsxPDxcIkntu9RruMOne0r3J0R
1Mh95uyAdyO9KtlnHFBYHTmS2ar8CwASOIe+ImCtRHW+u3mDaaEIziRrHcQ3lFHh8vJqvCbGqGqL
/xCKRPk9IF9H2Kq0aPQnWWk93CIH2A5j0H+e5ewUPzi863mhfUeoOCdckNVtiuU2JNFmIozTFLJo
zOstL08LnZWi9xg1JK3sLwpyw2TPpYFFuNP5Gw/tyPhVaLWpiij3IBp82o67tPg+meW+wGXSLSV6
L2EOr65pUikesm6w4rqiBQcY12owsPfCEFw8uG2XeC729aQC8yWtdsKb1XuxyK65QdOsqrwmWW3W
Fo7VWvYgSZ/Z1jcQuM8Mxev9pm2V98pmqeF/Fsl/bn3sF7ItZT3rrsiM+ZEIGlo/crba3C0KCcR1
S70RrWIxJo20u3BVkE3wB7I0IrbXLT5zOtcvWDV87zlD5uJq4ZIC/+IDKggbptDDctkflNXIkCZ9
yZt4Lb2H9NcZ4sabTyO7b7lrgjddWliRv6sakpGpQpPvAaR6XGJBMIzSFBgDDlI6QufI/33guc5a
EHvSD9mCURlyxHR6MVBDsWDh+CHWafFtTjDI8inLVDJYkl2B5sRe8FV1wDCx3foTj+wnotna5sZ/
4ivzSagzBmXyMzVuIa42docaiHn61PModqW/O32y5mnTmjDmb5NnsnX8TPvbWnoW2ytgAnrrb2ty
u3Ov4cgrcfFAaJanjsQ+F2ST7FFdhQN63nxv7vCZGaBLQcjwmT2Wrj2rOJMFzZjH/XGDvo3Zb25v
bXAlTvLa+sXo4KjKsIoqr7SiTTV4wDLMJGy4jMfWg+vXX+020wTaI69X2bBlblWmw5m9HRdfsxgJ
3SqLO4uJKzlFNiYhPGnHHdlnzsCssqOJtoF85nJLJm+4/y7alQdPj5U2oAXagnQreUbXGKf9wtLz
SJCp96ml0KMg5DilB5VFad/o+OSronIykdExuzNaCWjqs9wGgHUlQtrqLlFtHsi1x0Uox55FpNFS
sv8FEhjvW2O7AzoGf3dztzbJx6cii1zzIENPjhGb5OPY5+oG3tD5RBwl1VEYospqMr8ypqXHGq5q
sbHfcOLv+La/tIueAqpu+pZ4gBLEwroImawZ5KV0zuL+LqogD38XdHVCqs7jI3vvFSFyActyYe/B
5jbMRgZzdCCJeMk8NkNsL7LaZOGXMvxqa31qiYFf82Hbs+raivUKLjvE4Vt5V8fyi+ZJ+eqbzmu7
fAmhhhFY1KlM9HNhAG+jWkVWfk5oMwEQJh1gx6jWLTJysDVpL9/9+JUl5lkPJGGDRt8YUFsQ1VW5
LahAsg7f+HivFzDsYPUJW89ZrMMQ9PIWz4ezi+b4cbrXTlJcsKXEk2gPElqu3f72qLreKgY4pHkl
bisTySJ7Hg/MGx160KQwhgrsGPpdDSJjrRXggS6/JvzBrUK5Yr8uyBCn0Jro021vRAgU1JG5f2jo
5Eysc0N+ACaBnka5azMUakR1j04h2Kekx9b4WROlbSkSwDagSYnkr7BnG31hK1LhYaN+lrjqaMRt
M7mYwK+J5ke8YB1GvyFnUufy+n11NHIbAAabIW2qj5FHW/+Prz3pOPDsjKFrAdiJTTZwCV928XVz
tW9SJa9xsaa/jTpaTR2c3AS4U/sk+RA7PFBKT8w0gUx+tc7sZhjB0sNrPXA+uNpZ/Cpd0sPzQoW1
XR+eShYUlf3QrAkJEN7keW/URxlhseTQWyF6WNnhQpV+xY3g/d1KfK8OGTLRlvXTNjxKBMBclhxu
HZCLwISCoDd1XhpLlKMNSlrfLZRgftb78JjEGfNPnbcMDOpMZQ3kPMyaJn+He69GLsuUe3idX86m
tvrU7nlM0yC1vkOcjnQi/BWqO8xrR00UVswyCiTXTTuKhvsc6WUjLTC4VD61jXqcNIoBfxZ/wUuo
hMdv5beRhHhlbtZTQdFUY4bjZdfc9M+dn+rBTkxefKrzqTXcqQkiGvxG2r+MiVolb0bGPSVseAlF
hg3dbtWY9cNXWWDaQA/c+j6kMhFpQON+ClniKMWEgmaGGZ4Uqyph/Z4BaW1mWGHpP61bmeGPFzSL
yDVg6ISO1NSfbb+a/B/SzFacIevgfIhQe6D8NlJ4PmiYBKw48V6klj75HJoccLl3e+YMqQAWdUt0
IAnobQgi2X5R5eqFJfsbPFKdbFRNrG3rJfBFBBjrZk+1ufSV9oQ1pLPDfyli6/Am97u6vM9/6EDu
Y60juwQquYzruAGlKWbVvNiU6oo7i9WA08oX8wtaThZ6CFTwOkcjhJUs9yI2iUjXgjCpWDP93pNo
JWI9SMaf3exswVYq47gOvV9iPHNcFg6YVVLFab04IApORZLI3vnXFIeSiQ8kXQ1EMnAIO2gRzapP
1r4gGTt5TLQ7pkNAROJMWo1c0TI6DP2ksxHJkJ7vXpeH9jK/NhnBfxx/CsxYOVDCP2NKTVi9zhDf
J1Lhby4axZhWZDRfaj41tvVH8oORLLlSbrVX1XtHm3hlZCQ5FzzlZg+8JmnzOH757eXsFYCpgIxw
h0gIwfXq/BXpsvzafjFVAtAwPXBVRNYXDKQKyi1gu9buYYzrnH2kU3BX19RvcwHICsNMnTSPqgX6
nAuA6udpyG3daFNUnph4msrp3h76R4FZvHvcU3T3i6coKQnkIUdYI7hYGjM7nTDFa/WnVrXRRs4I
GgIuKuYzbeSKiI7NShZGTnN9WQ5quoBTKO7Uk8ihN9Ox3yFpO1V1O5pIsCqydJZs7LlvuLtKoopD
KtmgUGkj3YJwfQTYHLx1Xx2OGwLko+QG1kUVIeBAqFTXArU4WeXSfKWy2mIUi58NtKMALzLzbvuv
00AtEbOLlGnJZnEJo4mTdQf9ya6Rx2bvkC5BqHOdrNzAPK2TIaLixnTX6Xn0eADQAnvIcdwaGSet
RoyDjO0loR+HoU7kKB5Iu6JKyyLPBQqOJx4NLu+ZGAMPYGTysxc6xb+NeXBn+3p3duQ4ge4r6iue
2jy6QthFR+noRO2aiVVWCwKeg56Av/i/D6dcFoE2xOR5SRo1T0bWY99gKrRVGUoN4tA70/FUq9ff
o7G/5MBwGcxWt5mIWmX3qkP7yGkDfDXFtYTnjG3BGa8lgc7a2115d04okPvbxhgI5XpOzeEHQzKu
L81pvUCVF6Rj+V+rVOYcHD8DNenPJE/LC6WUlx77pIeVHwebp7TO4vXBOn8M+5ITraee1zStEtVv
dT5Nrn+eWyibhwlFWFzG3EzaBX4EEMbZxQ6RAIEMKul7TcZJQxXzKo7iEcw7vtcrBkjw+8GdiKsh
yFot1kN7inDAHvyvy+xRuOyTSdiOvXNwqhjIF+rmUbCHXgtZiHqDEAqPfAjRdZgqA9fOwDl72zp5
WYiUK1W0FhrPAKoNRfKGQaQpD2VL8C9fheTOoUBiNerlC/5Pc26tAdoJnuEU88aD9+znA8DVv1pZ
oM9i4wjzp0CbOHx+HDFkJeiRMraT1q3UxBElME22fm754awm6DBQF8A1DE00V1sUEUj1bLmWB1jo
XLEDSn61EkTH+IfKrKg9+tyH5w8xmMBBachJ2ya/RmPJUhsYN76Mu4jGL/4QJBvOVqFqMEpvveRq
foUJN178FQtXl7jMsRQV+sq1adccxM6xW5e2REw/UOjX2xS73JYMSob8QNGF/7uYvNJ5fwSu0dqk
KX8Xw3DA4m0f31caAUsRcLumFhDwMlQV8zwFV2TrSIotUQ/ohuwym0EPk44h3ZWZxd5qfkEhMD4t
i2KCvm7Swm5YWl4QK3SyMRoGWCXn5YKH4zjipcCZoBz2n1meBpHjsSBu08NTpV0JQYaaDq7nZNsq
OaIH9IfPkWTsWfmMSiFz0EGORk1CNA5uoNw3JP8qpA6HGsERBtiWs+rYn4psFNdzEIrGEfAWJLoa
m1x0FJWRSWNFjO8szUbcJOrEpXM4CLlUba9c47kR6AnHxZpFemUyttfMNOmWp46X5wyQRroIoevW
Cdt6OTyqKEG3UiX9YFbe1FtzsFQWzyCFY0jaZNfLU7FnlsEMyxGhh2DJo57J3EJA3s1HPug8gmLn
i/Uk/0fSZsdHz8kvTyyRkx60XLVdfuxiJuMD69x2SZCRLzjR7rGUMEOoOLATdT2sGLKJpBL2sh8g
xtY1KPBJN412JvpHrNcUVpdPL/f0VJ/opMC14ZdUDaQh3je9l2+wGltnXuJaGZtURTGCpjUxSDJD
8yTUakAVcZws90Ge60egNlJYbME5nDvnxrJCSh7zLJ2zYBPDYfw0BRdrZYenyexw+BUvVOrnZMYJ
pSKvR56nmxjZ2Kl5UJp7Dwxy1GFRv+/eT8yWXi0wDUwMqYFXZR4hk59eWHCZXu8c1nd5P318W+s7
kd7eBI2dMPow0+07VQDEPKpfaxpd6hmKSXwUjFN6xSCVkEROZtvS+D9riLFz91p6rACFbjXPNl/p
6V7IYSOVXt/6yRdeXsW9wGaYyVm6p72hL4O60m8WBKN5GpP6HMRsJwGMHwN0+j9Ia/8iFjBPEc49
aNkzr5Nvrc1KbF8insJTTh12PgTfotlNEdG6LuNgB31bUdA4ukWuY46Rh6PYOJ+OU7ArpIjVUOGu
1ywtzkXLyBXU+LHY4l4O3lbHqjlBYXpJ4KJpfdBciDMzpQZJ7irkClDe3xP/hSyf7q1iLPs6ZvAx
eD97+p9EAt0QD0GoefTnOYYLk1ZaCn08jFUDAVzcbV1/6Cxtc7W0F8adOYr8XHreZymAcmlJ25Qy
lC4PAaGRK4iyvN11Sc9ZsAF171ENvtYi6DkboB/h4745YLGsj1sU2Hrox6YtuklWmvWBNAJNp1DI
qYAX9B00aHlz6hqgEv2IJgbLUGox73XZgjk0ybsceKVT4rhgRUKaAXekv6jCqaxKh37ShZXsctGG
U2vu+aSlVlHsxYBmrDSCpszqw3/6rAHZuRUlbLPF4Ft4ecCKXTTv6R0BF/FfXisfMet/ekGUFXg/
E2LZ0FP9MT+8VK/VAielb9vBuOoUFq/PNE2SP9u1/1cp/m0KImF2vf92x1eF24iX7jqafDVDHRMf
vljoXoUPe+3Voz2AHM95kEqdY//3D1nBDd3+LPeLkurW07S8NHm87o4Ql04qR2bHdmHvzYcOTNAC
eSvlSt7bti1uVGtzERhdu+yeTirk1yHm/UWygtqtTyJ8QJSFj3S0CwLmqs7AMvTiVIdUSZI8Et8B
SPYTaHWs9yBCAWxThXaKtZDnvaYyKq76dq4ONAqmd2suhinJyb2PpV8HOOH9aAF8MlM9bvCPT24J
yhudxNvl2OK47I+57gsyCeOmHjeXXOjReAARG8azQIPUCAgcqEZHEIb+hmay4Mv0ElRlvHlvzwTi
314tpChKGqA/SszMyZOUHPlRORulOYgLQSMENJVQCAQmV4n99TsTqC6hwBVcITMXFobriZ9lvcs+
8ZT+VUDdE9/e6bkjx/HMrbF8B8eeodmkoOCh72UW/Ue6+oB7ONkqQvvFvgFAHGT6hgEzQ2kYt3zv
TEs6veWd209y9v3/u7D+0J8sPTwpLatNUZx/H1m01PfiOojiwwFG8Gp1BHIiUbzdRdmn0hlT7+A9
2XFcUXfc2p07bpKXo9Ep0Lb7P50VrXNqAsfOJKWH9XZY9ZliKxih7RfhwmbLnLoKrU9v/6yzLuQV
FNA64yHOFfCyKMAnfEwhpBDr5lARk3rkDFwcvg64XG0KLbIxv/m7NohbmCmIDCnr0JbeZp1ggXPt
HmXAR1rSXPim+rn8GznOaGEYp32Y+Ow1ClqiXUWbSikiv02ep37iTQ1HaWBQS9Be54Q0mY4iPmH6
2Om/6yy1m3FIIVhMqJ6UoLu2G0HDSJhUQB5MzhwHOep7T+QkpwB2peX5PgIbdvoSJV0lxUxCKcIE
19H4V6ddOcBkGFAMohBU5DIWIs+n+YYvw7j12uk4pGXG7mhRjnOkJLroV8kN1Bptix1aQqbmAi15
BNQpKCVVZ8dfXtcxo3hx2P+pUQEvGidncQ4Wgp+6YB79I6kSc01KJEIcu4PyZU2ilqAnoEg/z0FF
ys7nwnHSnaXmIKDbEmvXa1v1+VH+JKCLiH5fAKKk7ZieKXjpjPOK7SP2vjTbRSIbem/OR667c7mL
9TB6I7fY9+eyo63pALsjFeQ6owah4JhaOcevHcFh+JPghHDXugDJkXViUg46ysmXaSnhZRXS+44I
a4iTWfvi2MPwyvbtX/WVT/nc+XMm+oxsH19ptgQEmyzIOII/SjVNAW0tDEgoeZEfS9gY8EMJVPLd
Stb4ATqG8tCnGZZas6y9M/l6pGYorw9kBn7xZNTTuCZTJ7vO21p9bL9u1MtNIsgvcxRQGMfxgNfU
xCwe7N7+vpRlA8Sr1MOz9cvCqAYFMACpem39d/oN3DUH0FCOoaF+PPW7crusivDJPdJyWe0eT5XN
tPjPrF9Ar1IXWHiFJgSzROcmeEDfO4/pyH5TCArB6xPpI7+tWMUAZthNbzUfla7lJm+9+6bVjlcd
m37ifyVKtXJjufKT1QP9JooWvDJ2bdsA7zG5aqgxZF8bgR6SEXZZw7f2O9vjqkyBHnWo2FV+aNQ4
OU8DKh+rUHtwJhhpivrggCJxZRCNxxfA+r+aEg9B8bvdOd+mzd947Z9lkNvw9KwQyFmekB0QdTuy
Klzf40udUfY3LxEb20ZGv4Vba41xVNHKyH68M2/gbO3QX3GNUBcULzArmUHd2arWUXFaQxZTRQOH
8gJ5R20fCXwDj2pOSrYJ9lPdF68hDTXVciAU1HRlAYEbF6nVp2ZCrj+SviQLJloqnfAqFiu4Xsrn
QEyltxfLc4iKlW9g+64WcCB63HbZEf57EUdlCRb9AtFHhXlF1Nky64R9ZkxxYnja+3wK/uZFxYPs
d08SiVW2C+0s6hdFAuTHwfJEsyrLO7Rhg0gR9o7pcVSpkZ/6CiBDlA+d02JUCpD5PFOqowv7M8vJ
9tHg9Pm6tFjE4KOb/40LKQY+NfFu1OjQTUeaByS/4GeyFrIq0R9h4Jor9tjAuypBH6VNOyZ6HmbH
zjDt3H9sl6KfDdqtS5jT/sKGrUGGh14o5FiCzGlCRKoCnYbSJR3xevlWR9rQga1uuk1+ujd8MRXA
EePRiFQg3uYtMRv93LqK9XNV80VD+CMKSwzHlqOIRUiDJQvRkGsDR4DcK30q3MIrqIWDPRKsVKpq
qtjVsfxveG/gWJyg2jb/y1chWM0AoRW94ncjPCI8mRPy6aHYkNJYndWnoDWq7v/QOsZXsRQvpAdv
ycSUp/W2fiSdQcKe2oGO32SoYzH7WdAOq9OqJ3CAnUYzFwjzpJd+R0UMaAeO4l9aBS4O8P61duWg
VkKJNPfCuAnA+xqCr54jbLHQ8r4di5uUt2FZvYoTH2hej6GNi4Ik3PGcaOhbJAPUeNzn5wIuzmGi
XwRZI2xJraIqDJ2YGP6uHU9D4OX4OcHmJXrw3IppGWjwmxWg4jR5X/T2X5kyeQ7bWeTKbu6sbqyO
apcmjpyRJiV5BmZbLwHuiYGNjTTFmC016pAwjRvYfQh+WO8S/qZzTCTBrCZU/N5iJuFsdffBNC/o
cLi6OgBbuHa28zxrMKVQdPRSpFRFORIbeYr40goh5BviT9mVuxgAVmcEgCUu9Pspdba/TcQvDT5+
IlG9MUMNg1+QpIrdVNvoYLbW2rA7hCH6YfRDh/uNfvmAiqKu6IbMpeGmJVB66QaQuxAL9ZHw2i9A
RqAsPS6opVEeUQ5JCPPcx/AzxYm/PhpJ8kp8gd9D6VRqVSy72vKXEoUB9mlA/aYMDFzAIqdWCCm7
3IVqR0oZAB73Vm62Y+8ro/2J5sQqV6+jGYAccYu64nHY7pX4j+8foEZGaIUXNBNyj7O98W2Bqbu8
ePcOFLF32TvCnTdaOqjWvobaTjLu/OnssFzE6lpTgF1JC73AAMEI4jzy8HnNYg+LKZzvwR8dSXtp
Y1pFJ8iMP3TOKuPvQNLYLuiqOMr/lT1D7Mo7SbNbuN2Qgze6U+rlb4IXI1R4jSUKoDOjyF+wcaMI
qjMvSBqgEtw9ddDui4fSXJrtI2ULtoTpzdfpQ8VCzQ3wjw5rJKuDGiIYSsnzJF1pbH3Dioc+O3w8
mauMrtOzo3ikvz/PIjFmKC/Rb92CZk2AmnfaD1rfKa2okUqrAlca80k6VmGEiVMfCrI0DCsS5xhm
aYrtJwT24HZzeAwHSD4KA1wV3EHPIRHJVsGzOPNqxnVZ77fKubB0pBzXEoFFZK6ZClJ2wTehZq05
utyHG0pAkhAPsQsdyJnj5v5n3BSSJkJFpD4uNxx8SgG03aDicz3dcjXohHoiT70k7SVktYCyozWq
YpLfM1PHkPAikcLAZrm0czvkiTp6QJS6GDVPJWnNSOadLdRgwLK1xYRmjhqmZ8UXRiMtYarMRZNT
TpdYOMhBfOnOZzQA6HVA4tw/2bufiA+hBiLv1CEZ1qEwPX/L7DOh+whqo5leGF2RdVnuJcKBTJPz
y87Cz9sjTDcfi2d8SD/CV/6xgTOWhzHR1FOV2Oh/VOIq+xiTiGm0/SrsqJmLU+m/UYdEI1CLHJvm
O7MJFnBHYMaijzzyicOvRhSRIB0ZLrbSelHzPLHM8mo/+ubPObY+1eAlNt7HxeRf9c13a7KyJqKA
mQJyZLdu48SeV87unYSm/1K3sMZsFNxOGoYpPFYy0KM+e0yYtCpxjMBfHKIf2WpslEMA+bpGmJan
EXXfYaKOn8S7On1fypOOqztGHy8RUBQscskfa3P+aZRYghzpL4ZIKDcxGclXVpLv33JJQnGf/5nv
eiEioKZznu6bpsDt8TvtSZDK7vXTdlk7xf/0dfT2Oq8380OZe/08zWyRhgwfUoEVqdwcULWzOPWR
uEyzBZo2lDaW62hAYbPlBBNnidQmn8cpb/XCsOT38M+13iklHwOwaFD8SFPwqJeebo5OxP4p6OP+
92J/DTIji+zKN5m10kNNymY1Cx4qNAiknVJ6IAlZToSetqaCwOhR0vq/7D+P/G45gCytOKsI/aed
um98Hcw/MvteIjyscSd3i886skah6lsh6jNCNfeWIc3kXrvp0Cny/tqUKngol1Rw6ed1x8ZTj+bC
wRoWcBuiuYt0zgf5k4JH4jbHuocBl1OOlw31VT7vKLM+Fr3LikVAzm3DORr3AKctrgJ9UQ0eNp6+
cp44i9StNfleoJqQPFEHA07mu6935PVEfR06+7tp/kJccVl659Z/JIvv46FZ4NudLcaxr/FNG65C
EPCwKk8MbbhCBK0W7Cd0D1UwQBiMOxTWoB20+o9eXvttjDcCkN8lANdkihnn7u7ISxutfkUyw/W+
SArcT4gexWO+9n0Qpa/6L9jf++EZzBB/ip1gDUlEbo7IPjWbxRg0oWsThdFZkWAT1cjABiRGPXBM
zzyDPQ6OTlxf+JceCjkcFOFUsNtvQp+xKu1/q9Gbfp+s692n6OXJXVj+DTbdx/dYCKfEPB8N5BhV
XyOC/3p696H5mNuYJjGLrevN1K919G42CfJtNy87+84X6J0b2eSahRfOnsfb2XLDgxeFMLQ3OLJY
n9PRQO2s6Yx7pKGGmULy/BUOiHLDGoXk3SCT74mKaqXY++TVGGlxaHAD2vd/JrMC087SSsmHja6/
qAB18hCoD6dbbqnCCcBHCSaHHVlY3bb8wdBpY5DcbjgOXrjFuDW834yFwLDd/wAThDeY8Axexxt1
gVS2WxM/BHtAKobYlkOH8zTQ7Dz533AoEsP22tEVHW012k+0L1TLjEDF9KZguoPQqe1kI6WI1iLu
PN7a3zxMpaOFJRm0Qb7usMdQhNOHmWjsX17ph/40BLn0j8N38G11lDzhRFMF7radqeaN9pY6DzXn
TsPDIqUy3Mp9VCT4682U30VqAeeME9dTtHQCzn935Q6PPKo1RJQMGjfbk+mQ2sWcO6cF2JAsfrSj
elYqDP5gpnH9Oll808eTTkvjdWMADUY/a3AifbfcrJY7sPOyUUSeXZSjsG3141kBkzkab4zZAPqL
Y4tt0Gcj7NMx+Zt57Ro8Fk4vLGD/QfM4IS2Bs9o3IjskwMZZYXj2hLVe/gcSK2dy3ZRHT+Arp48G
LzFvLnCGGKqPtcvNVRjsfoIXLqorNxk339doonRze8aEVR0+AqHHyWftJMB772BcixEtdgJ6UeoK
5XNd1UYUd3KIi2yQhyOlHcjEq8TvRQ2cJ2cR48jn6AdtDzuWNgk3clXcOtBFlItR1DkVYbhHbKzl
ilsLwrRVMOjr7ui0baqu21bU0RpLj8PhHYkl8ZDoetD3BCuVFA1DQu2OyqhF27aswIkZDZ1vZtaT
c91VNT8yhU21w1kSuOYUpdBjBlcjmNMg+843AQ6F7xKY1yDdHKuyoHdB8T9MZodK8SC+Tj86cTD2
ifWhbELLP9FATU41De7IBA4sfYy1FZnJlE0GxV23L3tf5unnO29weHmVqAWR1KX/cm6vzxQP5C0z
ILmm9yIzAfYAsuy3t4HE03te64YFjIw2eCkt+8Yx6AGa219bgmFUKCqzQRs+Hl59aG8QG7zvXnDe
tSDc2w/WYeREuwTmsLi93/2M4pAym0I6DUDqtZZM7K+3aAGxQsJJwe5WmFJz/zh27JHJ18uWk6QX
GXF59//JTBdRItxkTcaQaN1oSxYnsAbAIuiu4C8QkuTTnfghF5bCzsfeOIZmhk0V7Sgo6qu6xjQk
i9aMFujaHnevXnJb6DUg+B/dKHP32ypqbknDWkvY0cEezVNV7LtBQCf6KMPqSyacqP/B1Vcmblzt
erWpueeAMkfFVl/AuEj15WOeFbytMp8C3rh9v71c+eH5aYsTDtogc8RsaEimV2aY7OFV/a9f3QVv
WPhzEloljmXzoIPve0uklRjy81hoa5d/y90voYazhxGh7ohBIR+98UbtBWtBDQm/9TUkik8Y9G1l
fgaDRM9sV5Jd796SEC70Jp822VhCTWCaULThX/r00Y4WMl+4BKa62E3oMVIpOZsPqhAVpSMFfobt
4/UMZ9BdyFw/JyztHePYuUUlWw4X9nvFz7sNX2vwfN3JvXyqVREuWQ/zwZoutDn/V19PhAryhPD2
CCFqYcw5DXCznMZjnzbRz5MtdMij7sqA9mjzcGWzkUd1wNXb7oDSgLFsKwz38/MmG1MoDjw5uslW
JrGvow4ltE6DTfSuv5apEXX9kSPvd7MfArZq45KBmw6KGp6wBhobYPw6Z4ZyKo3va2tFg1mnz3+S
nIbdt2WCJVu+t8XrtdVykyrSgIjtyNdbeZLlues8NoUYN4+QZDsU13pwmfdJcCEs5w/3pJkQdzTN
Y0BQE/5RIWOScZ5c0wUwLbYUkG15WpPljREFZI88XQk83KkywgtpKtEXotY0MBPn3/0qNHXPQNEE
jk7xgf7OOvzMGQDNs+nHB3Bv3Z2S3lQkX0utYu5X3GSvtfY5QdRr7NPWuIe0ziCNq7FWbX6DKGD5
zmLS6QMHg9dfso8iGW5D+htYPIa262svaxm7V/5qYuJ8VNMYhRmRuNIQAO5BUGARmFRyEikXopLJ
waSsycQE1dWspGbZQbwpF3yRSv6sxI2DYBfskfJDyVYSjsqQBvExHhUE88Smma/v4pfxeUep3OYa
QFvNS3NIYGt6MMXr0MA7P/aiUOKvrN89TcXC74mxo1N/xRUlxkXXKRUFCMQmhDfpE3VxW7ULB3X1
bkOumxwJgp3zPANqwo+pKEvnCIADB31SlQOWrskSrvfCKrmhsYH/C+4iR8V16DEh5WivAFtPIExk
t9O568WIV3CoqNoDEgKmxCSbDih5ayxY0UVRUPPqDzuuDKcHLADB/OC9bgwgaxonDRcLwrfeJlVZ
kiC29hALVvrgFf9bFCgQ8eCkLo85+Gcx1bsNxhoMsClYR4yHqwVKLYiftA2LbZV9bjL4qATAgWif
W5XZUE/qiRl1Er4OTEtWlYvqB7OheMWoiGK/lnjI9p6bN+E4j4cjAQ444Hud90bkCiEEHYo9du4m
3HjsgnIkLQvyXNYGX3ZPJvh/3Y9sHTAckn8Qw5fqCXVHf7RLePIpWaIRStUzyAh06FoehKubLIjA
AIyUvGFdXpAee9WIoZRNM41GCLVsLOjhOQh4vjXWEHbwybuQF6Jnb6veqBfT+hRRCSIBRwEMT3yZ
9cl4hTfmdlzV0iiC8zbbmeHCIokOlXC4fkJAfBFrRF8mA6L80xMcZFeK8JTagSoKPGjCOpw7cuKf
YtKEUE5vUXC9DzXxBS6wIpVCq01LHfk6ssjQVhe9rFjIDLHLa+E53LRbfJZxJek1Bcz1d2J+irOb
g2qaQnkqufiFZzVyLS80ZP1m5z7Tpfc9TCjYxDr5rLWB+U5MbaMvf/X2fLT9mB8q9WO5oH7utKpZ
HbKfCjgDrokWjTKXvdVh+kmv0/imXYttnoAzpGfOaoUhZ7WlH37o8EiyKF/FfzHtIpz1ZulCcyVH
6Ndw+ZqT/TDy/izVdQPy7zuam/4zF+F6MS9N+Po0iDr318P0sS4+x6PSOz/LmUct6qwm+egvqK20
jDbOlHik5KAmi2PkWT0ZhHue0PVejpAgYcSJ4n8i0ryGtHC3zFlVShSHK/dSgpbwjCfB301MFVzH
qJJzzH7YwW9a96MDcRxTNVRp/oMSGsoORKD4eZzMJwd7+Q11C40dUBupkoxOT8cH0YzHKCb3tX3I
lbkw0S+APilQig/lVDAP1hh7PXJu3Uml43krMxO77Fre4CT/yt7p5Pt6h9UGKK5c/h5wfIFba31A
PsHdSoqpn2xHrigctmhUtF/fgskuHP8l4XlJ3h02SN2VPH80T7FCJHvkbVBqPJPl6z86mM+yDC5j
9HYiILNKjiym+8yz4cRvZDJtr3Xk0X4rrEaVWtjL0qo3OOi20pLkF3MkitCcEF7UOIWgB4x1fKPV
6+sPybaWituPn7ACOY4jHYp1X0xUChBt3Ay264azX+MyMEly5B/2weqWcRcEAL5owwFNavv7SqOS
yLaLDt4T+v2l9wfoMKpG4nVgq+YHT7rFAatwKpP6yM8Cvakf53bGLTkm4R7nl2yI21tAFAjcSzji
IO3l6KMrW4TS1BNLUOfl9ufApMvbkqb8iuoUY2JdFVM79K4l/xnJlXyURsl3DFFcFpXhGr2+nLXg
JjcLO1FLuAUTzZscy2gruV5xvPfTkDbztzlNLffg1z0XvD4n1kEHcNPPIrgM3pX//lHp4d89/2W3
CAwrHTQNI1toiXV9Z16hSBbSGIhC0Mz1S+sPYyYrgSRLfl9/Duazwmmlmb1gO/y88JDmWl/jnLol
hDtSKQwH0z5iwC8HUVd4WrJ7nLG4k5pc9yKt2F0+91XDpfpUZAWBk28LSDnf3oUCPr1ExoWeELgR
BJzP8Asu7QjdLtmOwGoUKqD+eBXM/L/BZJkVMLck+AratZyWaKGYMVtYZaW805OcIWq+Wfv9LkmB
54RNLWBOJ7z2z1rV2Bmoe6i/Glu0Ovbjm/8nC7uL3hZ0Ao543dpXSSMdqR4ZSYUWYBCYvEKplxcQ
bsAF12n520l4OPTyXG3xTE8cjsG8eCYev1em5KE95V4UOkZuLieyr4U4sjfi52hlSBL5i9/e5182
ola99LTmTpzyOV/vCdZUPC6qWo1otsBGVD6rVMNw/SXOHsFIzxQW0eGZdj4iC6QHhbumebOWhjED
RZcri8D71b3NPtDg8a/VfnEW72yRm71VcPSVG4d90vreSh0s3qTs615RMArvyY5oyVY4gpqSUBw4
NmiyYubnsd3tt1ETHlF2SXvn3Y4y+/H9xqWLjiPxfcT+PCwrkmosBmBTBkwIH9mHYTour07aCGjF
ca6zfMZPIUg3Iv8PSxgR/NEb13m0j+KGNpD0y+vn9QQExyealpwzUDvouG5Uk5cKAylagxpXI8hb
WWzoB8uR6M7dg0ghvyPVdYKeQvDe1qMLgVt9n6IZxYVTgmLyj4Y9ayoGwQFfQacbxY99kW+Dc+3G
CRR7uLBE8yrQwB7n1EAI0Qnx8sMeL4QkhR6ZvKefpktgsFLQFpVG95G/tl4raE4tDM+f6y+bRlc6
j7FHHYoecSNvlAAEsDB5nW3KqOPWuPp0gKAKoD/m4hXFsjCQKY6+Dk7MIPy37u7A+37EjSi63qib
9qSgW92lJVNsrlepTEcMOZ9cxMxdkpCY60HIqRDleNrpu60eqHdYmQMJxRzKQ9amGqxWROccmnEg
xF4Gt3Men3LJOZF+6et9XRztMO6C6IDiBrD134Xnq7JfbQxGteCXaNYw7WoAlciREnTrkDB4cTyf
Hh7kcUOIQXouXvN5c+hd532DNedZZp5kpIKNP3PsWhLENmRDLlsA/r9mX8SnWjHFHaW9mnemhVia
GTkxOSoYJ/B7F+QIXHjgs+2ZjpZ9pIJ7l4jUoUdaCNQin0EbYiuFMbqgKlrXJ0RsdTvnW/NYOLaV
mQVmWNxBVbOg/YOYz9Q764lU9pZhtlSSTG/8fo02VOYkNWJq7FopW8V8IqoXT3a9kc4r4DWZOl6A
/zZ014qMTQ7N/+VhaBcwcTzm1rwI/6XPyIa+hYvxaui7/hLMRlAfDGIWXUOm0/2b/hW+qXpuTZb4
zyA+MkoimQ/vH4GKZUX3/gophi2UYM/nozFRVVkAouWYLcCOQPqUWo+W4popHSUgNXT3Okt47DDm
AOC8v60hG70cVCJfZQW/JhJ6pJtAP/LfkBld1MTHZCmibgS07MEHAAc64hO2All0Mf6NMUQW2BP6
eEWUKevU4kj0TE6XvAHdDXMVEq9z1azbCxJ9E6R9qhBdMhPZpXPdswzwarB9C4Cq/BhsF+HMwG8n
/4FjoRFndsJtu/YHkwRRAzGJZzlf/2zajUSHbi1dDyBho9ZQS9Kg0vmKcxajn3WeHp7k0Nk+Kk3S
jgIfNGH+2wBBYWLeUNbLdUnYjwXjAbW4/YYdUwhEfUqOX48OsbYbfvrl5BXuUVcHnFmAvEa5UQjC
0P9XGZYxgMd4iSwN/4IVf5svEVIQB77BNKXZN9nhM1rd30Ql8bUK+4bgl7TPHvyQkbaVVcuJ5ZXB
6e6gDiyPU7MavSLbiDpyGmGk+LaJyIEoeo37Pg5C4bjyaBNeP7h50KnanMLSHpmz9YqeYxJEwKxn
UffTN7Nqk77i6pcLoidLGkfMEqMERjmFb7sT2zRpEOU6ksgnRB5gI7GhFmMVrt3aoj+saiB3EI+c
iKyn/tNt/sZBt46QgzPUc3m11xji+MrENnTusK5uT51yQ8npOPtiEc8VqlsQXGYqZRkXyRMZayrU
TLB1MexwKJqI/s6QHxMId8W5PgXEd9lgZtdEolCbuB9+597z87gW97RwCr3HYDrMFLY9cm8m1SRN
uWbPtMGJGPCl+/IM6Wj3ijW/CvBSgql58YR2TPcnjSEljJgbXIp5e7BaUzYImQhCh9yU1DGkqMdO
gTmkMK2qBZHkn1AzL0rrAz8tFAr1pn95NkUdg07aV6NCGqrV+fGZnFTbqnMXpwv0h4NFwmKNWfbA
YhOz23dEKau0UpxIrADozpkeFO4hG1+yLrjczCiXXNg9aERr4f93eEh4PgVjRY+4NdmZRdKpIyFR
8+EnPOL9sH2uCeBMTEO39EFTiNEArTNqQVpnurJWnWQi3LzIGCGJpPNR37h9x23aOVLdGqXNtk6g
sVWxn+Ji9OlLfNoNlw1Kn1jZZ8SKYJmyvtQvXwSiSBBqEQsWOtV4M5GoU4Czt8GaqeeozAZ/yoYH
Xp125mSvVqfyNvmv8IcsWjHBhB4fXWeIFXlh6qt41ZxX2SLyZFraWpOscZsRGikfagds+Nvi0863
ytLXzLzVokh8eXLqPTNvjC/uK3ZlrWsc9tMZf9BfAlZKlTYgu9L2kamf3EXdvI7AkRgYOGpNcw4o
Pu48Vc18CVZu/FGp0ERsaTS7Yj75PPGdQQ+lpR5zHwTATf91BSZYWLZzLXej3WRXlGP9NgE4qQ10
jq4w44j8T6xtq9OiFkwDcKWtP3ztLJjjYvvH70MDEeTq02/OVBmCBprfPOA9atG6WwZQsShijoC0
HxLnwCw60UOlNrBGtrrrc202N/v4bSl7hpiT7BcZM4EXJLIeOaj1Ix1SZ8OS3vb1Zpw9AOmJ6nr9
gdFCwxm2+FkA43e5BIM/kXOo9RgL6H/LfAqiHjQ75SSTCpKNtZjKaChOBiAd/bxZzwnMD6S9mZNN
8tAWNMrqSJ9DRufvUhTZ/+5Yaeycm6evsoeLbjN9pb2snk17uH4OGwSAM5jrKL0YBeqLp1qT1cCG
xwYvT+HSalkrYxJ5wFI+ZLu5xYA2hVZ9aM/QDlJpQMwIpTNPTUn114eFtR1/hulaVJJPDF+BUUYw
qQrYMSXkWx8u95lyUXobgV1RrZjWGz4migp4XXpsdxGfMwkp7bUEr3bQ9W/Bxaf6Ssq/cJEOlu79
k0+jr7Bo5xJa4xrg2b1/WPJ4zqA7qQs4UGCw+mmxcuR/YEF3gC9YthA3bybJ6fNcoogCnNQLE78O
5dpJGVgsQiI138y+mkx72BERN+6pTdaL/t2xji7x9Zp+eNiStYRdXLjTBO5x9NwRN3ydF4V8sES5
D3OxD61GY/0ZQafPFEPUNiyjWIbf6DjzdVGD1PJlE0k7IyKwQ6PrapWw1IUwU24p7CVlAh8mk+dl
LTzPmcYaBl4piRTmRBRgXR+oLtnsPt0DSeQ9mr5kpYtot9Zc80OVblUxhJ3xqitUeu5N6Li1e7kJ
4YwsIKPQ4Kh0xzv49NTX0EQ9+G9Vhedu4kg+caFe6262qt8jA+th6N2UDmsfzdQR+M8YPP7u99WP
KAzIwLelEdHoEgFxllkHty0PttW+UaPWnom+85LonGx1oUdwgW3/kMcoLwyncEWhS5oMFEq7sVBS
Js3fkSRGgZdW2LQIADt/d43BMO39LkkikrpSPzj8ahb1G+uqMUveUW+XG84gPdyINxoro6aJMt5l
Vo8jqtWhIiXYvHB5XiLWSCInGiOxqrl00rGqhmZ3XhH0RwqjZHQzCd2fmnyk7UYVQeDDbMwGRF6X
UOuVoIZ96Ldc7rgMYTpJb+jDKTmkmjROpZhD/Xm1YQhwYp13RjLZvHcrfzxRo4JKUt1CHAwqOZ8S
yobtHBK3Gvew+tCpYWiBORZcAW2X4guY81RB1z3tirXF6JXVME5rRRssctqMWOZ+MnLqZWG5iHz0
q0HxcR9s5SO7VfSPbN0tTSfsI6BlNT1psWufkW1+QNYorTkWHXtv1qpwwDtJDiAuz9cYRBgtg/RX
tVEtd2KTcUFmQPHhPn1CR+4PNe7j+lrgTBM4BFiLDVLcZ3wHDnkxqIhO6W1n+gujvHGaVCwrgl6u
/UGMmGBLGzN3cyc7XEuDSRe+ii2GlaRLDbctSVUm6bQdFpdJkM4g/Fh3J0URTC9Xt+Ym4Wny5rp0
dcRmqnMyDv3f6r5mjyTvx8KymEZiCCO/QZF/eMv/2GbuHguKXTm9+BYY/1F5+kdQUPSf1+j2/Kgv
XsMWcS7P7MPLFKBYS5rqzqm7nj6Qjzbihkwq8nqRphWgZMv86Wl5fV9QxJx75uR/zg9yxzI7k14S
2Or2t5d7+2sqyQcS0iuo28S2QtKJ9zSYz2R7uMpsHeu+AMxLkGsADVqXmEdzrCyoMBKkb0WogCQi
OcxocgmNepdKEX4B69jDrENzKxVYWXyXX7J7hjQ7YLHHxlAgawHx0Sr07J7cUg5c5EmxM3SI+kXj
hGfD652E8QIebaWZXW129mefxw51lz9xIFc5wVmkmqvG2Pdzo6QuQbLnN73JaOhS9SursGzFI2qS
JvUEldCq+mUQg2fi2r3mCroYU5tbWN0d0OWx+UD0qJOd1oMp07gYtXsf0iGHpHB5Pe2VbR48XWZ4
UzD6rWi1nB8cR65eixzfUo+kLdMuHPPwR10imE7uJFeUsPpEnpayb7VgsmYmjru1C5fFV3twxe1f
J04H3zY3RzTg19TDxPhDzJt+MO7rT+MT4VClXQjm0hIqOwGSmOY5IkA/vATkXSaGMSG8+Sbhx7Sq
8raBVA6ShGMwERRk/Q9u/wcbBY0A9E+yeaGw47uW+MUNKPiQ+pou/UgWtLRWe4CUuuJ+Kl33uc1Z
vjijnvoDarRvv9KtgsBBtKORerGcpEezgkuaToIqlfD9jqI1b3boL4Hgnl8ztTu1slim0NfqqjTP
+f6YreyG/wXsmmxxI98NK8zGwr8Gpximbfs71GeKWbx2eg/Ma7NXrp030vEAEF9Z6lny6d8wbk1s
uSKgE0XDd/IAkNNYflRRYZjtFkQQZRVj0Mj+uQ22dOIX2T7Mm1toRgeyF7zGaHBwfN4kcn37xp1N
PRqxUYrZBOHaGgYwFtIC46H/J6+TWpWlBcezF/+WBGC64Ic/N42kB7iM29B3U8riAtJRUVq8Cg8m
mdySy/W+jLv7Olgz2SPsJlrzvq6NscQGnInkd5VSGssOGLUIKYWwJJnEe8UlUKzgf0HtmzOdbf0q
LOe1IBdDqNn7x0OwDKTlYlRBgEJ+34Mti4HMLaNOSrz22/uM2LbFa34A8BC7QVIhhWkDd/PVJlJi
4jumyDTIeZQcfJjOOEWnC0+QySZGld//PEsrZuC+xE/9tpEXAKfSzoglwLE57wwYs/ubLeaGeQhr
1VyGFR0xDByxw+XKxHrtyGfPkbvv4PPMKPktJrqJ//+fFR1VX1CK1M0YFKaz4YVycQ7HmY85Sc71
ZrgD09SW8q11/sXBvLKCQymq5EF03jeequJvVNURY7TheOF9AAIpPmaNsuNtc/nMjvANpy/i7pbl
hTDUhYfTqFPuy/RI7WOKwinWEuOXOo+Kle9NY5eMw7XxCVlmAs59+36WxI3E4wq3BJmWKhc4ojeh
YV4ohhaGf136NaDwJEXUi6imBHRwOIkmq5Fyjr3SzIhbQc11p8HxcW25Ia109KkbkevItSowfnpl
sKttTc20lLPvWYkgXlXkpRF570Yml6Rab49PoLAxuGw+kaURsmgdGyV7hO0019WXfJVc3RBgqHGK
pkqaVDgE6Wz9zqUpC0xXB8oaz4hOez/QvSG8u+Wv/+Bbhdbz9ZtpIc1bfBpyabaOX14yHqlMjD3g
IBDnY6juvgB1gGxl+S4pbwAwqWK8Ywhs4oWVLuzx0eaXPthX2o+VsDyQs+hYKSExDMlq9ZOs8dlp
4PLPTBIC/pq1yetKKmOwgQ1Ehm8i+x+XmU4I7pS10az2hSYGVhcsNJKZAL2YZN/pNiYnioF1nl10
kTrJYUlBVAKzQrXcK7AcSoX4+wEPB09GGUrVwfexiQn3y0XNiyo2Qz53cTNRd+A4Frx1c3zHXeGM
Ox29wkPJW/w3XPrco2USsGPA2wJlJlYmqhoC66AbAbfvFBbm1J0OQSmkGJzmPfwqw9QWems/NSwI
BRmA13T5XzP80W1wt5dJZoI1NSCZxAzd8JuoG0x8SJnB5ZUbC/+C1mXRymABrCRYgm8lINsx9nRN
XhtXt608AJeCF6IIxu43o8of2bj+bxKO6yJNx5A40wW57wpjhoy7HWmiwbHKV78NrkUj2iG9N6GU
BuYDXd1sadsADmhj5I1kF07N5tsPXMAraeHZI2heZ6QW/KjFgIMun8XPayyXdMvtZzzgJUr0eGtT
HModYUxVwJWKs8w3i4vq4dZJTpKLwB0LHqsgBNvHtH/h6bjNfCH0hfqgChxgJRtxpbhEgUWHCMxt
tBJ5co/H/7XqlgOS2GSGQrcvx8iI8LMxAzAOkmTshjJb43ePxd/6YCbsfW0ADpokPt1XIJnhpX7n
it3+iiP0EW1GsvkNDKHZdffk3m/qaMeh5yvTD4mU4gW4DK/wWzL5RbPqg6qxcS2TzbJJwXofAU8H
ewTC9RZ/kNjdMQjwFLfEsNvBMQTGfp5aiZdbdlXwGCEdLbrxhFpIXgpib+i1aMIIoVYi4dOtfIjv
39DC0stSRHTJRs635KLwBXvj2rRXZ7tBPitYkQaPC30JObgSikHx6KJJrhYj0FAWu4gjLtFWMg6R
IZSa7gi1jDHyJzFfNVNIQl0gn82Yrjpg2rFHrrGv8zp9ax4S7mU/lmmjEkmRovWyVZ2ee9gMdGP2
emdsw+XcmBlsECDwBGk2DS4NUEVn/dPjJ5B/yj0lEtNEzQa+DqBwGvNqefrCzavPaMRIb/Tcoa9/
IuNnOdLN5D0rCbSBEF6luklBC+KM10bXco/niCQ40FXp3OuXPI66/VCHl31R43XGp2OjWxj+y8pO
qoIowoM/63BHMfzKba4uGezKiw4VYVr+5HJ+ZBo35AGWvD1lMTHjhpMlVUwF3vzl7hRr1ebJYGmT
MivTiiL9kwPYYUHFOrob2d6Bzq8lUm/TDnqAGo9o9Ct0KZeAum5MHMMvKriZJhySF8pLPEoqIfpG
/4N5WyUgQ4iYcaqsxErw+cO4FljCn1e/8MAotSpOVxRgoj0wZoh2F0aHRQ/A2Zr/+RKV06MGQKPD
Qq+HHaynm62zfQGDRv9gkG2P2dNbXTRPrNIUC+m3UVa1eRiaRFIZGJCd6g6zoD++xIQh9qKaqr7i
kGLcjPDk1tkgkdXY0Koo0dqfLq3/U7MMQMIj/706pNvZTqcq8OiIdRiDI9x83X65bab3Wt0w8tDF
uH6Vx9g44j7z58AtFT1mwYp0WAzrMZ+Ip4L7s35qHU3mmhvdSBKnBZjcYGaSmtEUlN75T/c3uT4h
qpe0bI1UDajV5i73OcFtwB8Njcg5/P+F3fNmeHuiuhdqohfa7L7GIlZimT9DtfDgKZhXgUKF5/dL
AB3FosAtnoqZ898HtJaJx86ArG2Ho20TDn+xYN6/gSveGsRKL6RO1B3iGew5TDX7q07y117seOdP
/0RvcoRR9ROq8QhNGvEdNDbx3NOMXoH8Vp0q607GuEV0BgxVBwQU3slrQAK+0qHF3Fmg1ccREviD
TqI8X7H6IjlW6ptok7T8CRJtmDeu3d7cDWYoRzFSW1wd1UJoL45dVUveUc/te5OmC2vRMo2kMQKe
RVtPrnH0dJWULCSUD6Rd2eQbRrzLYUK7Be6T5KwACdGQYMC5Ek2jHyZrobevY46Ts7W3uWtyE9wR
UblBaXngTnmSbYg97mm/Gy1V8MJ6xf7uoJkQwVhVMHLPSL3wVWcdDEDCcMaE91mz+w4MbvtG2lnA
wvIOY/mQRr8/a/teHqsLE95nQf1QW5HJCSdzpvnOWH64/nveQoRo34JajjoYb23g6cH0NVDRbVhz
Xx0E7A+VAk4YMk9x5944AY6ZylcHur9+OeiAP/wyLz5O03X2BvpxsDTPc6U7QygLRmgK2B1rq2SX
At5wk9icqZX8vWzZo4iyVVs9Rkd664Pom5JCwfJjcFORfxssqIXQ5NI1Z6ntK5MVoquTD5saYvJ1
DAG7Dof7coZ978j6fQsAJWPoLrbOMRGGsTDD5a9z+xeGLYdU9uaO5A1xnnBZehIJcSru0VkUDZ5P
hghwLNj/5TMfZdbF3NNYQp/BG1p12v3sDWG08zlAFTAXgi1JjQMpbyMdAHvSe+GHskJmPWDDCwYy
F/v3mE/Dpi7R3z/eBzGBWiB/VRseQARIuCMCtK1GnJWEai5QAlNcBef6VywVGNIxCI6b1URlMxjE
tXgE+stRHHxhu9TzfgxdHDxdMUZsHlJKYoYzQl9zEKpRWcXf5innnMyw4Fp9yrxTTGTNu6Dlqh5r
T+SKlA9HSx9Gd9xsMnLYCaBi6/uJ/iRdok4/ksYMyA3vKAGhxNawbIHyltcr4DnhraJZGdkGY3IK
Wj1nzxbuXLLZBvrx4jUJRpvXVx5uc2XdfU/W6CTh0H6j5tHyqIOGsmHCORFs0l3BZ+1yODioQ0pl
mefbtdOjgQib8WivNmCjg7zgwctysaTN7Yc9UzPSz2Z7UilnG9Tcf8ajWVxc1A8fsRctdlrKUQlz
SvollMkRsvmFoixPN/AH9zdGtVxgHKXYhsufmafzmw149OGvSAFSKB01DBRes5LGJBUOJJejK14C
CoF8RDc0K/GrdK6vkY1rH0zyHyTnPBAOaXTk05IEm30P4Msr9ZH+X1FOlvp6FYPme7E3IH1NIbVh
TFB0RMmTwqwbKWKZLLcmcZdDSB8huTowfyQAo6VD5RxJzU4futzhZdH9aq2sbQVLXHw8S59rraBa
d9mpEk1ZMini6JH9wGZxSXFMF8Bq6uLg0wTkK2CttAmJbPn5At7sWh/NYZ3XoGVovoQG8m9Ivu5H
EL5+KhhuANjxi4xwYaUmkwb/Upxe2/lb7GkvDOTJ/tVRyRgA+ILdzwV3Fvl917VxeSUzHTdHx6HC
4S6ejqSI6fTVkMg9IYiko8/2XByyaQeU3hQfmGfR+erFSXgqEcjVksqvX8l6gxwN+ZDzgOCSEmAF
D5LXoWUW6dfiOY30mF6l6mshUMRweH8SpnHK1py/yk7s8G0Z0G0pqMeIPSFIHuur6uM3vY/g3uZU
53JwpADzvry0LN0noybZc1e6UCVJm2xAkapn/rJaWKz18c5lrRCTVJWkMeWr6luIFZp/EGAKCnmi
YyN5DXFeEoPmf/Lp30xKWKwXJfWZJ+WaT8LzMyHT6BUm5BgJS626DghiGwyoCMuKQzfyxPzLHRML
ORr2I8Fws+9u9BQdn5SbZ5lLXnNSXD/umQhNumfU38nJf1Z1MMFtxGXQbF+z9OwRRXLerlTZKdF6
jxfPJjXJpi9dUzNb9h3BIbYBSC4/DghHWD0ZTeN4NBvO/+xWj1ThmtHzKlpJGJrpQXDFOFZ+wmoA
MGFPyGiJ6wVk6zQwtQPyhlcVTQRFLFL6w+wKx2lX3yS+OnAmUIdpyvN8bMs5Vn4KuZHZFXj8FXSI
im0iGTOXbHW4tAAP3JCDy1n5DjnPcbLAqaH+Qt2k5F+xY9cMSZ+9uTN+k/BfUiREQkuR5G+j7Oll
y3nctGCXvN1N/fMxTDyroGy9NxIU8fSq5//86DdQ2GBGaf5FIBT/UoP/y2ofMzFy6xXZQw++kicS
8deMk+6ZYBAwX7FxCXreKZEGCqqQZctY0EsVQMRz1Mlc1LVFuva70NRYMGzMl6LeZCt+tCyol0bH
xGOqKmRSslpIYGOIiIuwV4obchw5030xOCiIy0Bwb605RyyRLlIAVCWvHvS42Ju0fIh3h4K8oSA9
bcMy3BsYNG99eFvE0KBzs8tSOE6QATm71DM8tk2NsvairGBJwwLgH3nicEdiJRuGz6nHVS3zw5se
xZPwR5cYsqMd56BTAhhQ9svEAepI9+JjDxGIh3Ar+horE3u00FLJupaD4CvB4ig4Hr9wFSk5IflK
kZ4y0/Q5tUr8RdGIrMmNn14xOCfyn9pC3VyfeyE+F4qN3sXGIR25pO1yL+Z5YcOIrW+LaSDslQVV
KjpW+avPBlqEzXfJAo3/7upUP/XlV2fJj4CveucOoUBqfHyLI5rcQVXQVUX3I6kGu6Ed8BBjhO/T
odBV83h1QFXBs3mH0e5XJrlFtT0OHYcsW4LLaHsUsYu8TAvr+vepmqrueml5xiFM4eBQge5Sf+/F
V9KsMrM2+L+RiZo8kzBJE8TCjQYHQ3BXf4GMBKAkYZoZNqWkzRSnejASojLOPzE+lP1DMpPrQ/43
XP79pryJq8RqCrS2aD361psj0hy0vPWEboL/Iz5pfVJWagWHE7c8H5fFr1w+Z/aVbIyzW9DSxhpx
XMtYulJ0SdFHceMwM4iaBxb6xvmdjf71syNrMdZi6v/fkTwGUEYBctFh/eBZVAn0JmfgsloTxfBy
cBQwmNJa9YmedxTAsd1kRZyS7ZB6Q2WNv4oPGuxCI7vRS3Ty2jj+xHccrv/nzCGNGDxUyyHd0jcm
4iv4x+nK/NoDBC9KMWsaK0d3bBpMwcK4XPj/yoKz6dXGsL1OLsLYE/tDakZ7rhmCD81UgddzNCuP
JLRm7+kKq3jMamk3egQ8NtO/oIRgF9aNhq7HbAeENPnDhOPPqaKQpro4a5guHOiJ+Sgxn2QUS1Ee
S1h1dUJ7lx9QXigUTjMoo18nPteUIeu+uNik4uH+fiJTU9WoLDpEIuZWvbC0tCq1ZliCpsaIwCmS
cS9wlOJMkh1gv0mZPGR5ST6V3sbhp21MBEN3e3y5pCFh7cNWinPBdUbnReNfTb8NZvkaIxySGP73
WDD+5cRtvksd0xXGxFlOALJEbvfT4OyliaAk5uypLILpgSq3USq1k7kORBVEwq8xXQcuu2LiSTS7
6kDaoAUsmebuf3WGMXD9hUKTrIz9ZazD5BC3ueDrux00/4bN46eh1QRFPn1KqOb6vwChbtNrTagD
AOhO5TC0WI5aXXui4dgQR0NmXB+C7Yibvh/y607+Zgjk9KwmafDzAQpqLnyxz0zbaF2vgT5jrkOp
+lSO9oeWB7/5ab4ny8+zt6Cr/xPqyjxyjst95c5aDW+hxYgCZxe64oZbtBMYwMnLM1RQwYZmTnog
outErK9A4Q3VdISAp6UutyABH7mQXKJQEQnWMLa452opTwFCWTWpvZlZkB4cs1kpZrLvR2cYBXOx
g2SlnTIQSdFgX29Y/DGrWVvxkrVpeEGGmG/GWGq9f1CRdtNR+NehmjHIGm5r5ZrsjRbg2+HLWaBV
JGWFgODBvQ+0SWHW2MQQc7LzKlMct6lfJQ/CkjMM2OsnU9/2E+839NB5gu6zkrwezS2zSCFw2+DA
aVfC4Z4zgUlCzdX3CciUgofidOgZlFffkaDuVQs1cpB3Rb0uDa5HYnLbI9rp/XpLqpC/5UzxG3y+
PnpjVtR6u9qfbTxkwOucUbePUWSpHlhZ0mwfzEpHzKNhoFipvVieKiLPsyiv+/sa4sFKjAhAfwIW
SqX0krr0jYfPdgTEMvUSMJJ03dr3zg3AXiFXloq5GzIx4pb33fzh0xfpzvGU9xiisw+ASoC6SzqI
fnjjmEOF22ZAmFb9cE4P0HQKIZrSAvWw118xbyCdn7QBT400ZFVZvGcvJWNwMUigKeHC+znodbV/
sfHml/Zlvos55YI3aoiN9YbQdXb1bGCBtbZJs9BNG2PhafVJtUSzceg3Oe+pKP3zDXi/mbm/Iuwr
E7xjxjQrTwgDu1JkMTTngtb/N2k1XtiU+ZKxg5+R7sBgR+VrL5MoNlYFV24qcto+P0M1FNbvwQUE
xaM4lg15t2JUh9MO/QbIx70IfzLWnFjhQX4+ff7MEN4zKmwsvg3YhXvXydULgpwYNMKwX1OwpY+P
bFsJTO2BrqXkFl1O/9JX9CdcvPq3/UUYyBXYa8hVz+uja9aekAAZjjDwiTq8ajmR0NAWYGZBAJgu
GfeY0B+gVcO8E2yePaPzSq/VRI0C07AoTprgfkoAXjdShngPTRltlN8StW40IPEx1xZFVJGzHdLm
ahDr40++C6VkXONSsf+zHqH6pcWjNWpHpx6FcCsootBI55QNOSgj1OQtDsFrf4+v3dFblXgaDPic
X0GdCOGQOQRVIRzoVtF3v8cImGpIKAG0qyD6bDRNlwpoEuTwVIfSb9qBY/vtw1S7Wic+rvMWras3
dl6ckagp+FoyTnoEqgYj0aK4c7H0B3/Y9HMtmljWp4Sh+Usg4E82TTHmW/tOKU1sK8Bl9KNJKErC
GS6W9xnL7n29Ywohg6SEvVfqAUxVHzhDs387t9E+xO/dOf+GHWH4eJKyv4dhBO4TTUnqhZnu8ma9
Ce4V5S0z8vWs95qyWfxxxEtSrmFxXDzZD1F8bpcY45ZXhHjZTV7VyJ2nu3L/H1c8DGtQI9qFVmT2
Wau/KYdvsPsevMrFmZgQdTP3F9UVrLphXCLvefegwGWdLNN6+JmhydKvnIBa0FreGDzCRrMc3N3L
Q5zHGtu+ZgPwgyyK7pPsKLPNlvw1/M1kX6bGZcy/HEkcJALEcZCh6J7+V1Aby/tXPb55nq+6JOZ2
z7vsV0yCCsKwAvE690JDatiLWgGNHGd8OVjU/0G56AO32PhWlP08KlthC1ARlL10tnilpri2Jcd9
kgtEr/oIHI8DCiSqDJt0kzQqyqzb9irkMPt1HvVKACsxG3SslYcKlGrtEf7jZArF3HK/N7ltn2BA
ZaS4sV0ScoLeCIMweFd+w+ZcufrJ9BUy0JHGJd3j9ITe4rWE+HAzfALKXEvhxlUyQS41+yQhVsxL
5Arp6tkeM1Su/gtldAMumkY0DaqZjl6g56ht0+3t4EB+ASNmE6+cT8sAFDFGET0FQZjbqlJaXN65
ZdhC+jKfTS54wH4q0fgxePm9W8ES9SW9l4h/bZmeiOgcEPEirsmvZ+F0KE//Q9UsPrHaOJUPmPGP
0Q2vXuXCVi3UmT/j14WARdnTo5pw2yaYjqmXUfZlIFH1c7Jbhkxlcj60YdqysD+5agI3MLzFumEa
x8EVzYOzWa/DrDKY4ihk6n4XkpPy7fdOBKzcsmh+IFjvhb6e3MzUpO0NwdVYhHVaCUPzJxUfsr6r
DDEuYYGYl8mroUzuwz8g9me+sivyjDWS4I4+5sBKwJEkmUJ2O1DQvu8HxHxBMYfILeThD0GyMc+f
jOtXGjdSEJK7sO5jTIm7A112VXqIH5kkVEDAOxRlNM8II5LQ/VXfCjTr+Jzm90+vLxZKpXWE3H2t
WMfiO3dNdQUD/9lctK7o7iyzJ+X4LDYfd0d3a3/FuQV1FuquTfKBMoIL+gK3ESP3p9H7X41g8EEq
CV3QCHzVc/fQTGftfAi4XyM3Q+01WQKbAElI5OzhjnfPa2h9jE8MPe0rVg+DgwSzaI1rVg1zVwZY
LiCI7qoAlpf2MtnQnCffUFwqX284pJLvuEm4blyB0c44PnxsPV+yDJFJFIitCOJvejJxzltCfTD3
hMq8dnbnIzgO2tm03XblCvCiUhnrOvI1cfrOGcRuiiJcJDNdIdDo8c19S2/8fyK+PwMtCdRoGHe4
5aBKmHRizslpTdNUsd6/DzDancS6S/KXSowY6X2gUQ8icx6gLp9I1MPNGZgi3Kvcuhi7t1Hj5Pbu
hLxOFDFP3UZau0RkIm+2gNHM2T6WSaM+cuy+dS4egPUlzNSxuu5x47kq4ewYintf+oXGpq9B2LNQ
Ukc25mcnJqcLq0IheT6g1FQVaXYAGMxjBIsQiHGWxgcV8A8SaEgW/va/ERug0RtPu/OvjeJYb8nX
TT0+PxNhLp/oH6cKVCFjZSG2LkKurr4lfy1wBeme4D4gPpmMbQ+QU03Tmj27V4wv6CtUMhTsOoTT
7fwEl4Os6blfcoflvVlWPohMan+jVu0RmEKNiNBOYi0+qUA34COu2XFpn/EkTmC669/g5wpXGP/u
zOp4PXJFydJkKlH+sNQUfNhPvvoqiTqjG8iCh85/w6uxpXgfTiCTRsht/sh6atCjqZ2k1anRYP7a
BoEcEMttAL3A+eX47/nDbzHK8MUTiFMVnI/cls3yufXIo9fzMJO6aBO/gv5OiQTciHMusCyxsIb6
wXhPrpyBG/Sc5tUdRS7pGTWkLT6WpYfvkmdZQRTji+fEOI8aczYgE2jcZ9F17CxcTuli/spq6nIq
TsdXAW8/frWCeLCz0A3JUrxQurMfBCqxTIYCmtvVcWOot2Njm04SooC7MU4EctrWA98WTVCjTkyd
kiBIywGx4nmolyTQ7KoIhlmVAhlS9NzeXG3/Yk1nep8JgVYAY7WG2WfBbfy1NjBKw34V6VKxtbKt
OfpYIBNkE4PO6L/eaaHwp0/V6225sUnFeA+pUEtKGKELyNbekGE2dy3vF5DBgUcQCAIrpQcgo4du
wk0dwp5kq2eASbHEZ/XyzKb31K2Kw+JWEsQhP/7WuFN8UhQpfsAVlc7vXbT7FbFymcd022CjSsEr
lApSyRSc0TXAeyH2h1H37Ue4Y27zfOyNlVgtUh9Fyw9jktUMTWPmxpbgXCfgH7JvzqEG/rUjz4Q1
PGISMwb1LLDt/pDIj3WUVbaJ53vIVO3B8akkGATC14lkp4elViUgdfuwsJhiqrcL9U0Xe72xDCYU
I+SgiVJQIC0A+vWHTWhTcKDUY29bEE1pSeUk7hkzuVv+11kGC2PX5KRBKM9OISCnZsx+pdC6kW3u
0hDMg2Cw4e0vtl5wPDGIp9n0ifAOdAVjPGlBImWZvVqSCFGsbk/X6Y6ZENZ6OJWYT0uHaCzyMI/S
WgdRKvnSjeEXWXmuyzNXblqewkBxqPkiz3jDy7f0uyzYT9sMV0drNhPXuS+uA5OGjP37+ncmE6cB
rRSmdkLoq08V8ywX0yJmLlhfT4SxaZbbnle82tpasOKD0MMQpDai0Lyg29D5X2Qd2n9K+/i7Eaid
e2C9uSdFR8vxOfs5OvIKdcm/o2PWiJosBMAdKqtKDdxytjxp7MkptvWY0W6iYD9bWpGr4FCzMciR
q3by2sQK1VDe7rQalglvv46dC+ktat+Nd3djNW3xj4YDPSgIdBlqlm86o6/QWtM9wbPdFAchOqWj
/HNHPBtlhadjksu0JCu7yfry0fdpsEmpGARnO4JVw0oDDkjJN/pFk72HId32ysh7YLO6BZZ3Rpig
CugCxC+QnrTwvvsXTL4ZA3fGaIy88EhtYe3ANKmqPnwX2smhUFltZg6Cgm4beoxH/vNRLStEeTL8
+juSadOTgOwPZx810AEHpqnYocKg0OaxQIVxatCy/cPlmZe9JMXJxRoMENr3FM5WLMZAWY/k5wu8
oE+4XdGHP/QTjR8G5UHPPZsmF7hdlUHX1YlNBuEdW8vP4IbZtnfHIg2XUW/2J/ydLpm9SdTTLkZH
ODxNMcyyeq5GTQ67+S8HWfcHNroN7Us0IkDriNnLtX+JsBiAa750DPG6gmzKLeN+JWGMQ72pFPxL
7w53SHWARFVtutfeoEAZN8F4sUdXckKnMMW7li2QrwSmSgt3uE7Apl1sGNSdyld6BXsVU+flgC+X
NrvbNYkoN6cJiM0QwMy3n5PdWhKfUYUcpO+tfzqlChWk8rwg4xzdpctqcOl2NiFMH/vSeIPuH81D
V8AOvgH36bwKXU0QiKQJYq6czaptfmWxBPGaf0VbvaJfUUhMrIaT7TV1EziiEsyXqfaa6Ls7H/MU
GNaD5+/JPBM/WSmGRH0iZsdomdmoblsseyvcElbvg5ahLvEcnz3hiEboW2CiR8FtcplfWOKZxIvy
x79iqXuIXWQK09vwYTLyn8SkkrMqzY7CZmGjd+bm9kXr2toJvg70rY4S9QCLY3+xFmFG7VukaB1k
xGU+9bL76xCMUfz9Z10+J2+ApFeytoNMMLFMJBJHM0qLyOwY4viRocN6hPC3uVIdftUu+/q2HjcA
a+F7ApsNAjhwpAicpY2fVmt6xbeknrsZ7C+MtJ3uLsxgYhaIgPY9aes8U6a/QhG4uRen0e+TXNc1
+p+lI5V3QRek2vTgrb5rstKAEoyZ7vJ8tgwQvPIX6igWDUIlUahP/bEjV8ORCQzdOSxOJdvRv3ng
zZhz4RE81FUwgwNAY5V8g7eEeBLXH7HWWw8N6lJTZhdONxS4bReTqLdYUXWv556q1PNLHX/7oXh6
3Ly9vlxjdhHGXF9SFJdH6uXfh/0FlEfg6/D2pYI+Vm5oZn6fnHViEg1JDv0SVN0aVBPIUZAd8xxo
KMF250jCfl/Ze1ejbCwpJqTCeEYbwUEpn4jc8rTMABs3T9kOL541DSK4/PvMfKRGAV8lM/ZR9Quw
jJn83RNAGOX8mM1Ol23IIYaa3UjtiVksfweVRd01XzSl2RQgLBl4voO0rmdhuVroPPiyhyZvLFdc
KkDScvI5c6My2hxS2FJ95C5aQXTkcZaq1WEMfh4ckHksWcGeOReT96Cwoq/fAqx6XpTxfZON/92X
7v70ZBbhArZ5VbobB7wVrpMhPIEa03a++W2XYRnD2YohmXsJfApQvnhw0f2CtEXr7B7SkwM1IOvr
2+6Dye+mXP9gGdZyMa2uHCVFF1AZo5U/VSLfDRRsU//M3SDme7kVVp0dJBB4AmLT4h3RgJTYEMAw
i5hJs0jUA2DARfYws0kaq1VBGVP53W1MoWBpyf8tpdpmJceCPYDkIOSes2RpKStCFTZ5oijWpZUt
goPIPuROByV3ixhh+EhAJzq+jEJnd1xO97Q5HuuE96p/8pd69buBLTU9Ewci9xRIMeD7Qq0s7m6p
6tXadKHFUrJVfZucaZBzywL83aJDpsFvhgIhCpQgUAGZ9PqgJrR/J7Vx+7x/EKPVTnaVU3UpMC4Z
iZ5gRW11onv/Z+UghXyvy5IRQffKi4YICZy0G7WXdUCwwWnhMqqkqPOpz83H+olhLQe73RDEhLKR
GLHhypg+KeK7ude/MV8KeJeJ7F2rIDRZ/twaGUhQf4NeBoQWOx0RH1WeBvGACDXLg9Ciuqx4BO8j
Y5g8j+k66SQxjxe4cwWwd9iqDzBH2UR55AeLth+jBMKtfLPhiOaIwRfTL8xAxZmQA3ux0oYNspyK
9H+TmeKlsrl0kiW8t853oVs691d52wM0VUFL/JB3q6pdk7Gf15qrF4rU88vu1IHN2VbBKu4W+cQg
WzWXRmr2mAPZhHvD/os8bMLybh2RnKawZViMw2HAJGHkGeX6e6d/pFj9wsu1tc+XW3SxpLqNCME9
th6iDDzyTiX0OPhfZShLmbAjIeaEw5ZmApv/qrya+/17+hGsdwDyWCe4qd3NsuLm0eqvQfCM6Aus
CoBTM3XC6zd4CM3H9VpQg0vZw1liZRiEYeJrPr0kZl+JYKFL31fFezbh/IN09zFbZ2vK9ABOLI7t
Xhih2vDbZoXo2ftyNLzmQZNYIqbA093Uz9Vvsy8xmyD4PxsS+GAW5oK5JwyfuQqRbj4SsGVBug+I
pJCzqPchRsmW0P7/VT51Pv9EisNwHuy9x7YHTeOQ8SAAmpg6/ALdmrjUBSRvI8/ez9e1n/fbnjBB
9LAYUYEplQz4z5Cv7N5FbsSDGG+/NabVIzC1hvevV8dqgmTtFKZfCxUzrNI3WowDAEB6KhOfAOUK
eKbmtYEq3PUdbXCNunCaTXliG7tN7k7Ujy/pMm0pZYhRbvPG85NFfWZ9nShf6PApTY4tDeal5TEZ
0q7ICtKyt3r0rHrFGgWfbiFRQTSVW14AUYw4x3ZPBRHjZNaNZWiwNKdimW8OJAdLC2JkJptwfruh
qk7mhUOsQy/zgmYSf4zXG/mDh7pFrHK4rWouT1zvID9gGemb1aCC2Yq5KM6DFq90jHeF3os+IxKq
cr+mqEAW6kZtPwUo/gP9/e1ps/JdmCTYAURYMv8+PkKQYcltSYfWE05wltcqkl1oJ+CepNuddLYU
RttEf50yZvi6jcRcl1fipKDV90ss/SXGzkcwU95BQ1S71LSaLSIqspGDe2tNA1dKnBK+C7m1Vrcr
7b6U98lFEiS59OeZhglOEvQHNuqVVAeUFjiR8vwa4rCwkQzOeUgK6NgUxrPEY1VOrUzZH35cJKCH
+0TZddVzKYfx0Ux8Xaen+ip7HKbGuuPNLA/UFcYX6H8cISiwjURn9NOCY2BZBDRh1DrRVbvUwhc8
E/mc+kIWuU/S1tjYnfoqztL2l41CUDzpolOFDuSr70ZW2IT1aGC0CQX3z+1eE9fDsbkaXVmXAIF3
ex8+JrnynLCExhdvItzXuqlBbnqZMhcsvfm2cSsP/UD1D31oET+qwmK9itJtF/l2L1W6gsCzXQmb
WUmJOd4p0mt015LAX8ki5PfQXnMsBNwJe/F2ngkX46eNkqUwZy5Oi6DGTPz7FJ6zsGGcsm7DjNJl
HSHd583HCm5U1ywlcvRDBI9acoxJcRKim9WZ/m5Fsh7lR+VrpSl2SvekQ0G3u7/gkA3n1A0N2SfR
owPYLfkybLLM8DQSZVsrJzedVUZFo+u8pjOC59c4xqrV80RN1kbxcIOuEnpVqo9S5Wtpq+uZbvD1
0REdwH663UT3LISHB39wrqG6Nk7bGfW0seyQBaUPVFOjKb2+S82ST7fPFEJvVGT+FYv0b4PK3cae
pLrj7roasP5kUz7Lv6kXJAQtvtR1+YZy1apBDNDAKWiyKEyYKh11hBY+UZYeA9570pHBqS4dZdTB
oFMugCg69/XykcdDbtOKMdY9mWVbFMAxLE0iWv4EkQKtWygG6bGJZh3V9lTdfQkM2VULobRdb5lw
xI4dC7588RdS6oLCCjd/VVylMzLbSuf2b6LhMNK2xfNeCM9YrXwmecEUvTKjzZU3kNqW8pUnRGkO
/sjpDyuwFWeGZfI4KuiQLURkstGhEfaK6RAG+v0t5RePXspVGkKbz/2ppmEa09TKgnowsVtH3Qt7
lSl/0F6RZzopGN3gzFsxyQj+8sZXhuD1oOoFT0xQ/2mbjOaDWVylC1qjyzdO3gg95vYt6mwN/5iA
5bo+QZGECvb81wiRj9dinFDnO3oPvsqxeunlTiOGyYSLl5Pr7oJx9v1f+friy5Akpdv18WqAQB03
oeAhASzMIDUE7r9Gqbv4CAvY09u0tj5BgT3X2Phf8n3tBjh2DkqVLHOOdIst0srVIBY184i1RDKf
qc9fjbmKykFLQHG7HrdoMFqCTX+QsNoA2iuAvZPyLlcMaDFmNz+711x5nrz7W7v8j1CnbXs2xGgQ
O11I7fktr07PPp+yXDvDbjgftpj7TCW+uJPtLmauauYQHQnugrPemP3+uAgEfNkyy1I04Q4Az1qc
xXNusO0oVXR15nOYZKlEnk4mqP4wd3TQwj/CHoxggYju+cdy5N3IOQcaiiQ0vTB9Qjgur0lLBWEG
lH621IoGOfZfW+XqPINIdtfk1fjqs2NtBTXLHIF3HbAB8A01FHfcPSXkA1VBfJ4BVlqqK+xAZour
W/sRLeLsOumgC47olONm/wDt6Xt3YfTTPIrI5ylbvcqu0v7dlh1BaLnDpML9q+p96/RsGSGiKabQ
Pem7i0VyaB074hpPVMg0MTlwGlnaLU5fOg1JFzyZgK5gQyEZtZXWTd80Ys9nBxCZK9jGfdYSpAg7
j84zjx4RrV6nRW/Bzm8pLYhs+YBpbfWHlaFCf4xaxczV1fboaJybjAOFCPWUY1Anb2DhSQm7dkez
WxpcfaD42qC3SZSd5iuh1+A9upMZD2sYbQ5JFRRjWvP2YeschpL2ztHbM4fZFSMerlcqJ9Ia1tWk
aoTKzrZQQuZhJ9m9o58PLLU0QaIehQMxzSsDXcdboUqrVrHEu6v5MqgCvWClEgmQDtoi/dH84/15
SVCUnU6D9islILdnNBIEw2tNzs2ojoJBh6H2uSqxiJiVeaujS5nHNv9FmtXv1U1X+4w12xLqqMXT
ZxSnOFk53MBZWzCWwj7y9djPb3ISSEzK1COfqMIn5KLRP7URsTIIUW56U9Fb6DUhUnCGipTAebHb
WczK5Si2TTKxV9bMss81oteThKhEimxXsi6EE2MkNnuHhDNKfs6NAAwf77xauyMbB6cBSTrFeYTI
pao/3NtNmQmqy6OCJ9fgTJLwix43zeAUB5wzj/acRspahkRHSl+GjhiYJNl8wCyQwQ+r6lXtWQMs
8n0FKfp/eI3C2B+i0SX+6EmkQlvufJxk1xDOrAX+J/+9sHIqHUZCoF1eTfOpZt8pRwu0hAZrMJyf
8uRgkmhy236Ryv1ySE2YhXU9a61Qew+1OuCyT9xNArKm8ioKQ8qH8Ty8MMj/XdR3D8sb7vvCAD2x
WPoNOmXJy8936gkbsOt/BZj1Loo7L23fjW0qwU0RNir9Fhg7A6XgTUIte9Ipy4akeQcdwWOyXFlB
WF20pzRPxOquq24kzaoCm+J4C2YdYj/QLKF10MnE8L67KlQOqlKaMFEPawC4tAYsRplg95VdQdIM
ARdCG9yhdJi7wOI9zF3fcP2IY9BOU54yD/WH+autyxAPuwOMnbHQipIXa6o4MfTPywuRNTCj2jTH
1qkzHKPX9TWzBloIx3CSSj91CgNWYZsWNJq1nWPYW73pk63sCbkqeAsJei0A1C6Se4vGWpj2z17E
zh72GxcXd8Sl2bDOobnNNWqqCVwQbpkxObp41i86fvIV2/LUQ5Vr5xhOgHN1Vc58i/0qx2hj2Yf5
TWfluAtCUxd7HcQ+M+Khf6UJGYSariTOH5kAeC8Aolida37NR5tReoVWluBJKojcTGc0ilSabOAj
BGa57SfuRmqDpeDqqRX+KMgNC27hyoSYt3CN4PuoQjWb09roe8t2LzLL8983YXYhlRvZwVfU7Yx3
VYuzes8GX/GzGlq0+9ESP4SckK7qxxUV/YrO6ugwE5SGvueODquNqBT7chJesKwC4ER7ijYnoQTZ
9VevZ296KH2O5Ke4i4zrY0PiVI5yhG5PTYtpThjnvtNmwRVXbzhsaMYzYwoLzy1zUOlKfvkqUsyA
RPx/RknHhOs4Wi+54aTMZrbai/3NI61RgIL6Enfbe50g85lYA+mmkHMoInHzY1mZJO9LzTGjqvOv
AQU+2gqKqydNglDyIOXEoFiVbVxaHg5P8aq0neCl+WD7N/wfVzVD1QY7kjiG5IlbNbInVdlEnDYy
wX8I0O9I9V3u7c7r2+njGUdBhTt8PFMx5QlgHZaIq+08YsmKEYqepwy5RVuO8aPTZSpfBCZ6zZOy
w+4E+UJ42NMBDhnDOZKx4/q/HjFmGqol9ZRivWDlyP3tVT2Xx5OxoqGalCxoQxabUNt8RP3wYIyq
x5Dyi69XPmcQRuIAROMcuAoATAAr8uMj+HpuIKAd9WqvvT+M9u9WaEG/yEwz8r4sMrhVsbJo6oMc
/nACmimNGcVFuq68ITYeJJ9SFE0DbUVRl5P3cJvgdmDfpGbMxaTKypRbp588G/zbrUo2d3TQuHSr
xrRY79cmO/PwdiH4S4JImnacaK/rn2vZDsDh4eNgdbzkMEmH9Sv3y87ff81OMDUB4sNPWxGKZnpH
v8rqwF1qpLDqpmrDtd+ShJW67IZXQ1Xl7864OwdhzOzJyhPL8lNwV8GhifNF/NSbFryDMVt8nOVp
tiXYRIaMh42BWKnJBv7grn+0SPt4WXVkhSO/0OalnVIR8dF/kGjTH137Tk2sAwHpCPasoRG4ZQ2W
7M2NK4HjqNbn5Jjbrs6g9mG9ha4ibg9hrL5S8bOm4muF3arLeAKFxtIoms4VCr1j6NW9ftPhJvYS
QGzaIozdAR9iUGQ6ejumpvZIR9ms/mdo0QBAWbq6C/lH7Gm+yA4u6owntJX4U2Oreir7Wp2n7M8C
NG4ZJ+TKPkM1IDqbEggQ748ijgUL9CR0p0mt5Geglrk5GfTFyCJzAv0529WWCUeY68NNGghk0d+4
Ru6czXsMoe3POFNtseWqvd9Zhe/GeVWfOacDPObEtLlD5d9NghxqIA+HL4icNarbWSUMQK2qGhRm
tLNW8YG6xeVyPWPW5IyvL4EeanD66RYRCV3/tQzsMKIieaVSA1tzEp0sG++GRQpQ5WuTKdvIs2Rr
Os47z+7GZLPHadvFL8t5mu0MwbahPI5GOlVw6+Y+a3Wj7wmOH43fs2wzsW4EHWclOKmdfiE/PUoI
yFxMnrzfrBFboeiTtkweXNK4mTqGcoTHFAPT6JDaE53wMjJLs5EB0NZubkXmp/Jz8+0C984bdwfE
3RlvvGcgJ6CMksyzUFCouVWmbt0wpKtzcjicN8NdMU6MKg7sf0UZ17Jk6TnCanPQyzOJtApO6Dz7
u4uSuWNyaeMErJsb0FqLaYJhK9bbx/lJDiXT763DH/ogUTj1wk8gLgHe6lSbxAESZX3jvelL8GNK
/IC7fWf5ikne0uwGhABgPPMHmN5N+jO8y40bJ2hcL+4/VSgOTO1vHGQ3xdtbooHgE23r27zL8XYr
Vgv9+y2t24VBogvpu8t+GpWcoVb/AUmlNg02FmafpWIGUwb42hPJ6+09I8zONqke+SyUOebDCdnb
ZVDh+vHQkLsaWI11zqEazb04vgCLsslkFqyUbeGNhFGj9QJeF5p7t9VVal0aWvwlzSQQWvXcb6TD
5CDBYQom2pLhCAHn03+infPlR5D5VK1nGCTw+F8D1wPzsgoEyxo7K9rv01NqhlGhOCWs2vdqBHFx
+Y1jls9XohUvHUwL8+t8n8GwW69CvnEiNNUYVyumGRS4/rpcFz8fkgNMjHNPpsfvrBxuhTz8FNde
tMplPRJ2ZoIsQiCvH7sV0iEtBnMsJ8rEWJVRfkDoPNL2j1AA+ywoFoPMLYWSRjCQRU7O0uALKjdA
a3XSyh6Y92CVD3XKxyarrj+LQtdUGY1NX1YTYAkcWCVY97k4VBK74PG0lj2lHwM0t3TKI/1bMV3v
ZJvGj3NzAcRt43u3GRjCORfmwfK4yEl0oDv/yCCv51M/UegdjQuCKvf5xr9LesHOx7jf0miSdGeg
2NNnsNea/f6+vxM+MlUCIA66wnYrMotf6x8qQbH72/CR24XeIeMD35prtLLwN59YoaV3YZmWumkf
LP4pZo9DhlUcWh/4eJt742jhpYzm2NrpQe3fhDast/P81D9ACd5yVdThjsH+BStgwUb6uEVg07w9
VSGryUcc3S5l+eI+umrVofd+QCPZjcMFRRGeFX77uHfmqhevuPxbbqcGJHKiylWZN4X+cKwvGuGq
ixVqTbdZwIR/Mm13tdJE01oY0gtQCYKwTEmADZ54SJu8OHxmFTy8dhbyAUkV/GOtAfVPSbmD+zCq
VzbA5WPab1WiZKasSz6WpGsSUFJ8bnJwIuTqEa7b67hu53PobbjuAZ+/JPrLcCTaPSm2h3FqqJ3U
ldtCI1BmVdet05P0JgdgU5eG2brJBVXrI75yqbZ+utbpKK5wT8Vr+JsZOvbbg1B5ntvA5Zo0OGwL
86/74oIA9laCY5EuE567GaSGIC9i7+PG0gtqyq5EW6jSVQz9GPqHVYzFwnZGe/qzr+kyKTHAkjDW
IKwbn66t5faksM4brQ4sxocLD/T6FcnzAzqYX7BKCBqQidCfDQd0n1+pwqsTPiKcfWCxhHQ/sHPv
MzYS2qQOxASIZc4gU//yXNbfbP2DTffFCtFhFjcF4sKx8CopbIPyjrBeNRZHT7EFFKr6fkvpS/G/
LP3uMsseDQNEzw078kpT9gWYENstRFH5nzqGxYtI7ZtJIeOr2ltQ2YoljC4bXmN8pvEPzDfZifQs
t+xhYoAAZiScZsYonwpftZ0GZY2SeDQi7DYC0+Vd02N+EWiS2pUCAqlt7rMfX3XyueZrTbv9ky/1
KzXaTvb5zn0HivLne+FPBIERooA4FNlSY4ngU5eEP4l9GTcUj3fBjCmR8OL8NIPnLof6vHPXXwme
i2Oviy9LhZ5MHRtOVQT8jFmfE2Sz7Z/vp6tAi9ndr/EnNaFeyajA9U1qvmld8R2M1rO3TgDSd+17
Pq4JJ8br8kebQ6VaKEtIAJsOL4nG7DxXNk7dGspGaZXxtQ39HGfxKaB1qfIheRhjnpUGyo10I66z
xZlj6OHQrQH8SD5OEu4yR8WAw6JpuV8QEjSB5NLoBMQiuGhCESxdHEY1uwL7EFboB8WFSwzb0nbU
Un/2yYX/jrqsaFKXzb7ywGHAbXLwlSpfBq8dMmVpETV9/VgMNgXL/ZXIxV6bGX782QRygKGcQemz
cot0TnZZGGhtejv0KZVFccEAjfxT9pGPZi4a/vJ4pVjgoHRixvVm7Od2r0q8xCYu3QX3ZXIjR4yt
Ww28B28p2MyeBg7hayBrMeBcV4VI0n63KD0qIzBUp+WygyE7gixembISAHb+4Sbecg7ZPfL3dhZS
0/3BKbYxbuybMdB5RGBwmhpvfuY019lwYTj5ipCJX5jha6bswiYi+R49f4IIk0RZ4MtPlbVCZSEC
E1v2gpAJfBKuFrxa/TqWR9xJaEckTwVGP1e5CZSd3/WUTBgP8Qp1yKclrx/2o0XKHI2US1Irnzss
IQUmqXzDMCTuJJltyUSGz6Zoqs6OP+ceO8+9EI5BFYF4pStzkT+NgKSejedHYr8uLg3BZUnsxtqz
uL/D/RcmlJLHNuF4xI7up/c8PoUldhXZcu8bhCs5uRni4AF8fn8OUFfSLBpxoAApdEzUcXf6mgv3
Jo2wjAA0DTn1nJ75gQQk8rMEOwKP3ujhu0knQ7v3Ro/HfTyBWn2PbfEQEEjT95Cjt1JZjdsiUlET
333jhcyqglFr7nsAuYnUm/VB6+ohWPIuP9wij8PUGomrRZyOW0iclMgXkhqfpBFTR+7HlBoTBG6o
PL2OogBIsaSu7K+iKqUJh3PDnoQILfcljdYNElbl1NtPrX0y2kVxaHovx/pmZfyenraEwOnZvAAD
8Gbxb0oEGASarDfLIM1oJY6oYjkRyv/nJC9tGttuGihFwlXKAFOcFzA8bbdNhYTt0rD8pylwOCPN
1rSrJgMsGZ8QberA1KKuknoAq/1moDk0ihM7ILKo7329xBsBJevtq2rnE4+gRUd6G025BlkKTWDp
fiUSCIZQygYMYSWZkNiypyG2X6uQtYt+T2E3uMrQQxXXiZwvpPyy0aen+85napWBtJXtonbL2P3M
ALDBjT74fhfH5/ocq//i+Rz+ej21XWAQtlvnGF4tu2Ad697mJAuhDcEClC0kwvp9wamG4CSlO1sT
g9rdqJUyP+MHNHGvuZ5GDarJUNgLeR4QR/WplsD3MgDEJzmZueeDRhYiEL9eZOb4one/DJelLFnT
jqdXeEf4p30KSvgh/aqlA6aKfkj2+xBOcTA0aD01HNV3NU8d7ypqhJgIh1cd6QJJgNsVeSGK7Qon
V+v8lVp1lVzgWtzm62+YooctavW1/pqeNynWMsozNW8OxFYkJrfz4UnUvSBruHrj6Pwx2DEnWDZ/
mxGiLLyHowKFRssUtc/ltO5D/DvLp/DM4yzSmbb6MwUN6T4M5EgiNHJm2gsW31pHLtON3SN5s6lv
CTumbjtMoUsLriNTzutlTwjtDyZXxC6MqVL2+LwpUzHzYtUkPo6ETIqhDT2dsICUeI3OTJ8RjqKI
4VCJLVH6HALCZTDsUn48fi0LRC+qI/Povnku8LSUOdC/cgWLvvJ4jqk8cFY3RkFjNcz2wVHkdEfL
hI53zO0AqpMn6ptQ7fLcC82fKsbOVhhYCUMFzyHJZT6nlrK9t2T74QF/DCYjba3QhwINHf2/QjQL
/2PxIQrjYhBGYnjg4Nio5N4/wlYkruSRGYOdo4mamIG4WhdFAyJ5etIfdq2LmP5q4nCcs7C1ZJOX
/m/q9O9YbEwjcEpk5onC0jhTsdaO6y1y2gJxF0ET8Rb2RR6nwzPP54jmADiTdYyl6CmJI3kLb0YU
71gsW8g2GpybRC7OtMwSxrjMEN8iYRF+f5j0tNKzcgsW5JMJmpUeYZGqgnedzdPKhqedcwcfB1FD
tCDKAWVSite+ij2oBnouqYb+bpajvWvg0lnlFvwISZthjfx2CPXSfRZ3Htkwnj6AX8x6BJj4oChY
oNyviEYa2m2W8irf/8aIBIwOiMFXI01pPy10h7F0dTYNSM/Tv2dFWvdgqoVXTtoRj/m+p6T9BbWu
Tcjl0i1HS8CuLLk8FNm+8LDHKu7r/DTpNcXjOR4ERwL3zRUAdixvXxoUvbnIcuN+trD1R4zJCKbm
QaHdoIhwTSkGFxPspE+MUDp+IdXxP/+aptymFBIkmFMffWXfCi+LDxyP4ii7j4Rolft5EP86TF8I
9iVEIIbca5K3gCncoKnpcOagtSIzVghurvQVo+PhdqZzHdJI+lV5V0YsjiL2B4CeqVsW2pQYq/Lq
4jRAt/EHZaRps8PalG5Z+FIEGVgqQS/8KdK+aW1ygBhCWSTyZUB0DDU3q83Ng5dDQchTTm8qrR0M
ZUDMMXcY89gwMmrjK7xTDGi5iKuSj6fxrqHCnDr01ObS7OqDdDW/3USAU+Yp53zLhk2+/RNPUL9u
TubE0WQxRIMm+d1aRQjdPRSSimD50NRlsWavvK7/jkj0k8iYtBvwYRcNLw80ReM45qVTSVWpxnjo
pYWNsuccOK3Lp5dTaS6FcfbHN9L4IBkn3JuiX6DAWZB5mefcuSYpsiqZYpQvN4qHprnD69dNqbPg
NZrg1ixIJcnOB412p18MSHde9uLsu0M7cQ7l5isTdtV/Mkiosm5/oJ+EumcmCttjQtnCj1B8ggCx
KouxnOjQIj2TifGG28vhSwnpamD6xPYRV2/0f/dlW0ysIsT3JPtHP9yhit9X+UTJguE38ll+RSMS
MVnwv9rcz2wOU0e0PafJBFVwlqNan0GF5BTxAIsajubbaiBovagpTodEaogSH/pBK3R9r1uYvprP
SMDpHqEVkpS9dFTnHRWp1j2Sa1mlB+odDhLZGrfoRXkwZce0tClvJPLfYFTFQIk4W75ZHaVE8GyI
kzokj5V97sXkjpDLPZtwRB9Wr9+shlEkVdLniwIFamt096MsTWwgvJgrjZJEv5uDY4ntrdZH+Jc2
0lo91W4KpAPnIBQND/52+KA2AlssEC2yRFv4yl+4/Vexd7fb/XJ0Vr6uXeId7ujMQiu7kiDn6VDN
79/U4vUJYJuMXVqxPHGiy+L0tjLah5kRS5SxHRSopBaTgirvA3hqGuxTE05OnVPhLQa2Py3WjdKJ
aKb2Ex4efzF2P9WylAa0Ar2Kie80nJrT19wJzr6B2nOJlSH2rOASonmh00Bshi2AdPzrmVInHzH6
sMkDOXdljDG8StAhWOGIkOEcw4bkp+G+InJbCAjf3Bur65Lle7gtEzl5N7WtmVYxun66sUKg0Ynz
fUnlzlTOXUPWfOAbpw85nYi7LPfJRAsBUOvXsJhYlfORlyAJE8YwrmudjmQZV7mn+P/IDkHqJIVx
LVVSMvLkL+jdMDFAdRvRagoQvK7hWv5zwqMMLqbaq8tESZ8syKRNgv/gua8Pv6Pl0vvOKu9SXh6L
XJrAQ4MV23C7yMZRPDwHPmylxk84GbWjYInjOoJMP83hlfedNbbIugqmkTqhiW6Zld3yS3hJu2TU
rOyhljLiJQAvdozr2KkKnbwgyc6mN86ey7QY1m3S/eBNmheCla+zWOa2m1hAivLJSTK8mOY7r2fg
g1l7qgZez7fT/MWmbm9ggn+AZ2sBE4EdEzVPPgt4Im2Q3IZTDW4GOhasa+m0C/QJNpKzVcpq9+Cv
mC85kgCi0yNL5ZKJvU/RfT8fap2WRPaIg+BZyVx66XzjGO4lUlfdWGkf1h+lYgplfl5VvAyVW5NT
+2Tbx/PycTMzc6id9EJAhYgi80hzS8ubDgl03HgSXeuIOT6NAU7COZ1L1IZTTxlRNKhAsYPUKtL0
mTDqnv4/tJu42Gnp6qq4y4F3SjscXvoshAZOy2C+lUcwLXzz68e/Y+2hmTD1QIo8Z92F8laSHm6m
/jqBb0DWX6HvD7DJ7eYDqgAuPJdabZEcUa56SkU7B/IzTqtXG2GOSwq2DcTV7IWXWztsD45WoTK7
n7IYM9dvdxzg7wJV0KDXz5fUul4gtmkz5QyNOQ8+EXsPH/DUaJAPH+JVZDJ1QX6Fh58HQB+jTkPC
Z4WAFPjuaUKiOH17fNFSLOrjIgenjergGEbRaRUmWJwCx5p5t6O2C2YxDbbUhfn9sQiqLDdluVAV
XjhxXZa6P9uF+3Exh+6gOelkSCumTIlm2/zM60YUF3+JPiGyPcUIUJoYUlrg9VoY87pO+8TTio23
LK9f1AcNRi9dxHj3pXXyyhfrp6UnokwE24VVBgOMSznaz3A3YOIaMhVKn9RzaxRXrE5iiVOZOnKX
oDnFGgWTLxyX7G1/H+4tOkagKfCtLROI8obga/Oxlvc+QeEsrOmrAUkY25RoK4GLzYUehI12FvGA
pjE3GWZvsPKufTwg0GN5SNjraHQjpDIUgxfVT+zjkCWxtLdqqaFEdDXNIvay2FZRxlx7nHAE8K32
U4pAMV+VQqfbRub82kkXpsIasTEP/YZUMF1wA+qU0nRcfRj3HP2UkY+q7GfvtWQPwV+4lG4/9EZJ
ydrooqMBkCX0rEjn9xQwrLUwqNbcqd8ygSHmfua6etzKbXU9Buiw3A13uu9kLO4pxQoGlEYUA+zL
sl/5UlVOKxxg/f9KB9cea6S0zGkxst1S8WpaCR/RE3QMtQfGmfsymS9mwbZGdCQjHvJXlB/u1TNb
kA9/KAsZC1lifSaYJqWQDOszqrzCyWBZQISneRaT0oRqyMot+WaM+kOlnu2TkhSzlyOUVvx/qz0t
K4wwGssiOzo21daNwNVR3wawjb/GlbU4Zk2sFxk2SRFFsWsuBifzyCn37QOc3vn7sq9WfrA7/NDQ
Vhc5E3blmTE2lXg3adOQW1wq9aiQ0RKCWLPAm8LTThQbwlJ86diMNKlxrQvECxHnSog+EJkyYsDH
QPBMCoELF5jMgI5tXltkgGYin83UnSMECGLSwgscyyTPutWQbpQ7suYaVB+crsyyzCqNOAXyH4Gv
lpgO3hEVOZvxKYTaO2+MfcT4B/PF/QP0aprEjns3TbQbE0eW35lTKJiilT8hVqw9SBZgFYM4+gQ4
ah8qjrdUqApE+ZsrOTkEkrs6r0rN/OziHlw79Y59mu4qm0iNK/kA0VuCdUCgh2ou372SPiQfWY2k
mHbXy9riPOSPIEMHm65TuWIaXK/Oix/KzBEW7WhfDEOQ/YhGhjEfAGDge79yhRrWmhfD8zQ9lAKB
po44VVQBOMDVqiT6LyGHou2F/RC6Q63Pcra26dKyFva2rBg/yz2g9zAfb5e3WLlTxxh2+Tp7Slj/
NOChosUnfYmXg++sTuq32zLO5qVVDkVDO1yeZf8Y8ejG2po2V5HKnnVyJDyjAamxpbNmQqnFiKEM
NWDfkw/QxI+/ou2ZrtOnGJTnjY7Y1T2CKdgWweHcTsZ+5mVZfB32EshGtTywTkuqR/O5uk/pXs3o
ZO7/F9rOg6VfADM8/budstwGaOQkWeA+c+AenjR6BjtmyNgdGmzIk8VWIp8/ogd6zrDmFnHJpE+W
NWi5wIwwL9pOKRbHfNYdqFDQjbmCGut5yjCgSWcziiVB2ufvfXR7LNzZiLBEAMCe3S+SMmOEqNbS
zp3tMACfI7AyMPmeK4IRu/UyXua6wZf+bugg186Ato6yU103pS3Hvm2+LooYvFO5KNAjyULgkPRk
8No4j58xaJMgHKMc8HFBWLkJIETsEtAOpWt2Iyv5/mAR7l+K4sAQ0k0n5MlovWmu/DQ59ICNrWHr
xdTDlWIjVqFtU2TZPMP2awJCnFq37+3uYNpf5II9YyzTiUH3l3LuLRoLkyqZREwH7huyIt9HmNM5
o7+e/FBKvN7su3a/QrFVJJhW92sHZ0vxeQHCr2aAe5y4Wvjn6yrncci1dz7pRkZ2hkgb2VbsEWsl
ICyHxWxyc1fGnQMYpQ9AYbA5TE1h5DMuLEOgqJyjDaqay47K1LhKllGMY5cbiQFkNKiNgqqWYtJO
pyTSk30q73GFNZJq+isIB2bmHI7S60G/O5Ou4zk7yWTT6PNAJudgWzNDi8TAErLNxF4XN49iPQ0Z
PCHQROX/YJW2Dxr6iGFhs5k85fuorAD4RtzHWg6JB8p8PZktoXSvynBiDdnS5QiX7RgokEuNggMH
eVtRCIFTZBtrkitEsz/qVqnhVTkoQgxiJOVgowJyfZpvyWiNGWYD76dwDC2TNbYoVkq40/dLLlfu
AhlPtl0qj1WrPwNAg/uJpghIh3DLlyE3sfvX29LeNqEIrFj814RkTjzGb05JDllxZyWDej1HYyv6
26OetLXswkOXDS9Yuz7XxTn/X028maFS0359vK95wFbdh2wa0EI7+mlv1DKsYJoxY1ooRh2CW5SI
fDBmVPizfy3Z+4pS013TKhflE2DvamjRjx1Pi9cmQIfjykr+aXK9tWOzq5CFnEXDXN3vpGdLkFPf
of1RGrAUB2qxvZPfk2aKwEzDOAIZB4V+f0LO53B4296mYll1tP32he9QjHFIVSaRZGlhN7kr1sR2
RfEWCSgg65vXhfaGN9luoYrTFkuCnJMDV4GKMIFAM4dvAsZ1QjvjGhZeC3xhu1VLUTygnwgqJy2B
C+q6rLDQWUSEIXtzaXwrjPz5Hn5/p66glyNKBe6OVmL2zW8J1tILyY/sukNlbhTLHWLkGeD9+yUh
Y/GNd05qU6XhrsdPfHmgeFV0vVfw7O5B+dA/DASYndUuMFmiMVZDHgSZSTBx4jobB19k97sItaFm
kNikUxcIovhsEN3NYQSzYA6doYUtFiJFjmvYKou02r79AvMo6v9BhnViT8oXSQOhUVkRspfwbLaW
qTknqzAPCX/ulLOKkXik9l1km0Fwe4eHF91RKbzldn9KtgLggqHEKju0jsXTvGo0W5pFU2/Ea7/0
WVjmIR2vMxqURjW5FipnxTUd+ZVw2WosUNc3tZ59yMKk+b6RVnFVAZDAkv8usifLi9tC++ZuWyFt
25NEJMLYdh2z4yEntWL7cpuWn2qMlZZN/ZRz8aptNXpnz5Jf0OUOP4cvoHasI+TTopitEzeMgBKV
lK1dtq/JE65LtHT0SsOrpi8V5vgK1bGmZcJscOHc2qi/6CJq2a/sscot/2+RX03Y/uqChXPGNny/
GcNk1ZkZrCp4fzzN4JsvUrz7KvbjLYLajjt/Pc6APmmCX1ASC3ZQ9cOLNjasaux8pt2JI3M8mZgg
1G1MaitnK1Rxo8zREHsgKXRCc8S+0VLa73beHLUSbd682v0AixXhY1/Na4//qWRkFycHx1bfu/pi
TuIfPzIH/LRYZzkozxk1ymx+WvaMCPU+SveVA6zI6fAhktnLcydqEfr7Rm2ROXw8LbNtsfUlMrPE
vQPL7ioGlqOHBbSa289PlhqbTNHoGrjxZgIxmNtlBKG8qJ+gibs+2ECWEoKYU+z/EVrXkRx4O8nU
moGd71jlcKuf7kezelyVr75TDGMisiK65ErkChTnkqLdbXHu++SyHV+/psKXFS6nQM2u076Y8qNv
Uu4/+JJ7YcX9jPQkUWawVBDFSoBxXw7KhULzNneiCEb6nejjb1NR+riQTmZx5SSkfW7G/CaxPm7s
JD1rogGSF5AX7+N+DGLT6fvRWqhkQvw4dcuAFPR9UvtZeaBh/2876ShEEAVcoVO6zCJORaPegqb5
zLAP0vUZnYaj8zek+HG6OA9jeKnIzVj3/NLAVCZ0Iy/fBvscRn4aH7ox75hWDTLzrgUCIEzFNk5T
872kgQ0yU0HvyjF26kjHfCR4/K6kDTwGCS5O9F1x9xVisZGiquDohO6ZObYjYFOo3lep4xlOuOKD
qslCLYE9pgUjqxi4ONwr4WyWwEOhXBPEuZoHiiOcOIjFaDdzmePUn/TPCQfgcUG+Dz8XCeO4pOc9
bMYU5GldalBEjeCclKW5miMppUynNV2+l5vkpwjJ1LnbmfR1FwhT6BXwXo7V56y3Qvxx45PKE/KW
fyAkPA57O5SMYgSUNPPCwh/sXXXb85ULnSe5NW4gBfeX0TIEnVsP1HablBPkjS3qCzck5oxx2azM
OW4JXUf4mRwqq73uHZKPtlpC1hku9pwvBiAxvuU24R+A5EeypThXa2BAEfOpYzfMgTTy8M36rilA
acNGefUHd/zacK8IvZWoqifRCOzaHuIWKMPacPIBNownYAZPwdd66w1fS1JmYWHks1ZpVoFly5z1
ZCq506CZY1PnDeGDO3dRZI3r1a/P36sbY1SjTtYZkREYHs6rpSVxIboo68mLZn/yOhXSW8Cz/Yoj
w49+9sqYTgH1DK6tscpy7bvczTK5QpJNBH32GIFyvbEXxjSnwjIJuIvm4rYwqf2gRMLBCa+7sku4
Hq07HTG3ryaTIsCsQ0KHp3R+ZZG2ZtAqQbJJlVwq9/lS2GvOnm7ZmMsprancKXkLuAFHgA8Rxgku
q1CNxUxvoKO6wCB48g15v/qlZGb0Cfh7myWfri7PxNA0tPeAYRJU0/zT3/C189DrGMEpNoBSLOhU
j+y/3RcbJFpw8eS1TdKsbR3gI06KvgASYV/JJ6TxLrqFmKsE8k/1c0jflOUSxMM8CQHzRk5x2iMI
jROVN3Is4zS/Uth/kn7mSsIfCwyzAS27hJTeZ1OWOZRjlUI8cyuuMYQ4RaAPR0NT4kBeqeCBtfZt
JMitQQ/wA8ZrOaSX1p8L3k+b+FTYMe/mIO8iPVxhq9bIpGWQQrkfBnLkwzY6xmmMN4s5+W5Itg5k
xtZuEZBRWL29dOhUTbUS/CFsS7FUoE7nB5jOedixkdhaBk3VuDcIucMeqfofXRgto3uF27aCkUca
TOFJUdeOpXui9M5m7Vm3zmuN2xK5gpDBnjsHYHjAT8F1BP4sqsBUmQfLa63pmj83auLgoowPDAfE
nS031PyXPJQy7UhgJh7HZxxdyZb+qOO+dn1h4tLBGOXjN522CR1I2DKM5JqohNdI4NEbccA3JroT
ARBO5gzTwXych6wMeAwTMacjWrrYQpwHywGqDETpUhcrL60ed9u/+P/jYgGWeIBMx4/N/tNA79Mr
osZd5QJve+nPvv8OJkqKX5inulQHLOeTSBGKbtl1rnA5piuv42Ji2yE2tZjj1WFIq5Rv0DkG1GEv
vTxdVHQ2EZsXtP0fgTheIQ52BIKRK79/CvwkJ0mv5VAs6BggK4yGgH7lHofz9vlE10yEV2QfEsi/
kWLdGFf7O8flHuUMUeoh26IPWLHMxqZLioPzyu6ZkIQtqseoBIJebxLAh7DG9xnqCtuJVzCO1cBv
x32Eia5OKHLcSiRfqml0L5dPLzGTQPBuMZ7iHyUD9p438Ml5fvML8/g6jab3Ags+GX9muJXMV4Sf
3lWdI9sJXmTOwf/fGREyaDB3Li+MzFeBMfuRQ5cs5UkxT/fKAtm1/8x1/odGUQ9FbCt76feViqol
rV/qdlZgi4+RzgTIY/VwlLvsnisPzsFZWBQU3eHQt/jxFiPkhbSoxk8jkKaOTH4iTm4Y7VSi0I7N
Nm8I+MTOSZiVGsdH8tFUOcCuyuOweTck2Etyi2GJmZHMBXb086eVJ6wkHB6zUykizJVIN/aewOHk
C12CHyO7TTlZ8BTspimGq1/2t0QR0Fk4VmAc3hJXeUwVBtqU7QVF18RInhqK7KrEeFF5xtXIMRRF
iW9YhOP/j8/ZHCtKAAE3X/JyTakNfBL8pmVbb8WqjiuFZK2nEOVhY5DDMV2Ng16lIa/LozVjTT34
HnmS/GaKE3o3NHonaTEQCUeVLJLKoQBDqCl8R2hBoiCiKdy2ll5UXaTNeGFxI2fc8AvLnoXpWqfB
Klyul9jyqGJGryzfyan5OG3nnFDlItYb19Z2NdmwCz7h7OeULPL1cX+fdnQa8xUWLVDXe4UTlcXg
uBr5gVSNIVw/0BJfSdsx81oCSPvXVdO0nFF68nZ9qokIxUUHxx5/ODFYEDtbaf9ZOMN2c4vEKYPX
q5A+oEK71c4dpMNQUiToewTXBQY6dQPZxFz5Z7pZ4hNMbccEAU6tpvwSuLIaco6ej8tkMi8uu49h
Y46ZVTOfkTX+4GIUFdeLAmFGW4gxR3zg4fNBxuF5vT4wK9MqTpRe8HMlxLQO1lsBZPsVQZNbFYea
n3Y6mnuyWPjeBaGHUp2F4ahLLe1tmZ9QP0p2RPbN61X6RdIt2H93lTIj78qFByBSGVg90kPMfYHc
dZy7vd7CCsoTRf4n4loJljiEQYpCAyxXZCJxjArlTkXgaCBC8evo/Bg8K8fvSncEJ6kWvAJHt0CO
gfbJOaKvxaKbtddMJF2N3V/Khi3J+/JCI5TiPDmLGJOi+x2GeEBRuAVzfnUZNbGa9I5zCWqdR+2D
1alGd4MA7N9/6pgmU3Cxdi1M5AaCL87/a/yYu9M+UdJZO9b+9jEnrS7lzwt53CqmSx0R07Th+9aw
OOm5UkVO0IzH/ED5Zmm45OdS0RkY74TkHsUp+QfMmcJ6shzMogwzWnpjFR5yCxWy9G77mo1wnaJL
NevUdGfZFiJhXlicoEDwAgGg3Ltn3p9zjQZDQUx26NGsdE5h91D9wTFgkWdMYAXD72DwzFl3c8Ww
y/6OwdLN88ZOMnKhtsXYhEgA232sgW6kw5lZVkK8SBY8u/+AhCynRsST4JZS4zF4fA+xT/zBGuaj
HOTvhsXjNPFOFqy63rEfvL+099Biu/K13VsXT7WwkR0GX4m5SquTzTNkcq49uV0gq/VxC55GEg+A
5JqPyj5Qr7h3ujdXphSvNElzjBirxo47wwzvEnS3+nvyviA1Hyw0SdxFO/DgkH3rPeYlvoLDYoyR
7H0JBDQ8fzW9hogtnB2ti4RRwOoRydDPyztA5q5xp1c+NPm6/8FUPVVPlYudgzuz3ntyNvY8HVTu
GqJiGNS3oEQ2N2A9qFhikhQQrotfA0WhLBqr1pN6ow+nrreFOZzxi2TeO0A5NCC8SKdLreouJFMz
VLAOYgNl2EH/8lM+vND3To8NcQ5d+XojreqobCdJMIVROh/zlH/tP/ZrjvEEFleUG4qTBtcDJ9ys
du3I49Qzief2hkbSz/Ke3Iu/dSI1AYd9UT5NK/aAn5VT4f9ixOWvhFyl2tS2z4TXTvEWF6AlzBGV
nshXAy819KSm9N3RQ6jbgQuvnTVfvYZGllh9RVvNpXNGzJhcezQixTkJ1kndIDezgjMJQvWhcSM3
r1UWGK4muQgjtJv4XE0/SwvF5olZSb2okeyDpw1QWTkg3/LsemJjn8IGRUDNeuxPhJrioTCOnP5r
hVaa9UUgCXESOcLdxcn59syDMOxlA+6yw18DIVTtkNlrFzt66j2gkGpnDq+vfY5tSTnK1g5tpqri
cl2o3tkRdZdAYixZyBbWB/E11aH7sc8/9TWbyZ/w87E011g8n5WqHn63BVvbQmUdtsetrDjiUlyJ
t5vBgU7XuQoztlmxTHbeoG0YAP+gl8IcDAurGnYOjOgwRqBa6sKxK6B9oxPe8kiNP9wIdqCaGSbq
3uFYseK0WBpx5C6wtJf0SIheQas57xCxec4n50MzLRWj4OtmheGG9aSmQp4YtRu8qIOWTbFW0NcI
MNt7W30tyQcloEYx0wMmA6g21raDfYz8+BVFoswX691nGxIl0SjQ5BLDCR2ewn7o7TP//+rOzpBq
6rkc/QfLRXxXtrDlcC6OCP09jD796WK6AZf5oYJvAtCaUfGfYkIm8BrBgpFwN0MLZ/tPSlL3E9R7
NzI6PDDKdf9OKN0Apm+QhspgUMKmRxm44Ll9s8ZGEJ9JRqhOkD1cNAdC88cdJAPMuuWZU1wHrIH/
NFAB94CsmttvnUh/ZoMFOFKLTLPaouKpQtr07+PO2qSQvu76c5F+CUuFZhBWDb344WLCHN1eNuYP
1z6tDvjlkKvveKoh6h+jbuFJqJwTTc3btz0JAGSGdgIFnJsh67GNVMxE3HJy8SIa3SVqsJ7u/7wJ
Kguj+/PDOvrFE74SlA4mmH4Aup2hWA9TqIK8evZJnqC32vmzrvVSFjrXe/ZA+95bUccSk4WD/2Ce
3ddJKq0nU+OitdGcmC1M+wAHkN2kDgr40ddCUvBOJoyi9L9lId2sp184Born+iVUHxRtnf7h1jH+
GmokgZL/tKHZ2690nRlIQtaQ0ENlKdCbsUPGzq8/mJZljcN04lWAk7sPbdvFgSU7wsLqT1xH/2FU
Re9TBhqcT1IIkdw8jIRF+M7ZbA6H1WtAMoT62w6SlIK2PhQJMKR0smpU33MYDnYTOn3ESKjurFjW
yIhpF6P+cFDk3IXei0QHwoylKb4Wn8eQr9tpUFJ7C1uNrEKZH5oW4X7zzr2fQOCNtC9cRHmKW+zs
S86jOK78N+LZqAbs3kMP48Xa3B8HeMVPHl1WsTu5Lkgb0uicaIZfmDVFlfwRUi9mcDTlbqvyHgzR
boSrL0igD1AlWxi/x/Frc8S2lQmC7/vZPzGqVDp6ZeRe+8D1SdSBnQVtQMoocAZugSP5UmidfuXn
ZScF6VjnxSQAK3gPYOTTGyjH97Oi6+cE8Jc+iijD8RTvPQICCHo9NSyencZMNPwNr/euS0AtPdkw
nfl7v3vJjPjzHCkaE0OtUSouelfdkLVmUflD/X3gCK48tzJxjynnAB4/qLLgHpyTWyOf/GVgCZjm
8+d5PgLsGasruqOnK2VM1SFKq2ehQlorSY+9WvDFo8M+8NFfAoV1MbaFzMmmh9+vWSuSdXqzUoM6
SBehBe0hbdOsAdPtQv+070+WZdgCnzm7YR6d5P2CvOa1UJ1RNFXoMAyyZSRqF85aq5iJw0MZ60BV
YccnjwN1CDeFLc36SZWgxxiM13buNA3NyDpCMVAbZut/DBo5vayPm/AkfRaatiKDPCce6FPPdbsA
L+pldxCCpuJfXtYBu/LS27KodjUU4OsMo/knb02wv+GEqTbfmUZEIsxTW6Y84tOzA8hhADCLyhQ+
S/x1MODQQWsU9MAgKfxLsP3VUyVprKksqDBDKJltTDu5N6w9/Ttxs7lQ9Qan1a94rI2diySsk/hR
w3VNYgegvk/rCogy3j/DLekV3Dj/lQbW0Soh+MI+edGYIn2L0fFGgLyQ6d7R8kEvJGIXfU2Vs0y6
oQzQ8i10n8fKPKQzgjEFBxYqeJsNCHaGDWOSeKY3HJLXOECbcpiHl+0c5r8IcKan8Yn3KCTVI9Ma
YPg/o3udmOPXJ9JQgbzxwaKXf+6L8NR6yBm6NPI72w/U7/7YqEvauYvwRpi3V9+chjEeIdBUFyYs
SpgV7bQmAjBl2YiGuLWOt7qYXTSiioVdxO8s84mgWSVdYR+v8E1uANOK3X/OIXx6iKFygAJ/POHK
WsBsxtjMo+WkDDVe1W+VaVkG3RZ2w8op8Px6XI0NFbTSgzcL5FHBP3eyIA3VFD2ep6yrnE/Hj77P
kPU0zdF7/+YimfzW7ed70k8I2kf+BPrhMOJEpEV9iiubqBSIZQQlypI9iFI7eR7HMfvNlizSr5vB
HL+sYx+h9yVHKox9eIRKnCUr2igAxJAX4DEa/RNItMa3geQj8ugo6NlvisWI2nGwNlFbokoLd3vy
xx77jR8pFlu85OeWVl/NMyZm5txZgvPc9MmeFQ4O2ECH8U/o1k9yiiEBrBTy2dxLa3v6zz1i/9Pq
J0jmefsnE6EhmBKY5U44FKP+73kEelUyxu3gSIdGTLav/TbU46IOpnZVhRptPsgFqqtZMee2W1bY
KQBM0nxkZbd2MpPFFMcSIfP6V7BGr01I95Crjo/7H/aM/X+iKgj9UJ9Mu6eNW2HiggPLy/O7M0xa
J5PWaD2SN6JdeN2vg8Nz1lP3eKWxi8vlGIEImDQxvY8MAwm6JjtqZQU6koljm3NrvFc7jLaMZEPg
4UmoHlYtqs4D4P4Otry90HpdB9+qP5LeMso3s8th4qSdi6R0s+e51eYuQr861ioXBh4SXTVv+jye
RXXqRDcOUpFBKaZx8UcwSzv8p5513ywuhTlBz51Fh+7Z4zHG25eL7hfbMC4ZPZIDBeog0OMeHe/g
OQvKSASVxsHk6EC0WiIWbBRqBC8cpWKDC/U13/OBG5CMlwfZaCISvtGyTkCU2IxPvYeoVmlM3z1v
Ll0fzucHJjIBRIl4wGr7IrrVbEO+B+2rJtB0uikoDUWLDZ2nvLUrkii3NAMOoTjxGMu2JnK6uBxn
vYnh36BosQ2JkVMtm557S0hFzYcSXYvoshylHAkqkUVYtg4zsItB6yCPkXBEiFbiBAKmv3ewSW50
kSVTZBu8txQeLlwajUQ5Y39OLKbGEGZaZtFAt9UqRPXIXlTOqKkY/mGKm6RNG8wHlhSjd6Smp5eG
ZxsuUX5rFxhAUZ/3UjEGKMapLNGyitudUyz7hBEmL9XYttBbaHl7kaRLV8XbxAXFuTK9OnWeTpx4
Og3fxvjxH0UNUAWF7gr0Mmdlcf1ujG6V3hniCzwinno88z10pKTikZNVOnD4Vs2VW2uW6OXwEnov
SrRJQaPnyJvnTWCytYVWvU/GS1re/PIP59Nsy6oLH6F2guNGBa+so/LLqcGa5fWMp6OqFhVsOrMX
udGLaWAymy3ItZX96124a+ErfjP9tyTJ9FQXPpo++A45A987/cwrCYa0VVDPKHxMLvrRacyvtl5E
nFiF3HG3wBkGSWraLSqg+4tE+ub20YIinoxU9C3bUpBAYc2qGiYDzz1bkrbE7nddUFUPM0Rn1o0K
fdCR6CYYVnrHObJQp0prKoNFwPuyAnCDCUCCKWSbcJ/epA4nWP2m6c1laoqXOW23iUzvB0qnP4Cf
2HBlSCdU9/tgOSv7tiC68n7XYODpwXor6UNxElMw+grUEVknOQXr2KWThqReZrSlppJEHZsG+rqR
SGirRSeZRbPZgYtfY3bGXL04CC5ZKF6s++a260lW6xwNkb98B73chvk9uvHIZkZ8aMElXiQVzi83
we6t0klihvvAXAzZ8Ni+ALCAoUE+64m5e1NEm57g6dTLCC500VU7iXqDXeJ2N+5xCGCNrusz0nCZ
mVE10U6GMMIbwltcP23lyMFgAxgFcxSFF3Xo81LZO6A7QdFuStFFxGoaHghH2K69Nw5nHiikFz+p
uxHu2urI3f0cfJdTfLkQgIgZNxuIxgfI7K9lvGnerlKrnKXePJ4mM4edryegL49mB86Ey+igCIsm
/sFQhISagZJ6/LA/6mbOEdYfSD0D0JT0kCseghmquGH45s9RnIm/LT02J4bOa3xR/EVDamnY4vmf
WUkXDKxrGvTMKY2LsyCBu1OndWfz9Bm4++6IwWhAhFF1FkomlnsVNLpztYQdTYocAHY9uuyJQHhP
Cs790uFNOqKRAh9669FVQ94gjAS8xW55nWKW5yKvzZ5NEtlM4n7mHmmEuXBDsWGO3thpBfGLCfjZ
Iom+AXZQU8zOPJdosLE6JbkYlRCrSzDGYznlXGEGaW9036QxVwCu/gf5hWm48OADtIarAsVim/ES
AbITafl4H13+Z877ympNOC7zkOE3iKt05dIsZkKQ35G06T5iMBU4qJt02mJO2VOx0x1oGWyJMHAf
ekLxukN065n6ZxCJu0KzmTOD5CGbu6hPICKpbqE/PGsEdEhh3MB10vS0qlrJs9pV3v8TSCESJxuk
7GH8Wv5ZRLLzpmPnIJPQZuoRhOVfzzSHghUWgF4vHMGH6rDEq7A6MaE1ykq+X/aCj1ixGzQCI/PK
F5HlLhpZ49GEDHIVGWJ/XApmBktUqkWbImOThOHpBMIRZLZUUGbYEX/gCRsw9zou1BDXSAyzXmMK
S28cYksY8uXZoozOQrxanQCaRqVZLClrVLGmvwdP/H+yk+Zu7FJwsLw82nSCRL+gCbgxPwLEqqUz
KAL6fVD+l7JoS3WpnN7jrGEg94qHE53TCIZKYxVmTNxNV6jvl2Zwr8IYfgeh8wLrgQHlSydDs2y2
+zNGcbRTaSgoB3i6c4kpHpY3uqJVub3WjgPwrEWDZZmyA+H8Uz8a1sduGTOvKNn6rP9NJp3t4W62
yuZDds/fd6I1EDGKHq1qD1G66v9KPz3jdPW4ae09rftovejR0rgYDQzrg859v0u/8LGHkRL8idGW
XmIZsrIth8nk2qxqFlCDXWNOLkwZV7HbC6TIeaHvEMxrz9sKao8I5yUDKWGD5TBBUDMk85eki5bI
u+m2i2MPh61ebYHEtAewzJSguWGSGHyhhOsCsbUsij0p0Zuiqp0YbRHxldvosj/gvaq8Ls+Yd44D
36dZ/RgjRCPfToRyk6eXUaJnGk2WVFd1jPu5Vuquf/nCS0stFoWNylbcDx2gYjjgkB+wqMQvdNEV
aQEqTtBu2GAj6pmIMV+aZ9LK9wXR59tryxg6tE7meprAWHmSSWOAQfGSds89tMIbmwXF6taZiWOm
PJjyR8hb/kYZpfzUXJ/Gm0mhVeRRHyskp8FOfwSZRCLZv7Has4WwJ6UaxJ33J6J2ynAlCy3n/osI
2yALlpDRcgdjgE3M2cGNcIkNle+ogGEc/16x31MpUITauc/lnKzlGE4V5HXvqFP5MHApqYpHWjcE
6jvjqaUPl0hIbX881L18oup6IHJNvjAHb7UmDtrRKaJyV8HUQyeD6qumCNo8y2nDwWZKwkDUbZuZ
VVAR6w9EyydO27JvsGSwEGzcl4P6IchNk0eK5vD00iDzedDwyJsXBwOkB4ESnZAGz2znaalgN+IM
Ag0B/bZQJKz38xy4rl0WjTgvhivXAK0FVG/tgDjjMsiD7rQVipKnuxhhfDnaHJCqYRCPzflxWu1D
EKyeB08lqs5WIKy+hDCF1O/r8Vh+/hkNKjJyPOTkqtDKZq5kLPX90JbGSFHbxO6ejRA9DFUKhjNc
r3jB0GmBCbbvhQGqZASLGYdJe2v+9VR2+qEnOkcL+VMF7G+YvsXif2+7lqtaXNAXm1wXg0aSJ/Z4
MYzcvomst8M3TQrLt2+lch7TXgEDesDYoUJLhygV3L2LTkCBchUJ7rsVG2MBT3Sxe7uKV6GJGl0/
drDQTHjlTKmfQ73TaN4N6GRHTiGT5dkI2DygrmeVVJbUkzIGmf4PLLJiGRaHw5vNcTMrK5H0L8ei
0WHtHuzpYDmYL8Dux98Lc5Y/zMjRadnyj5gCQADkIms7l8eD9bVu68+u+l/pFdv08nlBykT7lMTp
zjqO3ILPMYNn7G6QvUhOMPy5zCT3KMXQLfpv33WIbrTytYZy3aPxAlDj+xO1BbhvD55TOKfZyjHV
cYcx6JDlET1xgzzerMJ6S1BB7L8SEzwULW/B2b9aM+nlGdFPjZeQ7idtFnQ7NliinAXQfXSh9wFF
b8HO2jC2fP0i59VwZUQzCZrcXGc8MEUQAA2YqO2rFPpGQ2+/u6fEH2ZQltGhuMZDrVIWt9hAVtCz
QccpfslaEnKGvp/c7WofXnOiwfisX3v/3qBd2ydUpzpliQH0vDuBQyciP53JNYYl6XXF65aZ+FO5
sgLILa7g8Ozpx6Eh9g3xDUyBt1oWA26aF5jQUpdlO/Gkd7CIurBgKMWd56ign9TibKl+GovYnW09
hXC3koY/RuxVmxixAdLsExlvuT1pItXIuvZJmLI2IgLyxOEGrLlx70c97RidapuWRSrDafheA1F8
gbIvmtuoGLMsY3ZTRMqp+r1Z+qZDdudNQx8emzBLSagNb6UpLEQTTxKh1I/RhwEJxPNN8Knm/ruK
SeoNJaQmFBiKrW/jkfhpkOhJmth7cds9Enhs8E/bivpFNTdag5/cebAKjxwO4rNLPyYZUG23lwus
DN5Ngr7Oc9FwRLOLms+FKnilNgZYXefr5TxNGAdhiUOMXv+YBmv/DLWXFyVEq5UlmJ/U0Fx0rFe8
KviiDKVuro5WqklMszOCxtMgOCN0W8Ir1JIAhxowBm65BGco/2m/leCWM2ij/BVueUZpS3Lt8if9
4InnaKuXxumk3sMnrPgEor1AqT5tKQnVngE9425xzL+PKc1GvgN2b7DKVmMUynW1f5Kt7I+ONQgj
Vvt+CmBafgHDcWOqkbH/G74H6fTsdyl20qli5A50/HCm01pstQbNb75y2Z9h1m7GA5Xx7AaCaA+1
9bY0nbLESpgiwfIg0TSJUb5rm7AJdGFQ9mvjG9t0O/rAgAb0IAhNNnyh4Smo59rOdsw+2mDQOdX0
RBZy8mN2wq4gR9PjpCQzbfq9ys26yCT+TAFeyPmmAFefCQur8FRHOkV+bsepkHrpXThvT0vmtt6L
jLult4A77q4+e6Dk8nezT5PLrSY7EAXuWxWEoQkptUrF6KsI2QiYYpif54Qj4omzAdbe+N5gxUgm
oQ33rEiz/UWiYiTLH/dRBnNwgoSqQBSIac+O1o0fSxYRf1jlSZ4JG5J0zBspGk95g07DAKQrJIDF
fhBCIyTy6Yj1ooWvQv175exUbmFyOQeetZ2il8mRKRHmVe8VCIM8Nrj5oFL3g0Xca3HWOdinjUk4
WJJcthnUruMVX1g5PG2qWCoK00QzGl0yUszXnI2Vs/D7jWQXWfZTVxGMWGBrDcV4COs17S+YjPK2
wUSTHUuuSssA5ots2SFy1rfftBVJ3VRHmLaZ/VbOu58aLISinT5RCEgWnjaNWKfLA9F4QRzBGest
sR7BeDEEgUrK09BGMfDvT7bJNIizf8ipiZkVtkJvSWAqhp13u8K0kYlcqyZ1biEwGL4zbIdxexdR
Chr3yeuCi9VyHKWTaUTLWDg3d/eDJ8rkw+sla+sTQqS0lyk4Xg5X7It/YJTLgTy+o6fHlwQLvIa1
fOWfrPdMFHfJkeEv5DRQ0R+wQazLavO0HNyYqwK+O3nWOTz2PTBb6xtt9abQQJd3oGHaF4HvNI4J
5d9X2hTYw2yb7LLkTZ7CIarcMaEk+IApRCWIY0pRS0oghL8cdWdGU1HSTu6MUks0Rf6CBp7zMQ64
biBExIJv6Z4nOWCUdcvtXeyFjSoY3C/9OYGKdqIIxu8yXORkyuXkxAGDySu2Y8PRl+4AZOnNG2D1
mrOkzQSrBit49EIdx7oOZaEHpiat/y6u3Q/hBNIvibPx9urvKvsp/xJeqCqHeQzCscTW35V7Dor2
J/CBfRlQBpyylhQg3sQ1/CkO2R6Y5gaD/jLGh/154z+Wl9zb7VszAUAPN3JHgjtLbB4dqaUSzDn2
QxPzPGJyqTiYMEW5LkxzKa6topzK8ePieOJODysLFbEjzfljaqIu9FDnx/C6496ZJJBG7fXTJbm1
chaMDjVmyUSCC0vVKUN8GOZZTlSvs3kPmqc1N8Mo5KUIRPxzLXfFp5Jz9GVJHoGhzc86LgM6wckp
P/VN198cRAMD3z2eUwTwgMY1I2gjv3T7TboiHPrs1StkhkVBICk2pvk9rpaZEne9uJmimr4mqiC/
K0ayxXRuLDtiyDRdosvfHLJkLfpRwhQfaqTtUFzGbK1neFDjoEzgBcPZ5ae0Sek6GyBJfjXo/oej
LQUTpOKyYwmN71VH8x4XP2p//2AfBkFsGsu6iJS0tFiZ0kkit2XO5dVqolqqMh/XIvM5dC7X3mTD
YNgpFlNOJZoREff0PbLP/Npks27bbex/xjKcsMXCVkaQIPmqV2rrtHIKJzvZzyiS1PYH5dX43xCp
ran3+d4qB51S4kK2o+Uoo9TMGSvcroX4Ml/b60kIwd+yOXmC4aeBe8iLqaSP/3b6jizgpR8Qmf41
ccatj57352gmh4zZhvtO3StfdbSPa9BRxh6Q0dgN29u93uETmAqIQmkZOHyyWfv+BKWliC9n8Bnd
fABFMj35VUQPCK/I+SY6QKlnLODMNBK0gcINHEytOIdmdk1O0UFBvraauZLMf5mJ2a6I7VoNNoTw
xigeDiEk1EDyCeoThBTiRpFXQXrdOoVCEnIkvsKl15Q/Y01kUd5iyFZEwrWyjhYJv6GD2p7VuXQD
J83yoNDkm7l1J0lgjRFE+e0vtHB1UHGbcZ+AFqV6aPufVmLbLG5JazP5yfoMeZRnfYp6UlLPKS9K
PHoZ9Js5Ur4EnFv7sd9tGM4v9w4Gmw0rE1IKNCFgqs0KWgXhuwAoopUmoBAilENiGTGp7WgZirN0
SRA0p21RBNX+g5ClIBsQc30iCBv8CzoB4nPDaquP/4XJAlsfsNm5td1TPQ8Q8r2pE0swPPzb1/F5
RwpARTRkemz6JkdQv6+fQk9PTQKdN+dEWgx1lVR0tcRpgEOb3BLW31OnU17xxZKwjwtwRv+nvx1E
klDG/kvaPGnDA1D3AuxeQDDZCEdIoi/9nAAzy7QGfODy3ILcyjbSp5WUH1oUdMsEryM3/LiP5o7Y
y1SwOyoAPw4WHdaOrSMSerab3grzjr3TFb8aWQ/C29n/MLW/ZnfaMbYuopTVtbxNviyaRlLgUvKH
bRlHPI1rhjKqe1NmWKgIDdLOGzlCyg5iDHUH8Rn5Jtu9ZNbiQae8Z76ffCt7ZGq+5xSPwxfpkM8I
g8KXlTCTK7/4LyhsXbo0s+2peiXlqGOPZJTlnt912fsUHgrRHSY2ExGwxXn8eWOEPirgnc0wtHUO
Mfzba5+x7w0dchYiZU2mHhDPr5qtE1BTwjhbOJ94yKuxxf+BTwoj7/3h4DO6aruSZeG3AkMtzC07
EUbPms8Y+JdVChk9P++3fcIPVjtMFYik72Y6RJ+yZUrUFiT1Oo6FhPv/PYHO5GAMYs41OA2nrpug
YFnAk+3/YEYYbuCnZJLIDhR9+GP1G/v5+TBXvuEYo5bWNr/Ev+do1Unlq4GVIWRItnfKYMxvBM38
krSi4nbA9KL9tGKEuZ8jcob3JxDGl2p9DJm5CNpzPGa5g6oTaw4gbdTyTQa+MyK8UAtNrLwjf35S
3MZIoD8g4A4o3wFnMkU6GfpBOztRffDRzoMcqtDaQK0rt0Y3sNIgbDvSQe4CzUuh1prKOhZhwxWv
soPp1bLyBjoFf1VA02gR3Zry1PtOc/rzvKaKQCXuqTK/Vmpzca8LW8HluXi9WeDynqk0uALCYhi0
EhzMGUUH4z7sjMI2D1CRnjfL/U//wzU66iehrjE8P1Ydkzba6HGZpWUrvWNPKxotk6jOJkhH2tQH
B+ZrVgI+qAMy2lX25MTBKNUnyuc/0dJ5j+eiNKsZnySO9k6WOyw0xyOZLx+AZflMAsTPfDo2OCoS
eSVlkr2o1D7kCm8RryWYJBuJh/AFnL8KtDokbFlJy60E5HEbjkD64EO6094SpPyMYmLzxwpy6kr2
YrXbqcK8D1D+3j+SnimXT5neSv1beqPzf3wITXZtJSgTZoYS+UKxYUsHy37v+46kkHOPljmWuWuX
CNY8MTmD1Nvrbj1e0Bxodl2SNLLvEXJUWdhzIKW41HXtmTuWS70dDv2Re2p4bDkkHL0vJwSSjgXj
rlTqBVA9XBR7p2ueoJwpWL7Md0YlMEb0hbUsItf9sfpeHTYjCPB0Wpz+IKx2VIusaVvl2AwJEez7
Xg3P71ZkFNBtNsrCSGnHqZmaiDik1h6gXDakeKeIohNkFLGOV3lF/RtwcVaLsYBtuweTSzvo+run
VxTD/9DlyN10QM6Q7GWumAIijCjroLinCH9QqdcuGrXjVRyQgtDJOkQM2JwbsrIOVtOCu5pw/H7B
tL7ZpZuLeIIELXVioNyePXkKaTxaNPCWJj73kad8PdtU3HFr2hEn1/fnddJMk7XaOzHDFPzcfVhU
+AQ9zryt1kOAkplCeC9VDa/vslwNCyopNNlraRUNBZNfH2RDHxCWe9iZqaAtd4vriP2cQbMuHB12
VSOtTKZCRy1rTquuir+G1I8LpY2AHJI8X0yWii9h/8/n0g8MGSFRCMF/iC0a4US3qcbqTFtLe/W5
pcyKLe2MK/hBtKIPPHW+QFe9hvbYPkNHokOGxh7HHkBVRmF83GZuGUvHBY1iRJyV4bfCqOWGMtAd
ZpeMB23koxnTwdGHORkzn0MO4ClyAEOmUBoAapOIMjBRJkTX2VzguptXstfuv6/6iaQckUp9kNKH
nHyP8IXNSRRz8jQqmKBGHoVm8xyCb9j0944r7GMvnm67+0a8Uev/m/8RseZ4yc55JsEQdXjKKT+4
iLxOer4xHbbepEUb0fQonB94SmC9mHwwEf8yvW6kX54bv+F+749dyXwvyJOZdQGKbAnD7aB0jEr4
7gnyqIIC6ejwZnLSXVhPvc0CJ1LEFsNzIsNb0WtaufI2Uz8Of0AyKSoEJpxFR85RIl/fuHKM3CD8
1Zg3FARoQUOWRWNC5zGQyTpH3Cz2+AbHQOI36wY3E1VXUXvfNgyW6dlRRQGnxtjiVcbbS0ECMGi3
GTUpVhjLLedmr0sZhthqYIpx59MF88MFzy5L0QCnavjKUPP6DHdxGJrRt5E0/nS61ClnfBEHiL/E
Uw974ixepmF2LITVfXuFDVTOflTdFeGvbYdRa+nobeQHga3oJj7YgPUjSNEqgxfO5bkeSaUA86NN
/vtxklnhBoZCGZiXWBXxOX26Ix+nt1Q7gim83sxonHGr6U1X0U4KU/EVnpperO9CmaPgKZEhk836
tS/LS+bqVL5LecLsj+dfvci4XB4K/a6qkEk29JlrsWfu3YPnMourrks0wKQ/dIaChQFZPC7bofgz
X6FeHb4PGf04tipsT7uNsuLhDXs2macdwkSs27PNCB5eqTR6SOryWfijMPOHGghQZXJcApQo9gkR
Xihsdqtutyc18qUkzP04GiV7wfoml/wzpvjUiYDOiWUeCKq6EzCuzo7qZpfCyqokSAb0qWBq4ymy
CQN4dpnG2zA/dMwW2N/z3xp56Tt1tuoTOoMsoidxFqFlv2RVGb/sb6LEsfniAgUHR2eOPxu4aujQ
Gor8kqHc9TUQbUajGGG03zVlJYDXlF8fxD317zGsRCgVZQCxAHx09tu3ksF7xFWKT1RTcdlE/rr2
eg/LLUU99PC2afmxth4D5iPHw4PbQ7AInidASpEk6kKMBKxyO6SHdHW70eUewYDFfD9bwtpmb6Ig
I3N/pIpPmCC6ji12VRDWSivhBK1wyEkJGV3JKVDnu6S3yr2mxJLf3WWb3wprOns0csl3EMJwPjNT
54KXRQfrMPyn9bfgQpEcX2MQ7Q+rmomSO/CWPy50AVGI4KrxUVkgJP/6lFpXWzC6+TxRLpdNHluK
WwhqdQQ4o+YyRBilAUyPURZm0aipQyy6vmG/Ci4Kl89tOR5v+zzEkQccUoAbRprd5g17lHCckCSr
qne9uvt19qqIiAgZ8do34ruIIE66Vi6IhxrelxNa6VCOxw1OWZWulpKNFM66zSwDxT2FYnO244jE
UfaRtwmMrbDg0bkpS2SiOCIMKoF4J3gYLy8n5JO1llzwmUr697XOQlreY8Bx2RioJ/X0P5eRP0V4
a664AyVgUghVqAWEqalSt9Ws0VKb9ehVSRWmSvQYmTiQWKt6X3Mamd5FgXqGGki113ZbAJYldE92
so4LYRbqtW6vBh1ncGQegVvNvH1Ds/n1+jBERaqXKzkqG6OwujCT1aBmFQur+X/dsfFDToHOp80j
PXfqehgPe++Wmd4ZvYjHVg9+LQPF1aJbIWvuyu5zu7wVsNttul4L9FvxUlBGfLriOctAUSCHcSOG
ziT5CTUcWCbiAddFqR94gyxUKjbDhxD23It+d1wlWDEYLLiho7UR3KUSz0evgSoyW5nOGkWjNh0v
yM0PJnfAAFPsciZDUO4F5nriIjFcVvIWHldtrnYEFKEfYakpnZVTnpQO3VBrzEpZ5hdEWJhXeCMq
dmOvRWmbKgoWC0Rd+5yUzLdmpHUxTlWZo+QiCE6hrE7go+ZvhDw1xFXNazP58fOPiNdimguXHgnO
nhv+ZAUzg46EcXRMT3GMgW4+Ne+FMW59/aAmE/o3IAVEgsPk4lS/OBeIdTGCdBZa3vikMK8jhbMS
mwSQaVgrtaL0N0MW5k45qABzs/9365Rv9JAHjqgQ5nPHWDJRXBdn7y9aGHEnbhs8A7PxlibrJ31Y
9D6go+lcujkf7g2rmmnWMczFSfxpi3hU7r8g0A1ZM2ErvkXlqmlOElkNWJNsgrzmMPBq7tvrGsCY
7yBqn+FgN0wmT38GK/pWalLWgwPYxVccUp9S38YDW+TQcgCzauLYA9V4e59t1I6K/H0nVCjsc9Rp
nFmtYHZaWqaHsdNWP6kPF++51gK83wqFsjgVcnuiL1ucO8htyCFN06qYg2FZ2GXAh8IHIrTtcesI
rq1LmS7QqiVd+GG8JxzyQVh5bDTxnD5/zouOthYQaQt5jsOwGs8grpJYO4A5v65lScBmoCy7w4sf
EGclAd+MjeaHtc3DrS8+61H3l0WGlDrY5gJrOMQ0LalhQjyfg0q0MFtsTV8Y436RsXCUuLfzxrn1
S5RRYQaHO3SMQ27pcRHjLn9sJQElV7bQvH21NeJuN6jqepwNtQn0Q4TldI6No7tvoYtqB0pCwqnJ
5m3kwzVPDxebwhM2ShmZwMzcyE5bgJN7lQ4kXUIEKF/GbksGx231sTqdW5Qp5jwsgr4edekqQ+mW
gAcqZyGCwzEA6YhVQjuTRQssTdpPVbx65Co7WXRIg51EjnmkfmjIalYolz2Oq0Sn/cdi2o25FdQC
Kynz+RVQr+n8CK6W10fFKybODAuzzH8lQpwGkRy6wYLEBYHoqbgYgUs/SFlWGo9q+JXN7EprHj5g
2fHGzllGPzlGDD38q1/3mpUrRC4jhKBvX8YF27dR6716njHQVo1tf5YY4qN1NSTIP7p7u3u5OUpp
bXchylXli98WtZ2lnpgffh/n2nV51LzO2pmf3+RsjF+zB+Mr+hwkNNTIacYCMHa7+0baSECvm2GO
xs3C/O6ubYYuKoXTozfLl5K6w6Dzb9hYq8/pn46ivt6RbqXVtiGQmwze/PNO2fzjthsKlrKE0Jc+
JdJIiX2zlHFrC0JtsMOZPDXtWvmFr1ynsgGx11Rt9YGW5EDUuY3Bw7vGPSBJ3lzI4AIU9vmLeZbM
oxH9h7cEbTlY4BFnUshBcCt4f2UvcDVzv5VYclAG1NxyEgZVt3udti22DahVEKDwqKGfW5bPxkp3
HmMX6ay1zzB02n9WRLbxhQBlnJ1TQo/lAlbzSLrCq1UMFSLdyPw/a6Tc1/bUoR/m6YcPJsurZ0lD
27PngbkZ2s/7p4IJfeEDMWlgYCta2MMcEAUhX7QnJoVLbRfnpDB39VdT9EgAWYcGKVfapjTJbDHf
p6vxQwYRJnUvN4lpzfKH9fJXZ6B8ZO00XuFjtCJ626BrNTcifAAdbGbTf0nlqQGbffTQSQ9lSGaO
wmLc8LN1agB+H9bpwtyLEIJlkfCwKyWgXlUrOAvG6nCokuyBBSOept3qBTD9z3hZz0FiY1iXofv+
Dztf+PUnQbn+fbyhiJrN8DPh8Wz+2lEfPHxYm/3ocRkdUE84kSvESXlSdWVXUeDCQ/FTlSNB+qSm
aZrhn2wEULPuHlMjKwpFfot5k8W0EPvVJGXaQXmU52xjC8KTW3UfYJltbV5gaxWk78jPap0xdxM+
XHXdcgylGBhqSb5pEVYuI/sCNPI35Rfe18ueBQQ/FVVyyBA2Lm9S2Y6Zq1s9NmXdgGR8XbCRYqqP
Pf3/N2Ty4OG5zYU5513FqjBPAt/Cncw54LpkxiXIVfDe02byfc70cEfn+0t1UCx3OxsZU/Lq31kt
tYv+ye1hlkaNALdYIv1a/mBE9wcIlFUItdgtFT9DjtRXkjLEXBTGgPhMOjy5om5Jl9ZH/uuZ8iUN
/1S4gvPdu6awyp9VEqgaXlnMaUy2LEtSFiFZv8hYb0tHaj404B/YjG0mqcZlkrSwQfhyrd1h082m
TJU9J44PDlRtq2+B3oRIlqaXuOfBYm759fR2EE1nK0FGDwwCOqixTh5iI+hjCh0pvYeJN5DiWsRu
gkKwki5TG2a1WFXjkZ0v2OiX1w6gcfxxwwreAWj1dBuFy3V0JhEgKzC6sZ2I1wb3i9yZ4QhxoRj0
Dkxlz/ZjuAsDGLAw1zeYaCu61EZm5ZUjcPshFbg015rB3767PpQYO/sF95ZapBr/HmJQ3AObRd+7
D3sv3p50NA/ezDubwziuEsHdW9ENCLPXvps2kLrACWJHGNUlENRFs1jGsgyHAyybuD5yavQG0UTK
IYME5awr+BZkgZpzIkcEDVVwz9qPo95hI2sqV4dr9dg9qIcAgTZy8h826VPjJ6/NvQiXTyPTQ/e8
CZyVVLBSUMFPOADH4g9LTaNkdiyhubihyM1a5G5zt2DKgzw7U3nrsV5HDKiDFRV+KQCS1hwJT8KR
C0uPGjGIuqiLT8dAjr7BTAUXjfujFaArhT3moCOd4heVlLyU7aI2fcgmzYlxZI+sB2bZpXcpdYZF
wnjJe8EyeUvXtVyBuYZB19ujb+YsJlTAiA+f3WfE+U2YAvO3uiuSOcTHLCGlR2Th0w5RNCZv05RW
9toiRgZcezjo64K0tp5EDFTSvUAvZZ9gfawAxzcfsZgU3um15Rjd8EOj/RjsZoq4RphkGT6gFyFg
aKydQsEJT5ksnb1syubpt3QvbMegXKt5kfY3dDs2495ULOUcxlf/8LQybCGNXy2KuutGqifUfBx5
w+xet5sMA85om68dkc1/LePqQJMYYSTPvGFiuttJlPtq6PjKummQIx4PaoEThkjwjZxTdu+BGRdS
nXEAfU+FRsdY4noio7OoY68Y2GtZD7wanxPPWgBgL9ygEZWgBacZVpBnkLDBOBnEqWvNWIwdHX2F
zOI9lkmbZRJIvdDSr/UoTsB6+8ErgZrLUNRgV03lHJoVNwBu5t5ddxpb/5o8m6jfBi6gObhPMIEa
17KfeylO8YC7rej6ZTvPBYhLILQf8HnB2oVrUSGzLPdFx+NtUjFw7Uz3h/O/jYyBe2QLFOMKnrgA
s6lXhTRzGR7k1eWd5AS6dm529UQYW/4OaA73omevAxpeeuXpH6HqBhEzEaoCuE6DKibLOokrb2i8
s704eukyPB0PCa3QrrhGQ//3oErAeb27+h+CPEog9Ju7JG56MtFKWs6pthOnSRV6la752Dz1CSJ4
2xoX2tv0jIP4lRY4eAnuLzpeCLQ6s0eQAIbq28e1AucKx9Icrr/Xb+KGuCrF0WHdCLx6enMKN3De
pxP2TpBPGKqVf34ev0jlihTJvPy6eHQFBdHrS9nmJtU6ce6QrwL56f947uRXF0CMjIPh4hsy1ifM
b4wPqj7d79WXH+NVr5GjfLdqg6jXD5v+2495PLDb6Yq+x+ZO+ViBK9icEgJ6IvO3Sh6qe8cr/GOx
7D2/6vOnL98zRBuX2iJw7NAtmYprJhnacome0/8/VKmjGDwZOuqaBPboWp/RqNtYaaMizdoe3kii
mRI/d8UaxJBwJUUr5QC0tZYozLhhJiyWa4GPfHkviafIe/Pq4WVpoXDL8eOe5tSuIyai7GclxZZQ
eE6WjUtnI2BtRxcmz059uLj0MKQbL9MgQAIWk1UXbl++uhqV8hAEtXyMzomKP5iY9ADLg8oRlfM/
FxMhhN+adukmd8mmxHOrLv0A5Fg5AQ4j6VTEXG5qyEjLzcQ8dSXBX4n21y8Wud34cLQM5UAJgSVE
KH253YdXSotsz0o/mSqV1TpbDN5/qwvUpgKqS/ajcnAaMCENNFQl2yMoOQpg+8j0S1fC2MpWSsZ1
GL6DFYDGvOj6tmTJk3HlQXKEeMqk7GodTcZTgAf1QqDu7zXTejASJlgZ+f5iKVyx4ylWOMRfR0m7
HmizaXKHxdUQbLLVGWf50CcsUQp6sAGSY6oh0m6Eu61NTbPLHPi6dsHlD/paWuB0UXohKm73Wyk1
HazxvM+cUNh/5eAbcVK1kTteAi+4f/aYHQGGXpz6td7L5NbL4nC0vdGcxjO02iXBQ6RhfpLs159w
vhcddDc5wv+16z+gX7crmZydMkf8qfREq+EFhQAzbstGQCfBQYv9iWBYSikOKE9f+IG62tOkL9b4
hjG82OLQmXUSYUGsJtzbgykHL/0iSfKm0bx6pW5XjiuCRuwSgDxHA4qZ3oMc4VNKVm7On3qUiqRF
S3rykjMC8/T4wXgmBedkkhquZKp/PyN6nTjh47Mq4eLiu8uOcqorg7QKRHus6GZ1VZHAt6TNerib
+Ds5r/K3GO9LVq/41M7eZfG9REJhG7JDm5j+EMVT+obS7dWWNnEZ3OehiVwx0tUPQq0a17Me+rzE
U1zi9orKHLr10yALOqyQoEbJSgHbRaYj5MRjZRg9ha7VOOakCusbn0BmkGGH3SoTxw59ANtO12V4
cSspo2H/rbKDW4faTrS10vp1RuAJJ00g7okziP4Bpeu7v91GwHOg1au1gdfmyXR1+0KzpqADYgax
N5Qq2qZsznguJjwokS8GHfOZ0KTQw4hMbHnCUZfJeh8DXXcekLEMFWbJpazuDl9Q9gKIyTRL9fp/
oR15/RrmlTdcUcH1Nd8EZbKHJZ4nuFZeg43OfT2kiID23gHICbl84ITtNiw2FsFw+pawjJA3SDV/
9gGzKhyVl2SydPgaXF04cN+Ei4QNM27T712jyAJcBr4Jy5Ht64XfbmXoLcpW3WddU3ug51KjB1tF
BFF256ULlb6oC0ke6B95d+QDGIYwH76pnIdfxPfIk817d5sg1jT3/0dBW8waO79fjrziRU8ANz2L
ZAE+zzjyGWredpbkMfRqdl0LsEfgOl1gKzAgV2nuSB+kXmT5gdPqYrkxLi9sq1qlaS3/233aPUZ9
VjzVDcyoTkq8ofpk3qsDx380I660IJza6AZABBE/08bbiQi+cSCWvf1e0bOhhQ4nL5d4M1vTIUDV
nlIdmrtYzGy6z2E3ly4RJydL/7R3CL7yLX4izjxjVHB7Kmc8cHyO5G+QGTzq4UGIv8fbInyx9Ccw
7CttB4HdpfqhMoKrUUS1r0m3ytZYDbhe4FtVbxF6iKFGcEiAbc0UjLgxj4M9Fw76RDIJIJ0AdK2b
bIutst6qBC4AXR0eMpck8BWUGAJPibt2/1kD52rVvZNLuC1IvHc2ukbxgUxinzLZy9pUTS5+jlo2
JjZ04TjoNMLTUHjpna/P0vh89dBiNKTmVmMenTL6eH56ULpg6kPPFwdtERU+/N9zY5MigtG4Bf2p
lxmiUdNhljeaavprU9Tywbtt3WWv+o4j06rnNkK8+Na4S9+XWLk2iPUtbZ0odz/kqxtZNCvKAJg3
hVrj6Vpcoc0EylixtBUkow0r55GoLUbUbUjCZ/MIWxF3VBsZwPz7rkv1qFaTnsTCrJO0/Of6Ouu0
evNysM/B8Q1RBAJ8nJV3tezl4by5ljHKT9UlFs4am1df2ciJ6uOTOuNhnNP2lwXLGpPUb0fXYGkw
HCFsMpD6xpg+8NNWNpo8lEHUyy2iSSgMk2zF92nPnojZrAqdF0IuWBKZCDWzorKuDQyMWJ1+6Tyu
xW+0E4Ks5Zir3je9XGYgF3WLU8MTrU2gcOj5oQDxGbvvdO7nKBhG5TrmBOBDhgEFKCmelIoYR7Im
GurRU50Jju4mJLKXXkMk+ziISPi+wKjYEOnNoGNWiQkdrxMFTIQqgBdk5RsuXSm+1gcFkDroSlVm
6xz308MjAjG/2m/VQ/RtDlmzA6iFBKv40IdwhjgvxG7CdsdIh6xeINRzT9C1fHzTUDoBRFe/mE9h
Vb452aL7fPUQod/Y/rtYVfA1jMtUMz5ii+ASrL+e1Kj/Ze9EDoxdEF03jSL1CPzJV9et4J1OAVVp
tWlbXmaQ/5iIHBauSswM5uuPs9yBX7WE4dwb2pIBCPtCzynbbBvgspLhsDeP2Th4RizO6+1pBjGo
mzgtgnXPjAR791ZJNXuh4opdaMBnPpDL9pzid4UmO3dLYrXHeQkLe0anpjfkkEx8w59ul5JZ7KUL
vcD5EXf+ki1DIcm9tlqLBWE22twP7LPeJfI80XQl1T3gbe/Z51jFZ/hwNUwedNm3R+yI4xZS+Nhg
X7hvfdhJ9+Oz1ZzkaOLaA/1iOYjC9D9h1i2pANVgpn64alENIYM2JDfPTcYWxCM8vNb8tGkd1UD/
n/PgN0ncOnRrCM7QtpDqK0AD4mdPkbfQvSVtrrE8JLHjMNEpOJX6nevwYtD/tdImN/ztdzmFeRPs
KK7A7siMhehgpgq/dfkDypmJ4lkiFWecDJDymoFWafj+m1MX2nlUsEFPUTYc5g9RHI4Q7lOGlEdZ
2DCfmfeB7NH2tHKtTsanwJ3R9kU+eXQTVyiTUMMxlLm/2SCGltOeFbFi92TocXtmv8I7tPI26vI3
lvY3f7hG2tG3tpJiuSp3s2MS0OR7DSKsRgxrGYB4uk4ZKSX5houZmRrRjZrY/2BXRoTNz8U0WKDL
XlKc56Dhu3c+X3eoocVZWhRH4ss0dNmaAn3VzVS5b6aS4VHSJgIhMVLD2ikgHkZLvNVKjmyQO16n
brUC3XK1UiefJuVic6lo3K0M8nGCFDbWsqdW2J8g8EGXwXJas5X4ykWSBEqiITLZlTO73ejx7AI0
px8bRWfs+j9BK+Lz4mYQAzmQ+/IUr4w5zEeSWzwMKFYRCHEg99bn2d1Cm7Fc4h1gzE9pbIADJZqG
bcEYrO7zZVAIaX8UbjFx1KwpbZldfz68b4FcS2iVkXV/UQy9v/Gr7tjM8N4/SJSUOUxe35yza2XA
n6VfacGzeifhnLqrvTqlrZGBt6y2fvsLwTyTTSolw7NBzzeuZVtsRz9faFU79DeRhjNWIPVBnxNI
/zjehpxRaIlA72v/2wgKhhFHZQsELFFmiw3Iw4vNFlA3g3IITs8ZX3x/HGjU3noJIfZspOxpdDgn
pdlFS5jsfxvg10dUZFGYVIPgz0iT/a2QJe1inlR/pW/lQ8fUKAgu1kytjqGmKXrDm7G73cKVAhEj
4HNH+sEBKFRRbmHqM+RMuj1dWF/bu2aP64IltQ76RB+WJRzygP5I12gVU3g/XWd2zJ0QHxifaHBT
Zk2DTNr5pw1vT+TKOR5aDS5nDVOqCjx3FMEV7exCnck78QR+Wc0JRXq/exo53akVJaGCnKHGYr6f
BrSB33NXrzE1pfHVadTjphPy21DsFgHzUsNTNwm8wJtODgqECplYxkagiFSfN8GZit8zIDEJEZo7
HsZw32j8Mjc49aGTvHRQYY7OgUHvgaQdH5OArRy1VHtTMIuTDa3uEKPmP/3dhqYSgJdABh2P+MpM
4dfEbHvU+W7EbJQGz7Hj6Dd+gSKwkJ64J6iIyAMbZ/XBBKMHbin1wKeTn5MhW/vII6POO6HuD0TV
jisKEb0CCsbe5Gqy+6jYWfIwc4bUYja4Zjzpl8woH3nWweoGYme3HHXUdAkS/ZNqrJRhqxm8vasX
AdBOh9T1XzrwE55Ftg8vyexfpEJFDsRPnVF/ur0J/YMYDdEHC0VWEOo38nfT9s0QluT1/vVV0NlK
ikPBurJeWje/0J42VKhgIKhrWneZwxbUmCUBv7uUVlNypDM9xnmL4069lM+HeM2N+AIjvfCEtVWt
Jqn8OlgrC/pDuAfbOuxKvIeAicyPrlJ3izvmtq3hjLndxwhDNzI5mxiQCy6RhUJv4oWLpLySJk9s
Td57WLIbLnj7Sk5aL4nvZn7ABJsRcEvAUG0qZ4kfE/aomW5rZEiv6Lnyk6lTJ6gr/Tb+ptN2kHsi
FBZRa5FogyJ1BXTaDPVQyrN+raRaBNwmrHdDACJHS4GlVrnldpBdXEHG5ThaFMBV28fPovTTXIx6
QKw/cMcLw3f+3Izr97TGVKDEEHjtjeRFq6IeTP2WETbN7PJ88tUsaKcjR7i2M3k6fZDa2DIbNgrv
3m6i1VYr+wfNtrL9s4UFGcE66c+HyHt0lxrchIqfT37DqIYMS7z4DOJ5xkJhgoa24yfMHkssRYrs
bGIXlqfIcu28w96U/4Q+hfc1IG9sDJDzCDxxI+kBLiwwjWSV+fVMqHFO2gc/DrLKJaHdt6y72mRV
4IY2246Sxarhtu4/ZlmF+xbzIM9iY/YWpMMBgMOkD7s8lQPY9WYstQL8ERTradECOxHNcEzo3+9a
zItZMQYp+VQAQaD8gWpECn+uBqahVDldRPCGMabP9gd/ifXl/PkrI05LuocmvLFHc/gcYJ+/6iqM
DXy6mq82Q5IpM3jak1QQ4WF6e6DuxywZRg3ER3p1+xDsvddXb1la9uVVB4dTY4JVCV+PYGeX079D
PlezjFv75W5uyNVqHk0Oenmc4IWs9hqgzsZCKDyf+qgHI/Q63vSy0qFmGEiC6gFuqTOsAWVaoZfg
ds2yrnMKpVZyxmJy+N9upQiieYtmWxNq2xZ07hUn+EnXgVCQpqHQRPpNH0xWHCbRvPQN7nfdLFId
5JT8+ly1E60xhpeENeT1TFg2f6ipygoVwwib5o+uoJ5GnXh/mOoSZjsQBTRi5azhn8FBAf6/b3bk
HmalXSdwLhrsgk4NwN2zot/zRLJCM/M6Jdbd37bHA+sINO0xvTAIRu9rrGi/jGI+GFxQqEorrhbr
BwKXw5OUzYlyLwbZQvplqMxUffgvWErVz2PXwPVA6bUneQRma3O1T4zmKbdYnFbb5R7v16qcb5E3
vPiFdYmOAshM8Cn2QQ4e9/gnchaj1nbIhbHTEHSBNabj7G0uBh2KxsGvVDnReoCk2l7Gn8CqAbDH
pSBZTaLoUyvHZCoBI82/lKGkSLAptrgH1PMKoQI9pKbsKDq+1dwib7i5zF+H8U2F6/Bk0zKj4V38
/zSANpJKvNoUKHHmp0DQt7o55aUVGTwxPqA4DI/xi4DfK45X2XeKbSzd/jQXLv7TrlzrehWy2p/E
M3Ms4jAFSfEcv2ZNbXb3ng5YWMBeqQkzozKYIxZmznPZ3TH7IwNjSLCyH+reLvnhA9tzax+93yih
qaD1TyVVCMnoeNYezqdDAgPMk0F+FAItcOa6dQA1F/fC4QZ51J3eRM0SmultFBwK5nzOc2K7eXHw
cIm+cIbus2R8uxEvPVSWb42NGGSgTc+utPzzaT4QrjsqEi4A+QFGCdOzxq2ZiR94hZBwLwrx2KnH
WYQERz1nJYrqHyLD+8P8cd6U3aXu2UyZTZ1yfuOlkbwn0vY9rZ/Oxp31iXPzHZp5ymosc1Pph/3U
RNzFdlVsxH7ehSafL40oV83B+dUexRxZAk7TWfR3IypAsoQRLyiWQVucR2c95u7SqPA42XdW9fq8
DkzghAhLAi/+Nh62GQcocEJg+bhwJbfD6Uxx8YBgDxiwG0hq4Dl0nzx8If6z3+nEd+kv0lnnXZbq
9hmUAC+Z8yze9zlDHah7TlPmTEfx2kaB1s4df8/mMtdsoIH2GyUrzU18cqWq2cfBBMr+bc+s3fjU
0L6B+HsPLgLg6naKC3w3+kGjOXb6j9fbkK8N3bKIfuC1PgEEbxiqMEBRIxDFtlEaInNOLtNCJ95c
s5gPv6s7Vc+f2vEvwQkK7aU5K/oDoKOA1p+IB/BbeRsKloOJu0Z8sEDyFWOpQ4DFyzGYtipjKKIr
aeGZ/5cDHFDOcjRO5K1YN/OyI+aVDoLWN1Nxrrncgrx8Ur7Vj8rIkw+XdH6ugwhvyj77UYrAu0Il
7DjiuBaQSzoe1H8VaVP6ykhMpLoiSiYLgVNo9e3kyOAy8Sw3vvt/Gn3HC2oOt9Atkojzul724C6+
7owmJ1NPJ1Ix2GpmEgOvpH7WphbN8P2lCOyf/XqDmKSWgpHvrCMGGrIJimYU3tI4rBOfRI9I5fJk
A1Yfq+J0akgIlH0R0uTc8yFsLE5Fyj/JTXiSWJLDMLIzxBiszA64B7WjGnOgThClaBsdIcC5913o
4sqf6Po8f4I0TmIiXsl1leJF5CVNcNWBeSsK+yocZjozGBg2rEy5kp3NrQB5fnkUHoVqE/Tklm+O
L5Axlj1Z/c/Uiy2/iSYV7sZHygwNz4tDVp88fhWlYnN8nypuu0afv6xCQY/HEq5yly1CcYssODWc
fEqx2M0U7/hxt4D5LSIM8F2HbZpoZUMtkG4e7ukNuC7SgInnE9DYYOJtRR9KBfO+zmhw3Yx2TqxK
8nYLLi4ZQYuRuuAw7zJTo8nV2qY3wGYdlPm/IPw2MXArQdHtnB4Fg+zG3TklDOwJSype8hU9XeRe
o3dMWQtugfAcOpbBX7RQL+Bw8xk/c+b+O0g2KPHHUkNYsAolxYkh951X02MqwJ6zoVelx5QiseC8
xGHYxenEvoo10j5v0t5G43gBbx9Agkl0Q6X20/LlB2MnqBjjwRAGarYF6sWLY5qcFTNf+NPqBuVd
VVHZaWQrBPF0zCGhcuJ1YV6FDN56RyfL1XLHDYj6DaR+0TaHBtJe9MU5gVfDHwZF9idD68DMpV6t
aYW+RbzS/MG269rk5s0OU4eaNUt1DaBcgjLUszRsKIVsINx/eFtxgWIzC4DGj9FY5iF24FfLG1EZ
0MQYdbBHayfo34HUSjbIRdG54kmn1uAfcotrMWlbbQAK6X3pmABwoXfmWTx/+vkkcK64GE5fzzuf
G2/edMknJlMR/V+WLcZhk+cS6f2APJexU4aa20uNsQ95orwyNGFfSWWL2wLKLZsMXJOWNmv6m/ct
LRL41EICto+NiH2fgZX1YsB+l9hxGecVmu259rYV9fN5qqghPZ9vNe7GRJrhcwejmP9KJs/CbbNO
VTJ+yZZpyb3sDyl1djNUQTcnvcn6rR6zQRnKowWRNwKnZFOY6+V3GuKwYK5KI1FkYqE+ZgIgSQob
XuPnVv6D9/BvZoLVdDL6gitT4rymb7sxSoAhPlZBo9eG+CxVhpcusH6xQUE4/uuEf/eUz2T3xr5g
fyyFSqxz56fqs0fCLwm4YPkgvDmTTdBRSN7TIIJu4R79/gnyEYxDZcEefbOomr/kMjCUReyYQhc9
uVU832GVv6pzJHrArSI+c5btbpkTvm3S3YLysoQlqQ8vJlcXztPLusl87XfGKbraSbNLS2ipo5y2
ptiL8NN9ntX3wTheqhxnPV3kGKVVrldM4i8tVDwdNo/mWTooni0YOFHICFl/htigBYeSgNpL3Zki
T8NxYtJmDFs/aTLYF9uRJX2AdvM7YnM6BsLXaffBWlaftsTggR85KXwSHAzPhgrsewr4CvbLWFoR
i8/EUx6OkzUCxZwWOmpDK/ULN17Nsubcmz8aBudkyjSvxntGomHxUKOiOPMAWUkYcjlS8RMMjuko
OF0JvQuG1l7MK8f+z8Gfd20PPwoCZzxMKNWokibUkJTyz7fH1pqqaZubsBwsaghmQdJgC5YpXNc3
D04bqnAmHBiiwGRo9Mpl+OIJDBQAhY7qlRhIwfHez0/bJ6OwMP+soCGhMjUmD+Eysm2lSaVv50z6
6aG7Edhc23BNbuw86/U2mW8IFhs5UHmSAX8+G8QmGqtr/cA7fShVWI/CcSByVJM8ZhpUtlrZugNp
m4rndsFk3kmncEnEHUnb1PWB8cFAYL4yetVtK/nx707FXz2eBQR4ukQrKHQjIId73W4t5zYPd+Y8
GF/aD1eh22raF9H2mhhUts78C/DCXTsd3D2JzQEkg2QZYkZ6SuQwJTN3w7NvEulKcm0zfdHSU64v
1wWpaNwh9djjyogViJOpnLAPjRNrmhNCuqPGp2kLm0ZMel0bYZVygs/PHLkioNa91V4BXAgjJkSF
qMyFgZPEMNfvvH0I3+JVZoTiRG2xIw7TSlO+Z/g+vT9P6MopscORwgogCuV/AgmK2WNSXxrY+smU
WXlvwYlCyKzCsUZsI9HAyRnypL4KCrLqDnCMM2TSyR8B0ehr/mJr5m6cXVDCDZrINkXGDHIfT3kW
4pBVgPKmY6ELZZkvmGWOp6bFCm5rwECwYSxnSJDYP4aG3cGRAk/uCutHGv/tRJLGw8wdrfZ9QWPk
QsAQU1SMLzQQ6ip70D13eemMzsUfYI4eBEW2PeyJFMqmfXu63UfEIWnQZi/YqvCvrYyoRVRmpq4J
nDzOHDqw+kx0hftdDv6mUkHGs0JA6IqJ/Ab8T7xjJ/Wo5U8snxIvuBneKQYri/ISrGWVMqMJC5hY
d8UOeQebP73MjCl8+RY/PLpsvIoDDMNf14t2VckL0ScQIK6JXdBChnVQm97GbsjrxatTcrru1EST
9aW87NcZE/yfFhGcTZifn5iX/8Is2MYl3xZ/jjurVT44q5kuLIWcH/EBifVYndz0rvlkPkVX45Gu
AuE/g9eviI8xbjvRrAi/59WgDbyyXv8qnVEwq3RFxUKeKTYYa5L23exj0s3tr8Uwsnooz6Rmsg/9
oI0Lg8rNJgQfwH9Fzzk2IWZpf1qCyQDmBm2yolZbcZtv1FodrWTSSKwFQQwChZZeD+TLJLl3V7Jv
frBMJUFSpoi0t/qILuUWAO3wD3QGSr+yZ6MH8FJ+53Pjy8q36/29MRpgSSRIpx/T858mb2ni8Mzm
iUjcKd0pNRDV7ZXlnqbx9GRbNNQA//GDJSIbFBG2gSx0BH6Y7szYaL/YTKNqFxRap4UGPFqh/7uE
iUbwkOOEN5BWPBuR+sO8gqaknE6s4orLomlntVbMdS05y1k0lRy39cuJlN8KtUQab056UEvgWLK0
SqMLy4L/i2mMy/PXrnwoqQJ5MToRJS9+x4cOjmymmQ2IGmHYl4+56wJ7BOZR9X2T1uFcu5dsKOLi
FrZ1l2LUA4GHv0WMABTz+gfNbAFukKKu8hzATU6ZOviN7fAPzHzS4U0jlktcYPieyD1srixALM3P
e41djovk4d9jxYKyDKloqRqUXaHlLyEFUMlihq+Ti1SWwgc3xtTd0/aKb2KzZ5ZPCpm9DM22TsqK
evkTN1fuqTi3mgdbLE9S3aMDAJoNB3QR11doq3FcbNWYFvlqIVT3YCuel/PUHhgekmjQofwp95i+
NgVliGfNH16CiRkZHLF8XP15uuZEdzUf7KwJUl2aDnrqbNtQoiLLrEuDBXst90ujL7Bzezwp38BR
PlQMWmgX9ewbeOx3fpom0zcJAuwNODHyoT7Sv6rrLMQSm0krmlBpHp2Y24m5YGDhJVaXqHrIq2CP
eVvN8o4cBYp8l5hjcncvn5WYUzc1Qlt7OkExzGdY/dM5MJfnHHUnM5RKoItlAJwskuwTVjO3baMv
XNrFQd0UdMRYmNHwOKvp0C+EcqRhtY5TnL3sNkQk0NMI/AFR85+v9Lp4Uxa6vbeoiz7TiHDkGbDR
gn9vVWlHXmxul/aGr7J41RraCUDiVVFJl3EuMzcasim0gM8KXDIoBLMd1bTeUJ9194sHQPyKpdtk
SvM3Ie3a4h5sg31D/JKXgIeHsM15dEX5qNQ+xOUvwJ2euzVUXrL7GBbaszP8T0K0FhKYSHHmrs1T
5xfJioCoUTrAS+BGXeUizYKGgKgg9tMXThp5s+/bjoiBwnd3SpVXCezg4enNYjSgcY/n336941C/
K+LztGEiL6UFu+kV5UbkANLty+X5oqt616wp9PATpvKVezubDtjl8r6JbCAIw4j9hzRVml90hJcC
R20Z9UI+WK5aj18zC/YsJXcoySF8EM17jOtcBQrHVkFM8HdF8q+wUQ9ZICe2Ba2aGIVytbmW75Mk
OxpAIGLfKMZE/ikYCnHT/fpryGHdpcpWkCWDuh957hhWoYeofwF7n1SAefZjUBSuDxj44Z+ypucN
VXCVLslO1Z1BKItyfNB1+rYw+qVCn2VEt6CGOCMIATgCRAphBAogDSo2+w0Vb7WUKjEt5aH/cdb9
c0EakLk4BHr2aSVrt+jNew4qM3sL+A9MU5lqzrynSmdxsusUqw+Al4CIddyRa/4LkW0om31mK/f7
EQf+YTagkdTYBCW5w9QDCkfW0UmB/teaFmmZ2VYqcid5/G89ifC5To5UTFIyoMWuHCazEoiyx4cs
6Ms6U5bL40NgAk8nMdHr/ZVXHE3f0zct9wUNAZ0eL8OpLsy4CS5mZw0DR1rW91XqWqyqJJLUwg8M
KqyLnUaxnl+F5WolNslhtVpnbvOUDFvJqaI/Bv1B+F0SDEkaYlwEr0eqCEUE3zsDPlCkyN6L8xlo
vvS4VfXY6eXqdgRzj6Il/WY9wo3D5+0W7/mMh7+6NFBUFd/TdpWd91z0OSTEaAcQ2DdRP5JMlkFJ
f6goFMl7Jr1BhHcUqf8UfhP9h+p8pUGNdVvYhXKM5k+W9eAPFYep+FJaLWgn4qzWfaR4po5bdT+/
WIAxSX9eFfAExsZrgyfxrBELAvNorslD25U2A9yhtFT72LwEG4Rf+6pZGynJ9D1y9Iv5ybQ8fVvG
RTa8vsSpzOGkGh5dsyjAAJXtsEpDmbyhMYbM86ozstyp1Qdw9xhp/aC8iLQVFWI3vakBTHzByb7B
m31FaQkxsNYKDx7GqBpS/9E/EgIRYBX53ork/9C+FaMT70iuYRMjV89YmZwjGrS/AXDxgVMlT9rH
ZENf1NTpdHQ1HkJ+LFvdXmrHWfBmnOWCrmHyaX9zpA33xKoPaWngJFVC+6xLw2hpsw+ucLackNdL
wOEg4NY/5ebr7ozFi5u0grWDuItbfNeu5clxGUTzMy6nIhPk5oFBZoxbgzp6DnNKf+XrL+M7xfAE
/r08yE8yQvOfwO1OCTA1zwUgLk9nQ2iDxVVauPKqFlO2JZmsSlF0p0JxjGhp6hvhrr+n20oygc7a
heCvp9sCjuaOuDM7hX1RUd0l0CyMOUDNWqUMeXJhKFzzoo9sNH5CP7Avzvi8UgXXlx/0R1CnROsi
kxPU7MhU6hbGoSV+63CPLFfvArgbyeXw2kfVyEAnnsRV92HisTM1Vcg9XUUmSn2qTOnTfrmU1MvP
d4FWqZtDkchAyNxlP/x5+Xv1VcgbHciuZ1CBdUpXSJgA2X6BmofNi6tVSIi386oV8SBYv3ekok+Q
U2tAKEketgB9tV6pa34PePvyFj/a3m4+/KNbA/98YfWycfgqHuOffKIoxyeJmwJMOT7xFV1AkfRQ
u8MksesWMiQBa4VWWuSfHMsnCFKN/FDg5qc2Cr8TRYzpIVpqz/ol6+BJn68uDowJ17v326Lq65Wc
W0nmjGbgiQyJw7nRgcqpVWhylenVZ9gVe7hxMt7DxUdkUdKPLt6URamvxccN2uoabtlSVEU3bUSq
CysS04XjApRtID14Czp3w8SOFVen0B+/Yh/GRPcBYDnNPjSLkX1CkdDw3pHJMmCFdBdLiiwV0mSj
M/sNVklkQCFzRfpCNlTLpxhRAw7URJW6t8XMjAQVBoiran0eriRoKMOF0idh/x5ufMxzyxwTzkdx
y70mPAJDFYL7vJGkE4DP1wmgExaYrTuVY8bR2VBUCBYGUI0TORGPE0nXtbt6eDQsA+X1S3IR7y3k
EAJVkM8ZiaqZJ7q6UEdT63C2Iw/m3vjx5BB+rcZ+B09Zr/EWb9YWI8HT5oIfI5VZHWqfab4sCMTr
1SJVrWAQWVr3W3OCWreuuUsj7rCmcOqNxjH97E/XPucjZUPPxwhcDDcJBHhpi+AR75Z7PtrD7gWp
MqeFk5JAZaEWUCXs6hDuKTJGa0OH8IvqMA75iw8MYt1EtSHMOPRZDWnpmlTGnd2BCPgwpu9xCO1W
zzXaCy7CmSwKimMFEtOwul5F2Wk13FdmWy7j5x/rfWBbOdOrZSmM1EsgS0rYwKLc/+UiesoHKJ/Y
YtuRVEeoivn8WHlelSlvJq0xJiyif2dtMInA/zgsKuv1/piHRXMjtXCQGGInVdplXx159mhLdVzp
TRRi5A3DBIM1NbxXvoAGSQiI+m82LA6Xl39IHXONL/v++B3Yw+i9JzGBK4nRqiT1hMnW0LTpFwRG
xwvaht/VfYNSP/sN0nymV6qUBqVukTFXjIVHeZ5VIq0wIIC/KAGfWLEs4fysxm1omxaEy/+29VZv
XnBfTNZXX2gmPFjH4paZGKa82Jfkdpi78jkqPJ7cYn9vf14ptTlihNVr6aRdxaMQ/JK+hg/a2P7j
GTxlFa2M2PpiQZOxa6+poBO6IuAaELC2GXWISTdWe7sSH8sJJR3szDHB5I6DapMCP2i5Pyi0JGOS
avQ+JVL8vchiaJqhkmA2X3v3nNPuKKp3D1HzI2mngYID+h2m/1dGR9Y1hx7FXUQtywMnmz0OUpzj
27CJ8zncSiTNNVEYbGDtVzlHxtYV6gu7lmR6FdU5Vjy3/8kck6kt96PyShQKjm3w39ZHJfJm2kne
fP/mnrzMoqtfuIgIPEWNgr3f7Cyy8yGR9y151xUY8vQDaOlZhIuU/EeaXoiy87OBlyxobP24sY6n
Pvp4nVN/UZXXfoMIotYd9VJ+yd8B+ESd+05D/PmSFUxpEX4/exVuVWAJj/EX/A68YggW4rBUioNe
/ASPSq1SmTWznk67eAyH+W159RYcTJ8J8DbJQgaXlej4FUIA13O21TJjLr+lSZi3i+vePbipbiyw
+M9gjBtBy1gTF5sDjM1BU72HOt6d6G5AgYZpABTh8iW6OHRSRcQUpZTNfISmq6mgTA2xdFMBVoyo
iAo6fLfofu578j6TaXmqda1zV10P+22EG/QrusVe4yN1JTDlzeaxsAVSLRJi5fANdU1+GAHefOod
/XcFS64zeEo8BuR+F1iYBcbrrdBWehDgAf3wkywhjdd7TSM0AvU2aCcd4NHAmSjYqGyxVySbGt96
F/iFi6i7lc4pJ/TyIc7qupksBgfLpShIHp0ur+IsZjlsl0B+54DYITSk+Bciab9YfD7iBKc4dLM2
92PPcEikPyM5vAnheKsopKkAp4XsmeZRE/V1Zc80MRyCje/q4L+mYdzRM+sLaWjuomnG91eNY3PL
7sCmo1JpM/9uzH6QrnKU+XWcYs8/2mqm4wOXFx0n7b8vWlVfyU1fLdMvu1UiNCueBbsnK8LoceXX
NYkKnvvtOUiiCX2v2nTKO85DPYXpqO03M+MFl4dy6epmVcihCTrt/ESl3nnWvSWkjDePAodyfwJg
2qboWi9p/2T+MGVcZp2gDejyCHbc8XAnDhx1DKEEDuNS1c8+zskD26tJRNRypCmYqHph7oOQkWFz
MzgH0yi85ru1apA2sGpzbRyc7i5bZaaTdJPrpks79+yIthxOxY2P9rD516VY8vT9us1e7cHELN4q
7G64dt8e6yB0ZMQDqr6K3X4ZMWmLeq9uRCVJCcdSoOzPQL6S3CtawRK3JI2KIwZOUC2TSn4m+pyC
1WWeCBZ9GTHZkf+bSsnfOM9U5unVo92j+0oO7LT3kRS6CjziTjLhAqwyxXVTnfmJ3OGmcg9IMZhp
fhO/BG8p49NLSkhTD7cc5P7lDhF9wXSU5lhp64JgM7pEGsXeIC/5A3zhGK4MdS1r6NLB0RisSXeD
vRtgmnRLXV1XsyoNF4XIOLuB9n6E8sQtlMzrcs8YWjEltz51AG3BV4qlEyR68XKdgzgAhFk8c1AQ
1I6Cl9MooPpWy35VlI0O9Jsygj/V5cxpAHG8WYvhZuJnIerE2fcUV8EQgIewn+Y0gj/jEzaOW25M
mru4aW1RyXMd/W5zvvoAfcBFE9BZFr7e/1fsv9CHP+ZdKUaokfBqLdfYdTaDIHTnOMdkEsdMCOdh
gFcqq3SztJFdkDC7HIA50dBXbjMaklq9GTeVaqigdrMxSwmC1dmJ2/nkQeIU65tlZpl2j0l/n1K0
gjeDGUYwDR27qpxJxjK4IyeqvFWZ1NXMYLl0GZfJ0RkTCw0pLe1jF1p6r4di8EOiWuGH1Z0m2dcg
f25gXcAwI1WekFSkpLIjk0IJ7VXJFzc6ULFh3H7zcFRWTSoxn0aMjW/B1wl7R17357Q4/Ld1pEDD
1ynWJKP3skFq3giZDnjoi1hePUwBC3JFIu+VpLKfNZydkRwMpIYLirS5LSe+JJA9mxoUqTibLsF+
78ia8bEBCCIR+RbtagL7ONejh8DGjAiWHHusxivSiZNWlrMUEYYrnhnZS9Q0qSnvnC5EyFYF2YpG
uM4wAIyAAeSS5ix0lWRJ+tu3dTq/hVNHkbNjw4HBWSfDImaH/gXNIL9mJDABVJ/Kl1F+JOWZetQh
GZKlBaeVmBlyLRJ9C+Ef5r6xuzHAeF2v+HuQYW8kXYcIQefDe6nBhX2LieTAb2bWHlU9IyGTMiyr
KyKu/SYgNe0VezgcU1wWme9KdZDPyQzGwkzf92FbZdOB+jJzSKoLWEJohdYhTHDJrgZqONVnpkUs
VWoAULkEDUkezUJ27lWukoTgLu2h41LG2QiQ94mDMogaEMH1TJNmy6L+WDBGq2p+RUSUpk/MfoXl
NTdvW6Z8KyJ14Xt/JnrkBNSolnYjMTSlaFFmkROXYoCEFmhG0vv152l7y5740htusGzQ+o01Xsn1
akbDSAuFmGpyYniIfDT0TI5dCWWfn+x2nv4cTi5Y3s+w2Wsi5983Gwu8ixSQ3O4EZicoCypov/3r
41vjOt+XGt1ow7gYjo+ahjf+F8w2NaZpCESkDMWHG+bERv4VQwOsq4dv0GJR1u7+oh0QLqcBx8l5
GKzGdza+/4R4iiqPcED9yhkLBqNvvYx5oYwvqp2SGHE0SBRUXR1McZU6COLiE/FhLwo2AK17EYQU
CFLeuHOBvRwgvOFhPCUI8zILw8Skw2szqGxDCTMeEtdJUv6N8i0WXmrc4Jf+MKk0vhtKpfMszc61
z+mOmUwi0uBjDaXIRDez2gOaVgVZ8Zriy5pAmy1/eyUi2gjtnBs64tLHmE5GidaMxgT6o7N9zEcX
CE6UnDGSymg9fQ92DoSr0Kyo7TNZGjCqWDojR94LPQVmNAkAyZAwvYbT9pXiKVXLM6c2dXgNHiy2
n9eE4m78vAQJ93mzj/3KHGyFmSBwR8I96af0N3aPWtgWPkOuaeHd74cBY/fzovsqQG8HvrJTZQJD
6nHDr0yCk9Z0OfeRQHXLGMlUD5Qim7vn8ZfVaHC72obsAXs2ysJvCSz6qZPkKzRYhKVK2d7qeyVa
wmqt5VpnIojcQe0R1RnyDwzGMcIEOsWAiVmqnHVoKFWHRXa12UI8pmPF6P6rP+G6zAvam3ervJ4v
YK9Qmlh0WcF+TkaN9jN/tWNKs/o3Mk+4KW2nmo/NDPUCo/hkEAOBBOI0E3+DZsPuhmXyoTySgsV6
m/FW1stjgQlBryPyX4dkbKweITpYsJjj/kRnOjId+s/CfcaGgB2phg0dDvczBXmQ0jBJO20fYDeb
MVQTAoYxoqdROguJ9Z83Froza2nGmgHAb0C+6+cYw2pUwP642afsZQOVIO3jeGRwV2SEHNs6BHyi
Nfesd5dmGKTaic/LDyXqbvTQj1ar4UQnYYbAIMNf0DCfXNCruVofy+S9pIGKSb3cCgQ8wlSKXdft
UxaEHcuF3xtESrBMefGmhW27VgeDSqYoHql2biTI5yYkxBOVZU9aIGvqNEkOM9gMYwGE01rby7Hh
vknBSOILVAsa7c7Iqe9IoJFF1q2EQWg2iyBUoqFbEl4mReWjEOcJAVa0FvAc+29Wd480pyhxt1fF
ByZ2hIKLlq27b/+avnXisvy+GFHiej5TF5ibsWrb3YlDvhfDUZcPbiW1AA84e38jJ59oOSV/TNTk
Jq3JsiQgsXdR7UxehQig9wYHDznB4luhGsTumJex6h9k8MBGSBu5qVAD6I0vi4Tl8sA6HUiKiAeZ
GuTYaKlXjUDaP43MjOtzvj/WEDPIGnifikNgexF/T4AI+PT1aCkX+sRZepKkxQFKO533qW5zoXVa
1MvplZjYzot0Qh35OYmlAyAh5zVZf68saIjw07c8Q6egvNSFqVjgNIMhQ523pZm1VZuK35N5Lekw
oFaZvcKgos9Vw0ZElSc7gz+6AcXzbQumBIrd4szcT9ZWnOhLSg2wDYDxIbsCkQLEKmf+SH4JbLV3
VnxvKx0wH0v+pOQ6ygNV+so6wFMljuGYNH79WHmOmsw1+xT/GxxDCUKY/HNQwthjvYit1Z/Zqile
siDkgvpLfyAN2PvnXY5I7jY2wDyqZ08mM0p8n6EOIWUpG2vWk77TKQyoj2CWFo+sqXa4hkrQtmJt
/vaa2UC8INt/ML/RVdUUkYRXAWdYa/NTFwBEI49GrY3WVm80OIbJUtvH/29Yn+7zGtfoEoDHdMjl
n1U7LCbCm1eOhS2BK7pATO6lNRZ8RkOcEFXxFvs8LD642Ymjr5YzuzdT1SPEjSioa7UDTZnqqSvW
rt4FR/39rqmFY2YQWRYRMs4Lo5UmlPaDWnML9lFcNJQGlxVNiyBXOpog/glKQ8P9SwZ/sDR/5PtJ
9VYL/yPqAYa760yJDtOruhwSQHv8zQBJezE7EDTksgTTFTw5Oqw6B68Tsuq8g1cxcefVE+BY1Can
CP2qLuNGKP1VD4ndZaTZrUPs+DjBsbGlRwNWWTYQNJ1bQYjPBxtBAh3gFiHIi79nkJGZ52uhwVI7
EUTEIKfsWnlscboyL0FElLWklaBi/cW4J1pKUc8GKLKr5YZIrjanjLTxIKCtHrkAUR0RefRtqPqk
1JDiSDhJcGZi9gvr05O2Fx1HiZ7JmOp86Bx7/rtANl97PY9vKZGnapc/8RS24udZqsDTzm5ttq3L
/eti765eYUeKM5AAtTEo1IKz1NP5hyReI9pZrsPhlRDAawFeHvK67FHPIvJS1LbTkh9gckzUZx+t
8JnkdmTeZXXwaO4GG1aksmMQD2tHGqy7kDD3VZj0ZPyhspHlnLVIN6df601DE1yrHMvFZT715FwB
KU/ITQAyTopueRoEv0+5Uws2n4rMScznlCEMusm70EcMMjcfnxaGJHaRq4khNXZoNnT5K2F1zUcq
M1zYnRhHq/tBlcq6oeHguK9+2ARmT+PLoVOw+0oEZpS8Ky0jxBtUbNg0j3/j9C+/JGaily5n/gpc
u2EAeupKXNmbSRF5Lk+asS8SOBtLBLphCBKARJYwm0j8Gp8x4nES9RYg1M6ecBUe4TB/Wz89P+xj
6k8YSpi6uoIVhbsdWFa7Nd8tR+p8APW0ie/PyYNyQK1n6eRhzTNi2yZvwcEih9UW5csB/FJdmCpy
LognYnx+gFoMFxSF3MjQ8YhMTwsd8cJe9klzUS9PwPPl/bsTDDlWc3O1pWWyXv/zKAAETlZXpdMo
3nFTiNHeoat3bbLSiXNiUbygjZdYRvg9hdSLMms1gx8YLmdbldfr68ebVCIOxupMUEIizt/kq/+1
MGKPOk8VdPsChh0bab+rNgBvbuLTWxUUcSDNU5JKArdYqvH9+D55DVKT9AEcP8HKlBou6dbHuoAQ
ZaI9fL96ijkvj3MTJ5u2Ystes8T4aM7oZIaz7epYzpS+3TnO1GvD/BcEGo062MqKACpq8WFS7jVY
ZAgnl1rSL2oq/OHH12xV9Ziq3/N3Oy20lPZZhqLjqUw6s6ac8aoJxhPs7SOUEv9J5w8zqEu0fNPw
YCMOn5lRUveyeC8RekIFBjjrMgPsDwBdMHRCIfvCVrZGug7wAp6VIDU2UJdSb3VOChZD/6lFQAD2
yg9S/RgcKxczA7ZimbNFYuHoJkVCkmUBIH9U0oud3oUymnfkGQ18xwJFKztNbnp1ALthXcxObJio
GUHm8MMb5izTRYhrQqAquczpvjFtHpZilkYSJtENbqMf9j6QWXhKWVFOpIpCgWm3Apoqg2a50FTw
R/nVmMidCUNP97hNpTwdMCmv5fNnbeXaYduPkGTfmdxede7zc/na8lNKdj+m/n6DepSp86oG5osi
0dHckF9JrFSBI6DEQJbs6dlL9svO77YtO3T9buYH/rBB/YUxquvAqKQkC04cmTrsK9KDVmBBWJLZ
pFxbLYXKPmXS/B2BprYU1GMBihuJm5M1SS1/itoeI4w224MbX9vNBJbjMTtCfqY4eg/2rqc0ND5g
NnIOiCmdSa+t14Hm/cJhrwadcDKSZ/ntX0NosSPjyxXFSDz4u6LZewsbP89+XfCXnSE2+K82Wh+Y
4wJ5Cr6NU5JVLNDBuvyBALHwoWSns2mvHif8lyZRMMENzV8HCcJlOeXOWynr+sFRecjdxSoEn7oy
jqWlOYAnTjo5PwE4b4wukOWB7wFsdvSPVo4vwXHIhdifgWHEaRsITHcuK3U7HTEYA6ILeR9dcPW0
dNvNeodryAXhsCpFwElVN2Mr8FVjqmhRcZFAvINBns1B4n9Fje7fK18PE6UxzxoW8ER881zBfxEi
PhqOFvEN0dHWK93LU2vmc6UHRsNecqssFmwfI6vxnsdn7I+HzchTAVD/aE/PSCAiapiOia7wruqa
J22AGf+Ps9rgIrowsBcbJ57F4SxuPiS+hBY0ArWx3rk0ado5n5qBss2pxBy2EN54+oFKTw0GUHs9
YBMb0dx+nRyxIa5cOU+pe2pXoecJTLhNMD52lDdBAK9FSIP/sv52tHaK0Ukbi7IHJ96CPfa0Vw+x
pqmh7OfVpO+nw1lgigATa38JgPJh/ZFo0Rr6nyebdUN70iaeucH2bwK7ZAZTD/1zHzfKTP9VKBY/
7b/VLtODRTomz6A8f+3zjhFQfYAWArz4Bxxu1I3kfvIzxmRHNEPoJKl6zzAa19BoSV7HaBxpM4Hi
ku7oL50GzPg/KzG+ux0MOpaG0a1akJpiYYGaeoUluxXGg1WUyi0ZWdXsubVlFTlRIpphRdh8xPN+
7Vtch3pHA7XT1PcxXUdI9OfeJJpI8Or3hx/wJ3pcbXP/yOS9kdKQAAOAYlMTzTLHXiX59njmCQqq
wKRcMkIlJnuA5ml5jNafYsL+ylYSBoyDU03RHk7Li4YqGonQhY9VZUXwBZ1WJ7HfptWvDnS6Ys+0
i8oCHQdF8aMhKmXfUnUKZdM/qvhUO7DN9wpPv+BBGkd8pG34WI5zEbehm9tp5CBsmBoEoQ+7zI0F
M+ePfzBnrjdYKSlx30D4WkJNUrCoH8vjIdkFvC+lXyeMEKqtiFvteynZFk4FvNdevKUVnoGZ9be/
ZytiMPD30PsiY6RzTCdOz0IiGZrEMss8FkTgL75lAhBAGDEZ9uxWCRRe5h2IGgnU3wJqXJdfC/lQ
t2zWMNzXA4t48aRXK/BWOuBZF6eOlAolwW8M/9U2Wud+fSwcJ24kj0g/vartrjAavHCZPj4YVgj3
nO+h3GUqh4zpgmIiy3+o8/9/EvpLSeArnwZwjWs9B1rHMGZvhsqiov5JPyCMsUTDBKwUj8ziRx/I
c8pQe4MzwS8e65WKnok3edrUquzWmCaZHDN+5YujdAF0u7GztI/tywKl7dPW2Mh8Qw3nygyf7wFx
amylYa6GhpjP13bygtsT36Ujv/xxHzUEwH+V/VSki2tu4MRGngPRlC2j9GA6Aa51KN0+375SROWy
Vbj0RxsntJDaL+WI/fD6IwGqMEknlpbfOpNpu/hO/TwAMuKXG9D1HasUivUeyAeMS/kwa4ehC7Tr
3jwKBbxNnF1X/WM9SrFArT/PGp149hoDNL2sanECWxm2pr/D48bQoFse1DIgjIljyIJmpSYBu7sb
PUCQGs2TUG0jW6xB7TjIsRzYoiscC66f2nXoe5oijsjJyP0H+BHGvDguwlNa94DWUi1tS/NCVJj5
iq0P7hlAxXULRUR4nPHc3brxSlORjl5uobo7nNBmw2n/r/5SifrpobvfBU19tfV6Y8bl1WQcMAMp
BRKTYI5vOu4q11e4F+kMYof/+jFwHrmhKKqG84ZGbwloDPGsLmt23eS4s6LlhsAJsI+imrjeQjH2
fJJl22CeYJg+JCRXbt0mWXHxPV3J0AS9PgCIDLH9J6IxZodOsOJ8sZjarpboGOiypx0C//8qFhs5
Tg+6VK6fZzixGOB6SJ3h5rgpTNW2g/jGUAb2v4kPQ6HzR4Vy+ZeR3G6ooX8fO/R1kNPjAF9epjmW
Jb1HqIgvUP/z6zMXYzD1OfBSUrL1i69eK53MJWGy+QF4DUzeUCb3sPZ/AJTyPepe2S60pekgiIKI
5aWMeo9zdblCNedMyZz3BOGonDquGm+ypVBZGndvdQ9vVnxrZtjMhBhAL4Npc9R9vxfqLFVEqshM
WJ8dGJw+rDpt9L0rkGFJS64HItzz2Z3MRNFTcYE8v74nNOJK1WmIWPFqPYi0unuwivXbAwhVcrIQ
H2P7/TwIX4zmdN1s0/jtMyx874n0xRDt5diRT9DPjuXDXdf+5vdx6N1g2rfEAlluuL3uvwLd3lOL
6RWhrB4lsTSiAM/F5e9Q4ZJograjeivqNcocchQ7Qs3vGCzOdg1Ra59jQXTRsgJcjAeZ1DPppiR5
TbRSJW9WJeSb3KRMetPd07KKICzod6bVYdN899RcAxiOHuhmjL05juuTztpUBcFnj4KwsAr6bxqI
lUSJ8pcNjj2huAcO20qWkmrnoKAscXSMBHqNx2tSdfTxNlGMtb+uxIOCZ+tUSFMKOeOEB2G9jGq5
U4rLSi3ocZ/2M5f/mGVBd3NeqA4jSImava7MxxAuQSeoYSms3KOeSZ7oIaDqs87SeYDQDPJpucZb
o2Aqw+DNbXJPTuvfPwcP6zUBH+q3bP7mQAipyQgsPhypF4U2IZO0zDGkuxzsCS8TJWyxb1TiV1Rx
euFhbAcWqX4cCcgafKuSew2o6gWlrq7dEy5vze59X6xvBcNUlAChQuI5v8eWqLglju/ViRp1hK7b
Txa6HLVw/eKsW6+YTae9ya7GvwGRx43OKnTLYgmQCA84Pkv37tLSs25iwOvMFwJPumHrDv0GuMbF
iz0IVOcSkzkO0AWx8UvprThTf2uJjpVQxCwEZDZWoKZm+XN3jpaNHdPs6BKoJL4yIlZYp+K+JnW5
gUWaLkkgHfleZk0pVAW+PacR1l5dJprqypfNqeljxvjg/HQhsNn9361tqAG5PEwCW4kpLQOTG8AG
xRIySi/qUFpDGid+GUnY6ld8En16Gx5If4/bNMDeo6j/I0ntrb4e4rZMMVAQyrs9a6KcXcTUkkOw
GcXnuBEspMLtbEv188jcuObbMl0Z+SWiSAKSagHv3GjmLFd/Z5BiW+PpD90t/74kKYOYu8NwF6Z5
L9yA2a/8oVFlxaDGOnWdZFBjiYKI+TW8v8TRz4nM8ck994E+M47Mv2hvpjKGB8M0lijHj2fwyoZE
AduZnFgGmS8k0MQoGJvbm7ZBEZQ0pMuf0ZF23lU4CTBgZyL2Fv+Pif/Xx9uOKWJ82pmN62NMaZ/9
am9RqhDKMtZ4+LDbJ4piWY3fGYKKLq5Koy8LISyL84rbd59RGsyEHOGtOh/AU+NOsspDGhgmvmwZ
ElsRCmxFqsH+bIpc7WamrpEJzSC1uX7Vy5ig2sP4v3Be8UqaU+S3/GAWaKlw55Drs/imcGHNnTnf
n9cnimGj+Ca4gXnrer/dBg31mCrt7zj0uc6B64pSYgIXdAkUtyvKImXXYbrXOfg+8c4boanswzd9
koxw6DZALmDOxCuYP5zrpAFh9zVyw1jXw6UzbiMvfDeR8FIzNfvY2YbOEERWpHPYWf7DZ72STPOV
2uK1MZ8Z/j37a+Q6CYs2QHtDC/2BlOgCiS83ZKgOP5dsxhMzV3aEShgc6/fLZ4+8Nf3TC/VNzN7N
aD6e4sboRzS0TgsLM9LUB24ujuYQVVtAu4W1ALVGudYrMTXTZfNPQ6+9RfdqngLLx2/Q/yqIRczS
99wdAyTpzX53R1XkiiQCo3VhzpunqpO8N1p26S9iZ4d5F+9tg8CL7EzQyb7m+OnjOyemgS6fVdvq
Yn3rxTYlRmhEvwyv8YJVrtTY3FQPGu6tdP3d7kxl4izNJe+7lASUrjFbL6h2CdAMKwqaFPwIR7GT
3EmhlPh9VMqCAX1HZcWnve1indgextoRUsegRsrdWxwMNQY3N8hvvJ8l0UaG0ZpzAlfGaSbi2lL3
AoNMKygGezNaVdW0X8jYF6p3zuaFFEiRTvlYADoJ04/GIvbg/v2VmUFBDLYs+wttx+3+mNAFRyHf
5yCImKeOXUhJWElJbnA8wsUDk7MPSiYpa/8YBybsEdd6o4VnZd4n2lJnGGF8IsflK2pDSlGTT5LU
rgMmkwRLgA0miIWY+Y27e2B6qgCVC2AziwXxxhOELdnzMilFEwNuiYp7P1qTg4Mx+ECLq9RBQuVb
8RI06bGMBOWCm1HI35VEX17r2L5mS92c+QSkZWjPrKRBFI6cNdNw4YHW0thUPHa57XWgZ2mLuRum
XaPSP932cAFKasBMxyGpGtAKTegEgTzeWVj1yf6IEFHwSMgklI+hYG9gAzVGoq0/864KnJI75P/H
tHG0mDvKnB2VwZWrIlFklywrJgvFZFgBMCIRMaCjoVW+Ru2MF/o22l01x8X0Ss2Zh+D2/Z1aq1R7
nkm0tDXbHvg4BXa4SWX+SKkqyNykLjIwakxCfK6h2zjICUMZFEJ90O2wXdr/sdrDAh3qWKoxu1lJ
l+9gkI6htIv4Yal6qDIkpP2I9hTdkQp9XxBgXQon3pqfphoYKtq9fUA3vsankieBIdrjP5uZh69h
5AYIwDW59P33+kc8lhh7sD2FTUKUpS1LN0flNHPOCkorYjHYbLJoRIB5uBtUeuuMm1kA7SWhjsCF
nEV6liLBl+g8e92fjgdZfiaAbVfbDEDx70GBjwNZc1WDRanE+enlVsMvS+cqDUVPGs+i45CILRrz
yDP7gdN9yjDqLDDti4RU2530ykExG85RgXn9mWJ1SaHIwrdjCdLKJK0lke6KVo1KJJONEVoW3TM8
F7hP1b2WMFYJFbQ48JsXMTm2A/AYO6gw0X9u2kEy/0KV3uv0QMOU8TqCZhookOajSL0WVVVX4bSk
pNjC05hpS/L1DDNW/URzF2om+ZEAd+A5Z3+GK9ryUnWfNqScsDLrHXzK9h/5Tyq/pKxTcdkGblp1
WSp24cWzNrdA3fvktZJ8+3dVIZw1fgj9wDX8LOe8TmWiTCBUlOxsHcWUzidlUFhAnthia9V2UyWJ
Uy2qBBoJpDAV565yQG/1eG+wX3+MSdiAo2GLxkplXfivckJGSEVEpIuDONjCbTz06aDpgBQNhv7z
5HRfXsZOy1iSOypDHMtpnelPK+jZQzLZcRo/3sinkIbFM8p9yi6FAkz/COEDaednP72R/jysNh7a
xuqcz2849/0rjCO1XyHpVUuHTn28AID5r/jQnlHdIHs8nHqlidPv5Kw3Ly/Iv1n0vaJOb6652Ehi
MQXTAdtC3gqVkjakUoMjoqQ8td4Mai7yxhZQYituRtGn0HkiiA+fBqU81bopw8rKMXsCdlZBzJaI
XQCWgEBIEzHfmxNwt0Hv5He9dw9zf83ijjTMh4VE2KHUmDR5ZfxDFqvhEvjnljISkSeKvQsnQvOg
qvRmPu9FWCVNZSqbDtCDatpWuMz+efyOwY0TvRnaaGfMPputsO+uwXzWLLNunsjdpw2T5tZQSPHB
MRKQdKIrIhFfE6GjFGbz0AkqHYx69/EtvoIKlafqBgzMEjfU6J9yythDh9e6aYW2PVsjD0ej+nB1
w7go6Eha/HLF5y9nvySx4pMIafHZLG4M2+OWtURDZCijT/G419w0C8HRVfeJ+KI7wQOpKcA1f0dp
CLhoeOBT6x0O6ksYHIESAYBroE/viQdCh251sM+cqcoRc+ATW189s/Pr/7dAAPiyaHmYCfop5+W+
Goq4iKXznuNNP9yCPgjzSVwTwTnqvLTMQRRlzUZPWYYIImHw0m5LAi97qMrJ/bhxM5/bcc0k7JiD
gANa9Imaqmxy74vgT7TZX/7YoR7WjTWwBhgaz/j9pbwXSJDowRDeKsV8zs54S9EN6+WvuQm2awky
3hM4gjl5lTcl0RCzJuVJd2i2qPpe3NZ9Q6D1DEiw6KPDwUan+OF/p0a+M3f+HBHxyNcwpLb04KNx
A4Ru83W04WQfeQlH2AMJ4GKrOrEBpRPEZgHSJ3FBgC/dFaPmTP1rIDlX63Cvt9/RaYOpM7LofcmB
KKNmnbMbLf/cY/GIemRWdFe5ntO+/LeTd+MyjZn4Lb/1x+Wo6Idvvfz6aYkeNNAfKRG18p7snFAp
AejbpjXNsWJQsUJ13PYFr8D44dvqRsby3OooZLMVerv8dI7qeAIgFxu3UlAuDjG/cw9sMdx3O+Qg
FjfBUCPNOOqHehs9adH6I+4qUufEHU3Vm+46bgPCBcX2/Sy1yz+YXEn+3yxHyiDBmWnj0fkwqq1v
SoCIDSD26ZtHL0xHg5EpmLJAXTo3sYMeF96SsZ3y7xxBS777Q0NksxSDw9qY86r0X33OQE/fngVL
36hOmx/yyISB7P5rvHp+GLUzXtPDudlrxsPw7rmSn/Mpld2Z9oCfQNbw2WnABuosXkCGNDr2bQLv
Ol2ntyTXMJ8E0BlS9S6M0MZS31/C+McpeTpbrd2Ke+tVBNBPdEfhzpzDvSyi6uSHQiQuTXtUsvy9
u5qHNgCnDM5GWbXqipgJnID8hrAgdrdeAQxuT+UjQ38I9+ZfNQ3JwqTJ9BngoHz9l6Kyn81sIT8i
WcJ/CytiWgQokoubt8S7dz4wrZmlTJMUbI4soSBVFVqhT0hmOjEiT/wMqEuglYf3fGU02EVP8jq2
bkWF5EsAKuBybmaX/OCYoDjvn29NgHXNjDh7S/IaAd/iRX2uv3ZCg7kfxbXQDapSUm2TF0t9u7eq
cuZyLrEQiL8hTN4fl3ZmVnGTkmb3COLVL4Bzip5CRCy1F+PKZWcHofeFm05ASJi15332tJa9oXsc
Y2XokgsarjPKpEhR3ckCpFR49SO/xaXHUW2X2ZmRoHv5Mv6fI3Di9Pc30A8pThCzsGVDxgZdQa/f
EQEC50QpCDGJjSY3YLzlSeS632PGG5oCXlgGb5eJf98k0K079WIYjwIv32Al4dcxfzcJMI00oiLL
W3ISy0FZpVgnHJTWT6orFLiQkjetcYp4hyPUNtkWbOjCQ70DyHH6Jg0xROXEaXbVi9ri4yzs4Ic+
9AT8savlVPp4Si0oepCntuAh1bUShpUfKgIimDCd0A4HqXFv7okPRWi639yEoKl+ke2hhfnbiFFv
9js+umsICq9gFdk5O9dRQeHbh8G6AxoJ4GhHif5+TsihY++TpiIW5HZWuabQ63VjWlCJKawZ+6OL
JBmkXXbV0UgHiVatFEBp8Bv2SiPHn3cC/cKs5xaZm0cogWzmR9nPGqij/eTSGuMsmZIEzilwo24N
QkQg+Af+8K77xAgRJjjGN1J4j592UvXUkqM2FAsqNhlj7jQHXkMgBv8RnQ7L5+pD2DnSPHb5cRcy
oYRiHWNVPKAqKf20j06BBFYK1t9l1BaNaBZaAbCh7NcufXSGNh+HrmA0dAW8F9EvumCeBw5GZ9ZX
0h7zVVjcHQXWbRQh9FwevGkH0rLjzJg7a4AlOVteaAfoo111Exk6HOFEqTKUA37HKM/75Lpm4JQg
q7ma7wzH4GOLPgzLGX+ykza8ckbpYc+wATYZM0IGmR+WHs0M/SS3Pd8kqZj7tFG7RGEvLS+dMBcL
8vW94mgd9ISO7OFtzipADBQiMpQXSS4JW/PmwNnzN59Zkc38Te2hbKu1wdEDCLbFCfMNW3eBZdy0
Syx4OpDI3u/jMIbqGLYCoy1zWGJ0pP8rvFI7U3a3715es36nchlpMcf6ifae8NnC0H7tV5SthRr3
+lWVaC5wEbZ1PnrVR4k73VJyqvVKs4isJWHc2Gn9jQteJA+E9+/Fe5TPN0rAthHB8HT+4iG3uigw
Vo408IdS/jllUyk7HKuufJv4o4qEoLcojkiNMZWFAL3kEhdgHYqAjjoU5nxgzUucqQPy32qzrXiF
MCgtzb/z4U2pdUsExIIWjfZD/5M6kzgLTiDnzxf1HWF+Wjwfc9IhuPk0O8cG4SBk9rp61GkfjRKr
aT6V/MXtvQ+FDCJlf+10h+2ZnJ19QVgRUNm5+yKdEwqr9iP1oMauCPBL3YZjdpuChRlRPppNu0ax
4p4syMPUdQOL2CN7ZBjIXkVJAKM4g/PvYgwlQsI1vdjZKImTQ3LfAmcw1evfeYR/bDd5L4KvtEi9
NTCuYc5JKkumZOk0ieaBucZjo9Xu7bK3tERWDwLPatjamRjet9wOpkbYqK7gLYYjrkA5quVgqVD+
Pxyu/oQABZmbqc5tu8P0EyD0NTHWi4kjKXumUKCMHn8RhD0BCxDZT9ZiqOOO6DXWgDHCtVBXnb5r
Bfu80M0CO7VvlVjupqoDKKeAwsx5BFuF2wYoEJl7Po9i5oETQyRU9+Q1ijybJbcC9n4uitFIlbUn
TdLiDo4ed/ezem+8OblQMioHd9GtT9HmyXlqdlHPhuzQXtSdmTOa2R0VUBcWTjwEEvT9W3qZTKR7
MI1DixKKwseJQTf1ouCWfpxGakbXT8gL5mIXsTGWQb/0Yjq0KOsazW3c/z8S7A320qJNxcbkYL0X
q2Z5ej809RFyGmOhUVNBME3S5Lz4BRKg4ntNsUgUfrRf52o0v0XKSNYHWmnFpLLnkOA4eb1voH+z
PzBzH/anT8+niqLp4vCzzDuv8IWfH25sxV2r3uxuzAn9COXG6xu1odXPR8SG/y6XKO+v2kDT7VMY
9BBfEtIi8JGTF1fHVBCaSI3oiuilKr2wimBFQ7NI1vpkhOnY6K4bbZ4uZKQrfElnVXI9RWmPQ34d
0UMglQ7/WKgTnWIbOPoKnQoFYK53pqcr5AlySn1owKQvCVlnI47iKCubJOu5RfK+cGe9qE466zuf
w232ecY7XOZNTBuxDgKIghMCtMNpp7gQlYGdmDLLCRankXxGhkEmfWGso/Y/Px/DbhJBqb01yOO3
BrIAgZmmZsyS8SQVNXkTEPKhkeNKJo8tsIuDbhX4b/nHRo8bouS2fkJp8HSNbmfclTe2nv5PRBuE
KpvFr3bz7ObaNgzcyImt7SspBET5NRA/rsVMrNlluVF8+miSobzzNXiBR443O7qI9alyPGAvZNZy
CdtXuyq4YgRJYGDdrxk+HzR1jE/uQJ4dezh//RID5q1us+JfDGu9Z6k9zrBzKGueTCYxTrZ+6yVs
m1Pe7uMEYkfD8Khc35tBaGs4uEFWn/xSHhXRGm6N+UWgKB/nGHHB1qtvrj1N5sXSlKT+MRXd6Gzb
Z52bcO/SC1mp0hmu+cx/dTIYlMlKullnYuGRdTKYyTMQ4kUmkJmoBSvZpFWMD07kbKkH4sWAD8cE
s7rilM2T1/0AL3RMlLr0vPwBPO6deZdeWu4Gs/5TKN7CxRANA/okQW/IILVbEE8UlmLaE+1OQwqw
W6P6vc4AK4uMzQwgNNO2oTewI+1359If1tmdK4VlWm5+4CHPc/Rumx2X6GmW9wI/MNZAeNl4rcGv
YVjfeEj1YJXtAgJi9ws9C6VnXm95j2p4F9lvytYSUPpvwpVmZj9SH6l6Xu1tDXsYfKSAvw5kj5bB
6E+UhxJRzL5uuodg9dB5mJxp5CfLsIjW0VMPl+JjOsaAtGDKd5udnw0tRTiy5W+CySpbpDuySdYB
HZH6+KFEZftakcddyJmL3VD0uBWMI8rZcvJx/rL/oDadtQ2+moIn2C3F8Q506CKXgZajxcFSsgTg
DIj+mStmp/vouKr9aV4aDS5KP7GFvNLZ781l4V+MSUxQDRAWh0h3ooJpImGTVsz7QsdSj7YSDlHT
N6lWxKYj2VTSldLJnzDtQpL1cPODxjHe0YB4E3vKnHOOR/8d1jmrzdUVe9v52ciPBxYW1VuxP7ru
kch2DIyeyVsu9Fqjv6zOOef3DpkOqyNCRynMeBnpouF9RDhNufMQfEkG3EquXtR5JApxBpyZsPEL
E5J6PgFTuhYoi+6cMgZ+D4blMT8u+ce8OW+YXy93ukXp7+HhcPHzpmERHOO6Tbb+2Ue2bSJeuh5N
kyHp0S5FWMffd2zN1Oa9nEQr86IsXFezQC6v/Ee6QADKSbaAeX2Ccdql++dd4fiCkA16jzLthO7v
6ec/w+z6rjwscGrp99SaVRm83h7UwIqE4t/eLey1O9RmQxf2K2GNgfjGEBl/yUgwdJm5oKaSjKGj
k3Ia/YpIK+FrjwGqjwXg2AUFxWt+on1zeh+Z5h8B9pfDvw7ByCNRT6PIHt/6Gc+1uAvJ2vDIOsI0
6tp44sCWHEAsYBflNo6akY4fC9V1YD+CDo6rd5Ax4CEKh16/jamRn0vbBLBczx0EjTJ57YEfL327
w7N1uQd0byjpfl6RJJfHznQPxRxjmGO+z1FMgF6SfL4GSchYKVSiV3IltEVQbspZBDVDSKmROsiw
Q5UdNjnMOIJo+8cB/2hdn80fRAJf2OIcytoHrb2O57cbvtGNh9d1qBlTSpya10tjftLDhSGbR0vr
FCSCglVj5Taczku6TOYSU1zAwLco10wipWd1IXjn1IsebfPfH9en77yEu8PUzBmmM9m22cVjtuj0
JxM01DkWqkIsza5yRVXE69mBy7pOLziP08O9INfUmttpMpWj8Koc4gPG8gCuJDsi0xgjawKcL5JO
0SGNjP1YNFGE49XGoHa0NCV+ZbXXYI97V7rYpKHRx1xh4p9A0oKNrV9AGdsfbLlo8BADE1ggdtTJ
rnp2xYQnW+xb3EcrISyn4xxem+UxP+zLSSj0D+i3bqz5AdObGShzfCwSkXRLwOPWvUPli8SWe8Tq
JNlzhJbL7RUgJ00VmIxSQmo6DQu4woY88wmb56anOESNY0CrzM/zUtzj82JFb8Ofe/iw//4820W6
Hv0KBEIVyv40CHYi3P59jU9RcesLohdEsiJwYizXsgMRnILSgQ1YGWMAlKUXjJPu6bdJEjdS3OS7
pEAB7jj/1xyZjb9xQoHsNuYgjUyHqnX2oML3yxgXEpOXfkXwUnA51ltjjn3lrkU17zqzwYv4P1mY
5yfhDd11HVA/JE7gYg74w7+2x6UJE21XrKbmutUc3Bso5IBa4got+Bo5TupEAOHZl2b0FHEoK1Gd
NiazzdC2i7nKBNuImdRM0NcJYpujiePYqw7vJQ9zykcPwZz7B7B8/2iQt5e07QEpZcjxYi58FJzJ
KBkI7ywanpkOmifasj40ZiMNYerDv6ohC6JjFcSTQYpbH+DsP9Xp8sYSHirNxVwdaP0PO5UvPeOB
8DJDXYzxYbcaoSPjzzdhljeqDt6/7zwJdN70kdF8dEa15G0mNsurp2yen45D4oKgY+0R2YNvzjGp
MqbC59/LsH+hmTK7G1uKuNT5i/NXaGPmkIP91HgfNRoluTZC50yG+oUZt/JpEUSuRP3Okg2cwiKy
AjnQeGjNV84xrR6j113qQEvutxYht1zphHg/7sQYE0l3R4qPPT8ObqxHRrdHp3/SzRFEotB/g8bX
/Z/waFBnOW3NeIHuV6i8oHy34nLFUa5idFWRqW0BokQ/Eb0gPgivisuW/iXVc8yf5AqYQv6W2XzB
K505I3F78UxQaC68BxyVmmFoQNqs4WkvkaJ4XSsavftGiDrCjcEj270IbnsKb4iR83r8RjCSzoMU
3RF0mnVXV3knJmaxr0k1hqa7fyunL35J+h+Zt8l8y3VuCLdyzQ7ojGxxFsIY6/Kz8WYhkbgciVjL
dD/zf5/ZYmjha3UPyXXLCytkFZRBH6Ik+qkSzEF7xzL3G+nJwi4CniynhRlBPb9xdAZDgh+HPF0r
Dx0L3BkNPl8ISmFVE8fagS8P1N5SvwgFXnDjGQZKaoni5+mY7tSHychi+/XsD7Ne9VXS9b1/6D6p
3Sz/uPCfNvt/A5yYkDWNAFTZwR3GbnRXYxtQv7JM2GgSW3MP9ilcURA0WfnmGKP4OQcWCS6ZalaM
yTXQ5dZvq21Tqp0GdAGtCi6YJRt+ysE1rrKtFyvOvAkCAwKAoyYBjPjImcf3Qd7w3cN0073ysbPE
lDuXfs3yp5ifQg0ZklyaAExmM7EW9GmfajZZ4Kdgm1G1VOd0C0Y+kv2vz9jMmA6hk3NOSGvboQiH
Y8TBg8QHucj2mVRS2ZyN7IdB+53zAWsIGFmrACFY4ofL7K/qwXJ9H985Y0AzXRkLZdO9zdpjOuRY
jcvduSYuL9sLoruC1mI1OHinuIiYSgYZRnDKWx2XoeOSyTxgpseLCsrxPMr0pphKHyjn9gQi6yJ+
t7hyw/wU1IjJsTG/n4P1gKz8XdgC5jchQ44PT+KkKTosXoJIUb27yix7BBYinqwVHCBl/5g9y1H7
gVObBtu2UyWThegOA4zJtvetvat1lHPnl++zVw2GGmncBd6WbJdYatREpO/F+cQblsqRZAK8yw6u
ulA4qJxA88fFdeZg4u08m5MNpb/BDjdoEoiIe1egkdbjpEe3DNTkYcyXGkkdE3Ommg/eN+u8V880
ZvLw/E7sxnyo/MIydUcKIxR+ftQOUy0HPY+rReEy35aoVDURWuauSOJ4Y0Jl9GoD3Yh8xIGiSBYC
UPxpnDIVTCfWbUTKeLSQASrn2hhGg7WnXDPH5aTAMSvaOpcMJDV67rdmuF2B+08pOR1Hb50fxYeX
Wc0vzy7jsA0t+Ppr4fg9Z/25RdLLw71Jr85XFePuUKJl2uZf9i/wgngtFCCKqE1J4+6SLBUGNMFp
lEgPNeJOSthb/1IBZWSuaODN53mSMuHDejT28g+UvFL9jwoxnqyBmD7fRyiLsT6rJr4k7fb751XE
tweRPCfRQXEoFWOfhuT7tTa5B8CejUf9Dc0k5wOWTZZFnoTEqjYzgLIg4pR3fkMj1r2EMsGql26q
lZ4X47O27wVOTmqFV2rvlqLucBxAO3Xc8aDiaeK6M7eVIPF7Rc4W+fwEl9m1m2RiVBtvuv5gBoob
5B0wwlp+A+iahePeLyHbb0iW/DITzJ62E8auLLMEWUmuCIZ+J+Y+R331ClQgUo+rmIY6nKm2rSO+
io7NbudUwlE5po+Ted1At4UwdSs8FV2mgXL+phskykcPmB3XHtae4C/2YDmGDhOhWJhFpGhH8TJi
Vjlmi7/WCMnjCwJ3lhchD3NGEppm/v+uIZb1a8bB0+IPSYK9yL6ViMJ4V4Ywt7mcp2+sRybc0ESf
e1QY/WcjCQvKaTrBj0WRMV5eCk+3MhFD7iyVA+6xdEkkFJLLBb9g+XkRmRIkx/1TffFnC+c0nKYR
UXCuXJz+CRXJBOIIUQU1yZE741yKS42UCZIJDpLVkwRQMrwWbxB1HGQHQwcIRj2Q/gKVz4CF1nWE
WEdRe3CM0wVN0hiZj+aXByjGT6LGu+mZF8cRdEk4qXDbkBq71dAsPOhbLBVLz76CQCXPHxYLVf8b
uv18CyZGwpSTliZKwStK27XbvcEuCfMyO/tq1s45aWti7gk3EH3cuYw9/BFbyv0KFq8rNzvK/2c+
6ZdXzGNQti+bingUQYV+xLPvfNDk9GFiHa1PmNLcDMbADRWmK8wtI3cSpQ6ctYcn0uPvuSdmeapz
KqqzTYSNSr/RI99vydv+On2Nzl0fznLkq5l9n5XUtVBPpfwmEnz0QlWlOcU+D5a+2c0oFaOZwX8L
yhFsE0yw9hNThb8i01Bs1Lv1vQMuk+TTybxgqu6ZwtDYo8U6AvF9NHEGQKvWxVoiWsYP5aR+jHeq
5HSb1TFwT+msL0QpamcvnAGfz+91FbI3y1vSzrbW9A2k4euXU2Gv45L27gjblqatWQ4mSheZIPz8
LZXhWDmtYFlaWPCRESDo4mETBML8B4JqMri3dfUgMD7ObCfBdmgQUKL8902rJlLQd4SXuKuiuN/C
3ks7T0WCZCRuekmlryW97M0J7c3HUZN/mdcG/xJukqTeKqz6Xn0/XB7Gih30ASaLEMV82a8IB6f8
tVkgh0R/jIYcfeh43HEwgB7Yrgs3dxpOdwPUFnXyS6E3Zl6mY8ohtKDoUgi1PxKLVrjww7sOD2A/
I/e3kIIyQ2VhrPli8uyKeh3T0HgDSo1uK1K+PIsqHz3PUlgAayVRNAkbcd7FnXcigFw5p6o7LJxI
TmMh7NWBLl+Sb9vAEgffvgAYjvOz10c9YiDxYKqzpmG50YEDHlK9ZoZkQlr1NjgC8wYupRQB6I03
m9UsG+0vqyYr9oUgThR3kWjOT2oESAAm6JmnwmFntMGTfFi9I5lEw1mGzxL5N03lXOZGU4zCvTlm
2X1UxXiiZvqK7ne/rT0iXlfGhkF6TpsJlI8PvBkS5nDlXqGvnRkURooHrxu413GMaB2t6EoEPotc
ZWK/bRo/zjD0RE8rzrnhmYdC1Vf7EOB+IGkt4+vK/vX6/+wQSIXkM4GN8gNoTr4i0Dt8eIwnp4SS
tEz61sKhnc6XNYuBxQfFIpwF1+F+givoj4Guv+6KnedERpVHOJ3DBz/tqG18/Ci87FleKqzMEybw
eygvWSAh0jypTy6At+e0H9nfC6OvY/cgjAO8J7NY5bnSlsfS34IJ+medutQOmDY1Rr6wfGpQXerO
gh4tLGaa7kIWQR3CjJeEfUs1zruUvTpdBvasiHyCk1SZADYsahBIYp8Qp2u0Cmjb0F9vFL4PTh07
1s3uOSUp1vk4oTzwQHq67ASwwP1pVFuJL6DWAPhoKhSf+Kpekvs9GY7G2VdM6A1tfCku/V8I9F/J
zb9iX6Mlct4Dn0ybNehpND8daiGivaTkhdzJZMVe/zl9DfQdxXWsRjnM4BS+QLUkUQZQiVqr7RWP
mT5Yi7LNdeKJ3g0IXf6nacrHIm5RjMbm6TTHM0Eybjp5vmHXqFcY0p2Yx3kC76U3zDU0VpJjli5u
JVrd6fs0SwthgZsAaS5ADFafes/y2z1ULq6yQO2RDeRcMlmhDV6X2dXu4N8iVx0dHycpHs2FELnj
0QWoCe3XqYJi5hlpRM5Y9be0f3xW6vuGWMbluwG5aQFsSlGwYK4QCXHx36Cv89ihWKBaZkL4xVa4
xDQK6Z+HzDjxsnjvR5bMRusMl/qYdj1dPIcHUvnGmf7OhY9ZvPvl03Dwbr3H/WCo07FgJho0ICqq
/JXGyARVc9CvAqYvtWskc7ihkVQxccT4V/hApiAyu7ALSKEP5DBfRk+S8Ob7Rm6SAYmbVPC9yCK/
HIyXvchbbUy+b1hz6mknmYfCATAENTDQtaT8HSxwUdZzek2Etf4J9ggXB/jHETzTMsaUf96pcThq
csIj9DupUqwxlbCXFPtSp5E10upf+C95O8wFhenPLm6i96dfNs9wgI1zjo/36bRyMRO+v6U3K0Jg
NpUpOWW32cksaGb/kXFrmUx8xNH92gmO0xHty92ejUJMdQXsGAnACK0M9uIiaPNisUEuQwEXV0S5
bcuRzd3pTx1BFAvfa9Kos9VN3ALCu4ZqAvzsPYJYOfrQuQhOYhumsyqOSn3OkYsgLreChgGEPwZd
REQBPdt9f3ygRHpeNX3HOftw4FMpaUnectRJTul4FRNROXT+MDoJjc1ua2525XmBxilrhzkhp9P4
pFS7HefVnCYqTvYs7fXE4Ymv5pqZJ9Ifjj3kioZCzeywc4Xzxwc+ejafLEF9GYMwcc/+o2lwyUuk
XcCyPCnwQlMxowPA7YYeQPsGRUBeqbnRp1sxWmJmouuzTht+3nGvf1LVMVYkXyW4vI6074uS/Owr
y/W0I+3BHnAJjxnoVIsoTp8iBzLvp9gC69HU1iaBGYtBYr78sdRCBOIe0t/OPVyQM5ZXyASv2/sO
ASRT7ClbA6Y7S5m0RNgov5NcqksS1dJYleHFwiL8PuZ0Hn4KBJBWlwm+bC5EgYNicr3ZeXG93Gky
DEjPYx2j7IkK0CNCDJMT4w19ltBLQQpT96PANPP+l1hu+Whuk0ABiyFQyRWA60UkfdqpsOK6nPj+
nBv0KkZZQl8Sds/UpOdxqHcQ52L/AycFM9cxEO0iCht2He50zYkAah5CpbLvCl6LO2N4+S5PDlah
QM7f0h7QgDuwYct48IHB6SjCH+u7eGyZNnu9GI+vfDpiFyhh5ufOLceOL7d5ORvi6Njqk04djoPq
rjR8eZ7rU8V2Q1ygD17on6YNfTJY3U5gJQaAk5PviIxD96/OkBqwngjjo4eAG8rLCc6JcBbY3e8c
cD/faCpSYj8c+Sq2b/9IgV/mpbFtvoNqgPnHLbsk1valSC8U/y6JYbdAJu6Q/HhCQrvsaA8lFjkd
M7Gvxtp13K7HvNDMAYlgt6MbtHU91U55/wg6nUJ4/4r6Lu/jVppQRudMT5djC840lJPzOMREiH41
nFsnEF3oXMNvgj1vOpk6pGy4RVgg/CcDy63BuZXJa/8OJAkM7ME2CAovrS5VdpowK8yezGDYA5qG
lz1ixmtnjdxL96YZrUNSFV61IEXsCJ9UqT3qMO8C/0+cCESYPh56k3cPAXpQIHVGBIYK3/fEBa08
AFPROfuoReiR0c8dqaJwl5y5U/qbIWxXrlsGTtzhpjajDOimzNRrtUWiIH3GAJRkwFYuNx1eCrYU
19caYXysY3UnRKd3w9sQ50mtWFatcAdbA88iK/LVeajNma3zEdqeN1u+yRXsT2CSBpoL4RhyDT/g
MECKZJ4MgrX3RZAhkHfmenOOcuNnbhWlpRBDJ+YIEEBmxm8fmN+cL6jQOW5b5AHcdA8Q8WIWBGh0
5WfuQGX/9UAf7vmt5cuir0WEiaDtiD7ROBTqZ9iIK6DUsWk8t/QEOtC76dpuIY9kQ6va4jUdm9/9
fPAAXFFQG6A6LWPcdMzXABUrDxOg5Olua8/Md4+UUwUi2vJvIPTN0GSjUZ10gfJywZ3oAUNmLUrS
1K/a9C6KyoeQrRKno+m9RA5g0qB2eiyrzyzxmtp7ZWmuc6zD8B20o/pSAoRnkuCtEh4oogE+zHws
ioSuPWaznMPqPZWURpCVT/akJFqVVcsMdfndvuM4M7Su59wkbF4mtHSygYHiPVMUmoq82fbjFj51
HKnXF0S5ywZM7PVl/a/x3wqn2bZzc9+Z8tN0fRmuni1BTr/QgFOPranWwZM+aW/Yvr+RlKqYQcwg
u0JWTbAG6nIFHzxvBHJdoaZkBxev50h8n9Smn6jzO1UnuMezJL2nH38LkDh1LLunc54IX+phDCNu
vgo0a0xrXqWOCgZAwQdNnVIHEpTO6Gkfj87WT3pn5Njg8ZlHa7PAVehBKynK3zkyeKJv6yjx9Wa5
VQkVeVwLs56fIizKjCPLjSyTwMd/cDic9wx+he5K9rYc3rOYNa6Vd4qW7Lf9qbI1RGdJETgaTLeH
mzJFPBCAaEhbynQmsyWxIXEEtSnzTFHYon790Ljxn8jNZWbGe35nthXgQN/QOoFO2FQ90IeXjxBy
gDK1v9fA6e0CF52RvJUAc/HYIVuXkPkfUvo8oIpurDWH0ImzgqWhy65M2+nsvp8EUMqyIm9lAV5o
bI+PfT1CgBpXiyt7B0Pf5FfGIWUHMqXXR1doWI1gRc3ebaMCKORR2Fy/69S5bL9EeK+SNDIMAvCs
LMFoaGTRs/lLonXrRgNj2SabTOKOp6f6LG52IGX04LomlPv50dKMIngPIpMxBvssFvX50X9J87Ln
L4KMXBFzXw9jgxT0o3j87Hnx7Q8wC6Z+SNbeTF/47nLEnUOWZmBm/7UQ8loF8uz11ode8L+Wc5aB
7eFhN1vG5md6hNg6zG2TINjOknUh62uJBN+7z7aUUzH1DnI3Ze2dhncfzSzaSlCUMw+CoOoMMjqu
fJkxNVGsNU8tn7lENtkX0/LOq+PMhJqri/ICzWqoV7QqPh+WUf8K15lOLx2ygs3p69cjprMyhW6e
Gm/2MdIkPjf6F0T1K/A0dZJun141XiJibH/oVgV49LEEXAQVcRwmkeZKIosc0xJPuECsL6J4sHi+
tcjLhrQeNHCrArecPac9/hnFZ6xJfWML+oPFAfxWcqI8lnP4ja2iWw4U6xO+VfZGFqmZNyo4NU1T
hNQVp4rjPlRMDURGTqOvDiAPMOi7DwvXu4t6IfEGe3NuXalc1MDUwPPY7ck1QT8Qfe0tsT02/+F0
dZqr7VYQKOyyB5aI5oeGYQHvjez9fcWRkt+KmwClhy55Q18xtzE7DSfbONsfszEnkvUf+ZoMqdY3
B17C3TY70o+aMI/5kbV24OImzWMBkVotvq2BFrDNGptHQux4theqRtyR1BGOFBLYB2idlGdEi2mw
VFrPnd+F3QQ9EMTwZXf2bvxoMEl/+Xg/3mmdsXDpHJdC8d41VakP24w9leBR0bfOZXFfkwZf9Lvz
ZTi/C7fDCYcqcRCG0C2snvN8BuPhrUhWTuVknR18y+LrNVR5FEBJ7j/o7iD94gtonATJPI266kGK
Spg3A18VEMBc2NgnV84qWrCBq24DurlU11Gzguy9JXnz5kXQ/UMiJUc6ScpTQmcxod8vvf4PEmez
i3pCv7mim+TZ4Bn6Q4MqpKVTCpvd2Ja9cVz9WMaiYDLNxTXujK9sQOceEfLpgd5pHeo8/SdyBDvb
kKsjtZHr5rEeT1qkH/+TfeBp0cZD019hSkgk2gcokFDTEybdKmJ/WvLHz7Y7VPjfS2yED5lJsFAY
8r7po/nohywezR/0drop3hoNa/J9+Y9bpQEu1IA0TwAIQSLCzAMpGmdqnkqO72AUrWXNDvirJfuW
6gew2e3uCDz2BzTedXNsqkArK/pbRM488jRIbF20UFIUQeennU0/xgAOzoQ/7OqYcXqmtdNDgWAD
bNM+DhGfUBb708CCzv0PmlfJRtjLQdlHtM6jPRpqYzx1uH68YOIYvZA18uz00NrCLrkfQsvf4ZQO
pCjwsXe9+KOUj5ST1Oe9cmqvu+3ng7Kl1BshFm2bu3fxZr0gmyIg2xATj6jN28tjTlvy56aQsj3i
dOkfLlhZcvFSX/I/8ly/MnKXZPVBN0QMPDwyyptmdk/p/XIHgdx/8Lf5sM/jk9wpdNwAPWCrPopn
3RLvtodwrQiXCjkj574kdzHBpjfslsMxnj6wzcOPzdgS/x06cdwqX1PabXxUoMiZBgppEJnhgwyL
6b0JgfBDmWfnD0Xo0byqJrY1fkIRQh14WywH2juq9Dh5pop8hWwgQs1Bf2PgeWODGS765lwrPJgl
Dm0eGbHMpXiPVii5/7fc3HyOsvavk0ItHOhzhHpIRAmLCGGAjHfrSCzZIOTA9P2uldk5IX/IEORb
qzI8q9tifgv7s2mpQhPuOyJxgtOUethNXfeaApSx87wSwEEzXbSlyHSniZ9L+UJfV39uq8+d40bU
8l3C4lxsJyeEgpPA7IVkFbpN0JSwcLLzkh5b2GGRqtVlTZOgwNNVB5PUHye4m+ksHm4fWFiIjRTY
r4TYDYe6oNXwKTBnV0zOZrhHhctJESvuOwbTl63lD7kt6gFJ1eeAX3daP4JWGJIYdZjhN5UIshFL
I+Kp75xnTj01XcZ0hnDmBCc7ZGuGUTGTaR44gH3vatMILBP+OKdsSJjBP/VBeCmRxxCrpWLXI79T
N4jIZYx3oYVJUn8uLAOb/r/dhTkBx5seBAuQj/IihpavYSihDJ3AAj957UVRIoJyzbMSPcPB0dMC
JaseUWkUQV131DtY4kZjKZtfSIdkW3uSiQDwQliGhw54Z8RDVtp24IA8BBETn27YbuX8Y2JNJtBd
fUaYNxdTcuVUqgTF9enJWVRT3LeGqCIsk5uyrAI597aIByOecTYIb9XH0Sj6JNtqZJHsDR+cCeOE
GUSa3EdIhfcBqxbp4p0fSutLQe3p0426vz2Rusgr/6dELaECsZGRxtTZ5GykjrIsnDjOcacnfwSS
X8F+q/v48ZHDTooH/lPezifnOxhiuP2RRyW420WtnlCxunndDd0sF/RW4sP5VADJl86pBNUo6vev
yt0iHFSjdJcg28ewmmXrcQbgDzm6PJkyi5zsOVwIPtPwc3RQ5TylwtaTqwiF+YeNY9/qw2QsYm4z
dEKsqlaeNLja7/zHeslGsEaNq4bH2MsUiUilJHw6fgN+TdH/yLrFShWkpQV4x5myMjKzXo91Bg8b
+cCJiBXAk3raPYlCumI1JBLXvZefMn465bYW2OXR03anD9Xc3aJh/sbe2mXS/R/NmBIvQkyId4Ba
9dKuQWlsoyRWHTRrEKnhWRGcD6ua6Ojq66C2YdsF3iRSeqABfZv87jHVCUefiPJZxgL9nYgyxe1L
nCpmtjmSEf5xvIcFkrLr/MrbVf6mRG1ww1u+FkHvMvYjaAP4kEoHBZMPbMpLk2zSCoiAlSrky81a
yXExQDHjxiz95CythWGYAzp0WCxQiDfwWnK3xuEqlWYs9p8wxHnGGewyN+dOmn4RLPiUNEYtJC6Q
xIot92rr+/Z508L3juMYiR7Lsb+6Ez3rJSPyA8DXZWTcY48fyQg8c4j3WjBcSSkiRT9z+E5fiPqb
QIOzI6ZeRPopd9MosZMv13oCuTh9xIQxLjR9IPprk4vpvZ2qcwBbB9omuny492nCEQA8smQQB1vO
q92d6ejWtci6Zb7/SbNY1KQQgsfqan/G9LSM91GnouoF35Z5+fJEmh7F65VjIUlaxlzBOrX/Qd0W
DDzPXhNNhojCeW+KeHwcWykmxJ8drc24taZobe5RTLQ0GY/fVB17TuTRF62W6A5Vx8G95UtrAR+f
VsPTWZghvSCc/j/jwBDOO7Mi2RHe8LrLxHWq/px7XQ2DUYKfdi71rA9EScdXHAHc0APwZYzZOhLz
JEGYD3TW6x2i82BljIsp5rSeTKZzMw/EhK052bBZcI3rYG1jgZJvV5bbEqKL4T0UKeZSFU+LiT59
V8J3Tn2vghWQLbeC5Dm4YBSd4CEzT2CAr/Yb16Aem+hPf+kUca6Bnf5KQCgUDusI+nTcBDsriljX
+xBZys5vvyLJWojOlO0TtM/4lSEn+lwPwe+cNFsf2Mgta8BhZo57i13WYgma7fa6/FfJOu8AXe0+
haL+HO8DdJnM0qQEWPPiERMNqgk08Uj0hM5jIIPBv6lyxgSCtrOeA4QlmfDy79SXsf0eXXliS1Zs
EKYZZHn+eZRiLmEHthFxvks6Yk3aWa5PJHVd7STx/8lJLnmthq4ZP/rnurdI0IbUsyZnEf8h4xSL
ZOgOUyLPLc2Ea031mqlt5+0oNYwzJ29LGsHk471D3dmT42bDIhOe1d3dQVO7AnO4/sjkPswvQNfl
Mvnbd54GCQiKbxH5jz7wlibz4UBv5gt5+gL0Bs27RdLdmKSk1ebSRUI1P5ky8vul6O1oEcIcFEaR
b4lDFODNwE2RKbXL4ocgntFrkt5o3Sg5q2mb1lIjCLuiU/u22FGkw6xWz4tvJAKZn4aqUZtPOc1K
2onRlOnAmeBywt2WB5SmBn4krOejxCdX1uz/VB4ox9rfTwPDnj8MZzhr+wb4ftqUULw0duyRTlxh
wpGa/T4EMXG0dBsVThq0ihzEnB9+tfwDGlRDzrqxenKtQWWUP6quqNTKJni5ezyVmzZwrHzu793j
aP8qJcs0n0/CN5FYTPXZQmM0QHKJCY96ybYhPPeZ9veFRWBeoycTu1KSjf4jKK8PTVfBA/IZege2
E2IvekiLjR2mEtLW7R+XpYo1/iQz9syTKVYRYhjCXVUd/wfk5GykUTeud6BTdm+2Ln+0U7Iq7Sji
RGMNp/aRCPgOkUqwpI4LpFaZlGEJV07j4sby0mzm1Ueun5UJMw0TgTnvWyodj4+lotNzVSqm2G4D
J8k3cmyJtDMn6I5qrm/DGVP3OMZUThGizcKbAAnAO8fPAWeqz7BvFf/M3m8LBxckyiMZihJedq3G
xGnNbVppvuc4LlGMksFIB15kgbwTwRdwjIf4wZOW334/mXJsiF4e3iDPsYe1BlQo/JvsRbWi/6p6
cZ14bG5+f79ij0m81mQ+itPzW5iCTZl1x796nxSWzEkcEDUwc2K4/uQXwALfkI6EZyxKKfzrAMl4
vnQSTpBim76DtbaZLPSUalOD1iiCf85Pt1HT1X2aG2tv1RcaURaZPPsVB2w/wTuX+enHSWhtRvxS
mVgMrkqEATCkm46VYvRFccHwCd5ylaUcHCovZ2zp7BuZ0uUX8y8BGCyHfqgtGbXINOwrzpPq2YCh
rDZ3N767rJ21LAxeQTBY9tCsfffG5uCsSJpSukyHVFWcYwLEZYsVL1SNrvd4PD4zKZAmtZe0zYtE
sbvOnim4jz1BRpawqKZ6Wty4/agFdYsOYIvI/ib0d7P41m72zVA4BzFAp+Zv1TilX0/mQFH5Yc6a
ZD9VloyM4aW4ktzErE4uQKl/676arXRC0jtefxtWbn+4Exre58jqVvEh8i1dY6uP+YlCuNNExK2G
rO7mtiam1qS30TLsbNuTyiFurQL2AhsKY8n1KIdlaY2u8OnbUX8hYPEG1dsazipQ1T/RiXJCR62O
8QEt8rGNrwaB47PuYbchDvxvZ3Qd9Y1+xoF+80jVboGdLB48HyVtxRgBiSWfaEzHRQOtLHwikAVX
OPiD3Fyj+UxiD4YMHzKZTTx5UWw+hmPXadppY3tPDBvHkKZYFeEq9/PowjDoCC4BOy0PEPdP8Qtw
Nf40Vk0PtG5fsib7Z/FNC/Qz2dkGFkFD8suPlVJNt59bPn2cJwUPSkMXAJf+MkOLN8Lqdxl6bfuC
7P7Un2rGoNL+PCnGQnr8mPGximBK1J8KbmmcH1XSxXI1yQcHrAsv7ED0XGTGRbMXsZn2gqqFD3s9
Tv1ExPqofrJrPPXUWpzfnRAFut1dgw0PWpPks1CET0dZ0WscAj4jZZnMOt1b3/j7pvVoz29vAvHA
DqlyrEKC3SvN52FKvGvkhdMyO4FAoHQA46I72EFm/LmeT3D5jvBNPPtz/0k9HxOLjzgAq9b1wQcd
iwEiNPeTPS29HzxHKYQBrKm9lp9sMBUFlIyt02uk4xojArO0GukYsnP4e+1zU1SikqJF1I2GKgWn
If8KyMlifzjbH+PsydEvxfQz5F1wvFb8sjI1IFfwvUUWVKPkntTL440CuZldMmeooyxnfwld/KM8
A0dCPQl0oIzep3iwHtZts5T5uNdh+++l9CanebEn6SVkUqoov2F2wf8fDwQ4jJ1xyIS/Zkw5XeQf
WaJzXwN/I62hfHjw1ZHBasWUPYgRYrM0sWtlRvHhbkzXBGZfw1M+nhtxA0WbwXTZYbXzF7vyPTJ/
bjSV4Ryyt0RR8tYddbk2/AL4qHzcU0cEEWv02cZT8uKJbkQk6/zuJPr1TLSCIT8IxBEuH7IeEuXZ
DJw4p/Y9zaaNQ6zCeDzWhU8h2xGlLBJYsh92K9oQ7cp638aDc1id8ss0VFOLmNW6AoGlCw2NLGkz
+EtFbKwOe4H24LpjMXt38x7dlfRWBx4e2H4FXduMdd4Ih20BmdNrmpC9YT/qQqzcdwDeK/B0ZJsU
xu5msyCLr96Pw98i+EVfHIk10Fwb5SE1ox9aeo1xcZaYJURDlk77UvXvuTgbtE+NkAovqR71HUnx
WkTdlJiBqGPkGE8R+Lk1KPYtj8Oy5KUKr+0pIcQnKHF/kZeBxpkbbQgJyIKtrtcISutSLz6ptK48
Q5D5Rh00S8/CYnm5PWKpk2ilmG+hqU0qckiSYJwNDPdbt7U/nXXvp+1YX3fkNjeC+IQwYxeRCeoi
nMBc6tZNEARUcCTNFGeg1fVFEhii/vl8G8mzf183NhnXx7OyWMfDWMsj2S05TMXuCrFFHSCRkP2H
RSmyWzk26V9FmzSjSnkFGCco7IIsuzjGvxTYvnF9+ClqB+EHFtujUYI01dVm7H0Eo8WQIApvEZb0
/p+RnJMgixO+z4LnZQhHhUWqAmJhgs5X1pU0n/1bkvuhRjlwk3I3g2haFqPHSjkziFCnD6goEYUS
CnfWKpWJ3WyyU+m/YFrLfiVFrVNjlslrh4At/l/92ApO6L4hoUGmiyb4LccQTWpXFfgWAXgxWbkO
vmqvDlHv4dbVZqsf390IIxQaPhVgxGy3dY1jsOdE5rwvSz24SREJRfCY7YOp/QI6+0DYBH+qs3qx
Mw4V0gfYnUspZL1Pi1peWLaw3b8L0YnxOBXBU1NCH8Ue3gfUEyyv1NXzw3htfI9ZpaXybjFBw3Jj
kdHXrT+m6/rk+1ccQZ+NdAyiNQf2JAdDVHgyZ2BIrNGmtfBLsWBiMCC/cbS3xWb/T3MrXokikjKB
fAapO+ELqxjjEns4u2YawLlFWirPG++VUpc2v9pm26RGoifIY+jw/UO9Q6T1HU+pVoJ7Z7ocEekh
9JNjfjhHQaxcsyRxdsCvaeSd2DqPwy4+O9ztjm3J4eAi7PHRW+ENhdzFVMwna//fUq5SSs+7b+tZ
xRaH8LiJVnfHbjKB0O2rfw22FlR4Hg1sKQ4+u6LEY9/ITeLAMO3aTiOPs5YWsSgc5ITn09QQSNXU
L1rPlNVN3n6eilF25QZhxNUd/QBeVmH/TfLkv5CVeHao6ytTNNomcWcnlAP2QRFuoqa3I7qppTUj
sGmxW2WArQs+E2ccvi6BWG48FGwAEnYGPuUzx6lFwGhEHRe2sd7CtHbmUixHXgg88E6c0SostHn0
gIWDiTG7Z/tZPUYC4JIkldTAJ9XLbJnHsh4apqJqv7IfnVPSxFAjlbsWBg0o9Wg4fF9jZPIJ3zGq
zsy30NEgJCuonH+nVU1sEXwriy9H1ER1kmtag1ZdM58tjKaz31/OXhMk14QsYVmlNbwa9PefULIf
LJw1xlBn4p+L9mLeKlVC9MtRzGuI8jwOwuTXF7MvPKZGPorHrmJh3wNQ+EMp5+jxGj0D3iauacib
b/UMQq6+cmVJmeG5y+SL0hB3PtaCROn5/OCFuq+QTLXhX8K7hx/lMvWAPMTmsb9XehJgy6cYjz5Y
IXLcosa0GvMlutax4rfOq87zamxZX8r0Du5CFHXC6fb1qxXe2oNn1VGknfsrFSvRRo8iPNUjPaFL
pvpb+wM44gOeUKxL9Tra+Bx1rUKbijQj0VpPPv2yLhF7qrynN/jx12dFkvOlDCrLMR7O4OITqFme
pZ1KKsddjr63K+uOacCyQvDGIN5LH8NKHZgq0wA2yw4CN50lhp0KA3cxuyFt63ZzXVYHliJYOhK5
urM4rn/RUxGg7hPaIdubj2kPGsmTK5Qo36NV48ABZB09WLFuqW0FSb85PTPHACpb9LjI/eNNM/1z
TrS9lE56agC0jKopoS2Uudr0NRpmOLFfQb4n+1bw+CXSAN9wNTQBP5+x2E2swY6kUD3sxGMvJkRp
2k9wmKo/iKAMzjOv2P37I8BrHTEWhvCOb7twJawQWCng1k5umLTqfrrWVHc7F4Qe4oc9+OKRkh8I
FeZCPwVvEAvSjZul8jldnvycA9GeTzBJWO3XuNWPGHfS1WwHzCBpFltTDjfogbTwZlwo+pKY3BQM
26dHqHL0U9bTnTC8vnMMbpwS72rHY7wANBGegYpxC3BfNCgvsIM4atGwnClyKXRkMHutc94whwZd
gpO6oKrl25AiHE7VlUpPNdEFzAu9DmkHa4gTP+WxdjK0nF3S7dwIYx4ibPLSrP6x752lF4mJKJbJ
NlBECdU4xRNu9DlG0/hjuYSHml3eLAc406wp9QQZ/Rt6fzT6S2rlPMUcKWEnMJaW4SPaiFSogjbo
FhIm9kBQAyM8Qch2bJRDvbBqMhZonhE/VwQp3FnHnbe381ACwgjsrIiC4va5sr9tZiYBLkoxU2J5
EPDjhcC6ukXtJOlc3Yzwf5XOiCVupWjWnjcH+CEJvgUNjfGY5VcbQEZytnBnDb87ecYWirZkkllk
GVO+MF3OQIC3YYOIC/8KJfdc7mtijgK/XJz2rmCQBba+ryBWUiaPQMsHa8Vb1QxV/SyDGqhZii8V
iPfUa1QTkBB1hthZZsC2gSxjXHoWT1fkqSVM2Z3sKIgNyPIwOyUOgh4I94KRKW4TYCSSq6YeHCCC
0hSABWFV7+YZw31ps2EZGr81nSd5fXpcy89CMgfdqcdZhtPK5PhMpr4C0RbEzitxccwinEKqG92+
zGjkB+CksJc6ciZ6Fgnhg9SJnJ5EMPCGvmVQhHl0GsqKNbZWBit7Z/s5DGiLzxcZL41OA71huCz3
DdE5WSpX0rvdKCbtAYq2KOjQgjvjeHkN38bS0ux1xy9k2aXY4YIF7vzqgQ+RgTM65cNUyB4H+K0n
+gAvrz2TPzI1Ri/Ep/B1M05D5mrIieXj7eMqnkk5vZwUsfjRikQEud2DajNZXLqauBZ8UHR0vcT/
w49Hmvvi7qcafGAbZexOGwtnAnNEoPysJF9zJrYQKMHXeV0/7BFun9Oe5GR0e//oeTshOQtgW8Vz
MMc7zQXUQqurDbYnMaTJK+EpHbaZ/TkeCBES2szxe+jkcyt3mtO7qV8BLIR8fBfIJscgroz4h9C2
rDOe/Y4mYHiei8cZVaWh9wOOFYvHnvUYiMXS2y/gabAZlvpOO0Y3p78bz/U/JcdP9qkNOcd00RSJ
n19V9hsZjKnu23Igx4VpC+dC1qOskrTYWlc+LirasJEQq6tRME6lg5PX4j2licBbxjfomBKa0MwQ
vSDFaVHasTitYvSQ0wku10sJjqat+Gz6WV6HO3wTvVETr+VkWo/9Z05O4O+WFyFE/Wbg0uotCNt9
y61K5qgbbDFK0mfIs9Yu+jY54GOrDirc0W7gHB/M0D460VdS98iy0iWPOx7fHsODkYft2cl9FJmG
haQb7lzlMK4oRYeKM7YaVftw3EeAS/mmsOJXNuAidf40igNzVZdogno/Sl+nk8L5ii8XXOt6X+WA
l6FJSHggtjKmKLJMuk9d7rEraIM1aQg4r9Q0eKCxkHF/syKpI99oEUuDXoRZZBxNslgZEzfXs0hb
bQThQe3qS22RyMB/W7BCG5Y5H3/wmNlfadWL/NTTnmEElMItCcCX/LZaZhEuCESb3GJ+7TN2a0ZB
h0uh4O7aunZ979OfM405oqypu0FNpjXx7jzJqxunOyo4rYjoBlg9jE/YoAIiM08TRvVfvZD0xaJZ
uw/EXrXGZTcxgOuLE/Zm8v4r9+CbjyLgcQp9xKXvsaJoA+rn6IFLiug2E7UtqaZ33lblm2LgK4yB
8BPhXzyMA9lEK+nErXYns8v631LI7mzqrn0tO982BcmlC/b5LIEo9z/zVMMjo3K6Y1nXrsV/UAtd
A9XbnVpjNtUMj70wLixPw76lQoTKRYVboENTUV7yNpa6pBwDUN0YAJmzk4B5Yq/20R24TB7TLOvX
Ow4C3QmGbwEYkNWIlvvff7ZkyplFyDnSohaCtG9AuVO+J4QcR91TlrVtVZjgseegWSv+QwJB+0I0
tGEqYf7IwkY22IlqSxDfg3EssUlFhq8R5NRuN4gjZTY9PIpN/6hjaBBu7R5bRE94ipf0yLoaVVF2
qvbk3OmJ5zFnhmKWwpOPsBfdSDCS7fCFmEEQr/0WnV5Mfltcs7+qEaggiJzlyrE/YZWkpY1//5mK
BfIPkEVc/u/5JVkeN4w/udmDfOLs9h+yTHTpKlcUpWIs5UfKzsAkzNknfl8zhz2ImUVdpxElMEHV
gzvAEt4W2fy3dYbMEugbAI0/pvX7gC15k5okt2AQAm9MEG2MaC8IzoW+7EVSgF3cViQXSMSbx/Rb
YbTBgd/Thsx0+kCeF9G5RUOE+W7ggBJorlra4xXJOGpmG5IfAa0SZNsw+lri0ZvupObWMMrljR0V
IUsSeCF8QJ8xsVcdL0rc3JmfYtNomFbhE0qjxhBfHlyXSwg1WGfGJlxZTx3hHtA59M3Ii8ylpQS2
js2FL0DFJrXICg92/tcSM2Q8TttO1TgpqLdnXmJ1oDMwL8GE//8ZWkTejPNSegacyum6JEXBTns3
NViGYqBWJEOjDsf75kZCr801xOsU1XjAPr9uNqMxInLSiPuoFo6G25ko2ebPkIiw77v8C21crJRu
F+3350Wt60y/f97zrxjol4j7SfKoa9c7Y2zK/UZQX6xvavfWuA/YzfN2vpouODGPjbauohDYCVYn
munBGNx43wcWCFYzkOtouuBb9IuEAJoh0zPQlNYzcZrtqePQnCZkj3oQWOmC7kmc3iZj96rxuKe5
+yTi5tiTXt6lDpa1kDhR0o47ohFZY2M6rrgIUWnDYnA7o6TwjenhFqu+olXi+jEwacob4reUSGRJ
f+9S0/VY27ohNUDoPmUY7MhEfK+rKDGSTytAFGJdiACYn7A3CqGTI2mCax0kCpanbTsrH7vr/uD6
m01xdZ1VKfWjzAJXe7c9FWsFlpGOqWfLucR7xSpuSQkdM4tjJYCPQxTNs4JLuPUYO8+gEOhsP6/K
w1MB4wttDKARmaNPcwjr7lBL+Q768gsP6ypt8hsxazJEQgay38LHLWjVDp1Yhw4ojeLtI5COLNj+
2ufXAdsMbbQR+bnwX+Zb17dRFvXPI8ewSwCN3Mt8tX/QyJlhh0tkD03jLFuw2Z9ORyAhqAo0jBSP
9w/nNgZgmlDp5BhmhyCjjc6MFtfE1Ho539W9OImSlSUPReH2lXWQ84L09LdiR+7koaJqSgi1zWyQ
youpbMXRYZuG1It/XXV6ObQpu2mE3HDsHSyiomlbvw6BxsyKZdSy1/6gr+/AtriZSvfgsVJX119z
/4U7B7csAeaqKIEJvow6Zm+rba13o4I/mJjz+b4VsazgSnCCwruozZRREGe6Z73IulYrRgaAo2c7
dX837dHiLlnoeNktRAigr7NmYYGLOX9iQzHjVtRoXsY1efYQ9lojGDJ4z25Ki7xMJHV9wrvGuB4u
qdsKktahoyvg7W3gdnJSME1k4fQ+yxHRXsIkQylvYy1ZK8xMDk4k/Qna7OohtZwPEsZar2OxUlNN
pQNGHi5OGHAIL66A6SnT9Ps5nwXSED7ir0noVfsScXxZHWg9CV6R6bN9ge6kgFSRwjHgoJ0+nBmH
Lj2Lho9nRaq3XJF0F15iwAwCnZZ8tFOARNFsF66ylkCVZC7idW1cTDumoZOs6VGgXsYcDK6vTPgQ
zzSIW7i1g4APlnEaC4PpGOLnNKjUsI0OrKcVtL2PE/Vo35djrT04/VHpLuQlVqXahZuKj9EXn9iC
qoMBug6ibOBYKGlCEWKWKQxTa4Exx+m5SSGr6YpFO4amxRRI5StGVbg/q69i+aVfXgM5l13VCQkC
XOLKQvRMrUtuwSQlhpgar+CKioRYSBibjWE9QynFOtrg/61OCvANe9yxvosykeklfWmj6xsxAXeh
eLKUbMi/KJc3zhy7/0OQjqw/ncAwGWOcMZQ+NuzLW9XV4Xn/uHhWC8mk2zAwL3J+djkiX0KK9Yit
QFnVrK6CuJ/tOZtvbsNVOpHSZLYRv6thQR7sBxM5wFO/8hbqrigdw/QqV+1DgUnjRrSywe5mkP0F
Gj7EcAgTrPr/MLkQ11HTUj80+QnF1ww6/3Sm9B/MC+8ij+ij4nkCw2Kb0rksRJvwvXR3S3T1vjPh
W/VUgqOD4Fkw220nm3XvMk1gcs3+fl+4nlzKyLZftXXViJ9jTSDolf8ojd5l3M5pXJ+eWh5i3XJ1
D5PzKaq6sRTmWh2ezwOWtdmhtLNoMMapaehZbn3ZTBhSSxwg39OwADuidDleo2M6cKJA0Mezv0Hy
1ZSl3SQpzPpt8TraSX3LjPQHFixS6kL8iFvW7qx8JsQEISjAWpXlaYCLiQIT6pyQZLwe7LrH8hqA
VJkjSwxq9izeFmfEFWVbAluEAhtdsbpvw3iSbxmTyUXGwQrDtDmNs+iLAFvfUqsqZCRntl37nxf/
FL8oR8Es/xOUsR5ATfwKjBcJe2vPw2/ZHPm3hza2ezAkDbwH/mgXHhtZmiFpia68ZqrMguu4bMgp
K+np7BKy8WFgg2fTZ0dAOYHdA8HecBsfcz2Fg+uzuvwfleRKMUUnRiDTD7DHlT5L1pqe4sc5u8PG
J+4M95BlarIpRZizF+MV1CBGvpH18Fpid9YQS5dbbkV9eVQW2i2csxkPY7BPaYq4Jpldl5rTfz36
ICDtauu9wlU+jULOF+co9lWIWeYVCmzvD/9Qr2prCfqXFmdH1kaddB99s4U4RZKD2qeVLcb/ZB78
bNcHCq36NXp6xOVVFWwwruRr/4Px45xtOfadTF345Ir3BstlOVCLM+pwq0QbwNlUBisGtGC0+LSG
f4FuLrzR6rbyfiKfXBjJ+cLkYipkzaZc1LyMcyDKYXp5+Ow/BA8oghxl6pUkTT7+6YoAFWdUzn1X
+uXdzLV3AyB16fAWtCiInjSGxCrKeOBOVUQhfOo3IxrNyfHhs05MzEOqe+kcS471uH1WjCLswXRI
pE04ITvUHIxu9Up0bmryt4t/W7q3wEqp9kVZ+GPHcusl41KEEJz9RWOIptDvDkK8fII15/WJOWzs
E1Jkyzf3HHkTCVbm59o5XNnyS9e3yRdrfDXeRUcZFqPjdAIr3aCJmfsvy3+nzXUc+abS0qE+m+wJ
8isyxYaLRAnIhTcMfo0INq00xtpW7woePNx+fPGka3UXIzNA0QcR+5wJvs/s/1OYECfFE0c4ywGr
0dZaihuwvC/bucCRG5Jp5Z1R8AEvBjakMNUwWO8PcjlKhwBR4Bh/GoYm8PlaoPpioURZ5r4USRfQ
nTjubddlIo0rUZijD9dZi+syrFFetqn182+Xe4VrQHJnvc09LwwsxTudE40GTkbVf1fdozaIkIAJ
9IOxzr99jPh/mMvQYuXLEi1tXIFcJcQc5iAcvzIin0RG2CrGZvjaXLjHmHdpb6GVsUmck0m+/sbr
YOVaF+ug15JPJB545mUjOSvzSFElxfSlFSJTaj57SeCVZpyy7QpL+NHrHSlKitaDErltXzba1F4D
1UyxYOizMKlF58fIsaQBvK8omSvcmOUNXrp1po+ibNuGukjNhs6hbW8sut5sXGfZldZ9cZPHeyBQ
HwX5OJJySH0Fc5Ds1eeZcZKKajjM99zOKRIL0q5YTUMeGzYeBsqMhx6dOL7WixZRHQeYmiQa/Glt
v+UzVdYyBCM+IRJjPM7bDlEYnHx12JUakU4gdhwJ7fePS7jNq/Oxk+4kq4Pes2p5PXhSOrbl3bcH
SgLNCHMQYmHJfSYXIoIyJ2L9o99RZm9vQiCcW/rAgNlfwE0N2lXqapMGWLFObZDom/n0HcCc2gx0
PDQx0DDsho4POyP2Jf2G4gu1NHzKK8xQqPcUhIjFxIvZ+ikUPUpx345wM8fIvroFZHKGNw2Ryryw
l1uTDYesJybBCYg6Cto7fhIc/Hm2kN0IVtgniMMBpoWdlMfWNDvSymQRURhh7YxJTC2XgqHx4qCa
1vHXhYi8LN/8ok4m35NwMAMFkVfWckuf48jtMwMPZdm9FggUYN1f0DjoDo91FUBIo0X1J5YfUAb6
T8Z3d6KUdERphMirbK1goc8UkLMhfkUeC0ZEaAYKVEsjy5JnGk/eG+Y4oc/yojGeLxsce/AfI0oK
LPH0TmCCiJksz8zOhs9vclBCIdvw905DyUZcFoQfUQinxPn4UEjCt3UNoUsxMwbyxG8SloZpLy5g
hyNMtJvetX5FOXO2jrXRjNPMV+/PfsZm79i5AoXNNJpCa7GB27hMy1+tOGRNe+zOKxomr0eCwkjG
6DeRlNsT4V1FkGt66H2Fw9YSyGok5MFlJyMPY2J8KpQgOwugq7GGiSETfIthuQZANJRpcDkMOYeF
55AtBymeDh6rFOd1+na8AZamCMOdeJuxVpySHvcJCyzrBej5nN2ItytD8R2ByH9//k7ZYA4aLyZV
PRza35q2MauQIFgVMlz/iu/wl878LOzs0Yb2Ji66T5XhxxR37bmogl5f904+CDVUlr2Jxrya2AgR
g6eefMDr0ZPxWw8mOr7Y67YFt29hiC1dnMj1Y+WyPksxGwF2cbeiWnEaTwc9b95mgeVRwIzT+EbN
bBNYiFWSSTWjqHqEaGugL8wQqMp2FsWLPDgwoyBPZY6UBsDOWL26m4CBfBnaImY2HtlIrnHOe68/
QAoYX8UBfbxjULFunCk8TouryHhfkyaKg+OEhxrLvSEfBx1KmeUADAMa2yZHZUPITZ/rvZoHp0ne
Lj1uCskbT02yBOh3YLX6HrLmI0Vw6EeK9cymQHJpM7dQwGXjzfOVlsUHbzredmlKZM3unSmrxtFb
Q4+O6z1Uv/EvTN8rQmgM67lYUJ0vCqR/zQSA4la537Pu5z0xG2hBY7vhBxC1Ybcm+klGSepJ7ERa
Rs9YlVu9kWex7a3or0r4zkbGK7F6DX/BSbIZu4WnxXe2GKKuBMVykTPvkeQIpD9MLo7iIotuaUO9
RRCK7gQgbsT8xHmBh+HM/4sGUxOs/aULZITAQ54JuHB+uNo+0mQWULCdAKlon4RVQkhaMhoYCPcg
tEy/fPf8u0Zgu+lD2qO1iTuuKfRcfe80n/9tiTSNauoQmpS6Wq1qJDDiJ++UvaWcKKEEOb1n+Dqn
FFwBoE2KDNFbVzbZnSzh5EvEEorgTzgC71IC846w1cfgAL2y3Ky0XuimJzJrbqSpkdo8csWtwHE7
Rj1lTfqNaBszlPQtwetOwD7CWtupmmawZb6jItPryXB7o2XtNfyWABkYX4wbj38q+noYuojuRoD5
Zt8ceIz+UOw8RhTLLe1vi4rQVWnPdkpvGvrJTguxNwaMrLIhyu2K7kbyGuEsRWZmU+uemJ9I99rJ
QBMYCc0EQiIeZBq3p4MBi2lTK/w14GM4G1PPUTJ52yFm+tHm0XqsjyRnpJHo0z3ls0/bQ+b0Bcz5
Y74Eoe6sKL/UR1O4z5MfDP44OJbllQqILfbunE0gExU/nlVa9MUl+waDV2NmGH7Zeoe9Ep7kiTXA
3TrcciDH+tOv8c1AVt3Z2OKhySuBNlhxI45K8FLMcn1HTiEEmQjkSPLnch/0M50S25ChvGuX93fC
bqDD/QtVPk9w9//Uo7LRIXwrd497ahDsuYsFRK3b4qO5YNOlQobLiQ3fsfs+kHuc1yp8CpGgmzSl
OCgIRARWbbjt2CnfapR+GV6LXpQfcx1zfLtCWZSj0II9Yw0oxuJLaD8U0dGkTjp0SxQ9GwWvRGPo
tJP2NjkdeoQDQAiLYUZ3h7e7Rjw2zELUBbHwRdv3K+UBAyDwNG+AyeDiOepQGIDyp0M2Akc3lPKj
Nk6IG0dwMzcSSnGaZPUnPcL1qKeDzt6Ta4Ei/eA63X/UwqlenUy10/vKk7dTKNTFd5bXuTA1SVnt
Z+RjC9gfGcxKQzCa1NOptLz+u8dThbxjyN6K5am1F0GbQFBuZltaO26Y9rMgE4WUXhkicWSHHVmU
aelOCmvvfp05QkSENwFVgiLZ2cviyYsfvkjdr4jsrgWcbHtWxf81mXabo765rrvC9eZt789dxdWo
RJ2kvZoX4G9amKL8bWB2sob4Lezy3w3gGDGeTxsiRzJkUV+8APGnWGnf/wqkDCE3Ipb/nsne1McU
P9iO0WhxuiqJSmfHoddcPR5vAGqXXKivgMzQlForqOPyxZhoQHr2rk6Sh1/TaZiJkvmykn7YcXaz
qNL+R/OVIRm9hFNAMA5YKl14YXQCvX5yC6bYSw5/BDDW+MpredwZZ0f8Ay+Du4FhzeiMuN0uhGbn
xLo2ObhhZRhK70LVoiIXqmHVwPR6bIOCxhZf0Ae/+Fitg22JLJm1yg4JCLVaW79WdeQ6ogU32+dS
tlxwXJafbk4rEVsQF+WEjW3AideT9IWeD1jYM8wm8xSPjmI3Nl/wbfuQRz8JjqjoPYr1VT4tudla
81xNUSC/B4aXDv9zCbRnOrh1nayw54Q1V/6M6rlNHI88L6zrINdZTeeFgJvxIEdGpRsUB1YtJiF6
s9c7eFwomY7SAWhSoYDXaOtGQdXtufSSnNH/QYrNmxJxHZDsdz2tqkuHW7n994ekYtV5d1Mwmk5U
9MGXp3wXq0y8Aemh97dJvGGBvqfkMYJx8GtEHewtyiWvHe6LgFjzd+r5tguN4PnC8C4DB42bzJmd
9baVZCsbdv5Bw9Z1tAMcNwx2bZx90jPT71CviqwwjM2kHkVF5xmgEKHebbysgh+C210zxUQFX7A1
MY58pV02qCwJZ31dwTpU+8dmJ0apNzPS5OrpXYU3mZZt0KrFtU8SZZmg9KAYuomph9k+LvYd9vge
V+OTZZxPblPh2AXolC4flTIbmBfbS0kWYCeX6Pu5GmpIkd4eN4oFmCbmyfzA3ne00zHM6zSTsbja
7/Q5//oNyC17ATfNO1sQ2iV0EXolayZEKC8xfTIMW8dnl2WNErrZv9UYuYbhuesKtnj8bQzQ0tdy
YS2ERN5FpUlVl4Uwwc6AzdWpuUGi/IK8Z7OfZzOKXX3whinhXqeN/Nvb/GBLoWUSIfky5RqsijFo
vK/ND30/olaKE9d4PRUAQuDymoYYa1y4xctWrVl9POAJ7/OZ8prTdL+GwyT9K4JI0XTsFNeOCQo/
gYYXGKdhdCt3+4UYPpmCKKBxjQZiXT8Nw6faR3QRYuTGGZAZWHxr1u8fvB2UG4ooNvI4mlnDgbqr
R04Wy8BRpxk3J7OvQqXOMDVQBmUXhihj3IdWbSSQsfCb5a64CyYLWXie/cm0BN6IJc6K3lELhtcQ
ln3td8je88EOfDfQvB9/CpetoTEXaqusgGNGm9u/WJUOxhDodIUdJJTvQS6PpOc5KmdUSErLnx1F
W13UKcQbX3Llvog+XBOBTmVQRXGgeQuHPbVs3C7PTwXD3/xEwB/gGaqe6CgOABDfoB8hS7tV3t6t
hCvb8grKdpKt8Dscw+WRQrclQX9iDy8GRV/e25Vx7Tfq6jJm6FiFO12EXHgYp52sarHqeEM5Doit
b4Eo11HtjerlXXguPL1Ixo4Gj6cPFLh1u/WXWsawcSVGZX1Rn2jix7TyhnLykzdA36vrVlsaHlyL
x4On6Mz/npHjqFGfApbuX45o6K/sKAphYP95/VAmP8f5Jauod/GV1JQ8nb3zg/9ndn1Dt9fc0DNX
CcvAs/xPbTIcWZYQa2MejxbHi/fe8tU+cBJFAaUbzvnfyTj520/I20dN39FZtkakLwmFUoE9B3FN
zRqvvI3sZcRPpJ0h9LN+yvyXM4Sl7CMCdJdNWRZap6NK06efgUbIyMR4UTi4mqQ1NC82H6JbL5wo
a7qKATof7y6EDmfd2811dZbFJgsjtM89mJ648405eZdQt7N9tznrAGSStue+dPrsexR6ps+yn9Tn
6wzx/pA7AxEf3EhaXpOVT8e+kH55+EsGKfEabgwgfVBTffg9QKImtTmWas7cGlPp4xY/lBpKIfcP
+t8/G5+AWS5JlgjqINR7yG+8JBkrIvdd6MxwInBNu/WBUixEkqgFfzqbwIzwYeRGzPlb30Evncuw
V2Gy4HkJoDpLUWAlhQMWSgb4AJxQu8vTzpsqZMYYHoVuyWLn1NOvv5YMQm10fiRU9IYTGmhY8AIE
aAnJ1OBq3V9tVqMBl2M6QfD61OXu0Aa27cQwfhUC8lHiNcHdhTikwRyt9W7XobzRgjO+MIukPhi9
8NSGxCb6g+RV/F9N2HH6Il1cvxuPQCFBZRTgAXiVHH5QsOX1WZtBNZrgZJxI+fBCCIlEvWPAw3ho
s4xA5V5bAz/eFuWf7mJW1u+Td7q4tdR+YhoMpTgYUHQfrts+6UZ3TnKHOzc323XjMFL4BLu+Iw+2
fvPMeH0ZWEJumoOsfNX4LS/Y4fX7lw4gejowJiUlTTwbIrx7NzpC2gzPetYBw3+YcDwJPeRJZS91
zrbuP2xJ905OS/JJupt+/1gJd0IAshdS0kd2H3ma8q9BB3ZYdT+/ycQgjOvAOmH5uM8ZgjlQlw1q
NqjbHE9PpiP1/zOLKhEswE8pYq7f9PMtWHqCSXcvEkKG2kOPF/17VR2b/QY9KEw/RQJGr1rh8qqp
54Jc1BAC7Dcqgs0IJ9oksaPeZbjkXRR2jfB+JwVbym56zo/h1bk31rGjrNM1+JoQLzsWIMC0tPkZ
8N7vAcngLLOCe1U4ds/Tqisn8+WnCXicIf3ptqCDI+Xrd2QtXK5IWKOu34GowX0uv7vHYWTVnlTX
QAWNeDmMNTwROeaWAgRNlrV9Wjr9Nq0xUSZGkxr6BJw6+FmjViKCo7cGLgSd6yvATfPz1I060bIM
Kmze6K8Fl47d5TOfUj09AkNkbliHjkN97rCn0FKDcR92Jpz5rvCwmFnl7mHY6Q3jldUnixFBOes5
f/5CV1hutHpg6CzWVwsA+7bZnabsK/EaBF201eS86Iw8Jacf9M4KFgp/WVXR4vrEJ+etDF11nSyl
FHoXu7FVot683QK/KPhmPi297iSHdDrunt4W06aGZUyoAxts2GPznAJQLX7q7DkhtbBfeY+HcMix
loEPCxuKf3Pc2mK24HJbsqRNAEhBaPSrj2BQW9W/w9y+4lCKuzsT1ajGaU1/ZPppQVST46VFaNKV
6lR/yzuBSO+v4lTnF9Hug6x3FuOlPzP+w6++fFwNHc518cS26JOoMwEC/chTZpDgupKOvWTiGgeX
KXyO2x3n3XK6td3tP6HaGtUm0xDtJsfzgW0DkgM41XEMocio7aSc+8b8xO5hLBGSbPQKmkSjkvns
cHTldJ6IAn2apNgmNEAF5UEoEHmKrn3MU6Vh4ctJ4DSyEgaowzfylgRhOAMX5u1ufw9bTnNeI5+U
sChiip29qDCgglmSA/ThBB+8xKfUvaSAlVpK/Nllmx8l6wNswYr6WOvg6A2B2Wzq8ZLbzoJS+YzR
FVgMkeoyGheYEETVBYeedTeBAQNyovIv7TUGOqIP7zP/btg3QihbGJAxwQgwBRsL9C078E44tAsx
RW/WBDiAHpLa9i5ln3SdYFzLUFxEY+ro2O6jY2KFs3AH0+rHjIh6e6A2b6KGxZUAiGBINXJaoXJC
e06i5cDPvD4UaTMdK1lJOnINlzrMmQ5vK1BCjqYsJSh9R3f+QhSajqy2/FUBHT1/ui8436X+UBhR
Y0BfU9C/RozOhIUHEUFtkMNS86ZlKleGIl9JYjfC61Tsyo+VUyszlcEpjy40QB4JbK9Y8f8I2+S6
p94jeWZr/WQEe8K78wPZT1p1esk2n6I9muejprK2hTJrRV1+ldiTyBnmqeFDyBRTbGvgPytwxqEQ
nAa+gQbp8iRZidRKxBm78LHY8xAeDEcCXoXirzgygwzHi06JzHHUlzFTpYjXEh1s0DTdOj9gr5bA
YBSOIfTeyjOUBd9VRWIdOBEvMRftX1qnrmUc1+qDL3dd/1uN3z0u6l2JhFOM9jBud/ECFYeZUzdd
/kOffuDa7oQu/rRMlHLUGcM0GJfCOGNjBIuJ/AOtMzPy15tQA9XvLAIyfQ1MuLxaXVl2m3uPlKPt
qly1tuFawkLMp82SVgIusDudoPBGPpFxDJD8yMSRH7h+Hc4ZKMVk5n9WDapAL7svCH4phrWm2qLx
zzgIk7GqZ/NJsld7XOGi7U15FQCzZMmqTMyFygdVFCwUrnNd4Ot+nk+iAKJpl4DBI8gZ0qWjxSxp
6rfniJfqkeCNRzdqGrcO4rDkTtoI3xa5txSLqW+JmZr5ehc9yddND2/q4ofnGcEucIkSdAkLCOqh
3yd1f1ynBONcwmEnK+y8R2RPxVAcFMFd3tgCUMDMR8X1BHZJGNshoxt88/18b4KycCcDNe2xw8Cm
73H7zgGwkR7cR56s1HGn+wdTaU9+c89Ri3esTyV5YoLMbwWafe7TlzQau56KYH1yK+arxeW4IS26
OBPdz5I9x6MJnRZUb3rJXPYJRiEoZwK3OemTBcFhYKgpDK9CeCn5LZQzzZjNpCyMi43/JQvnfjlV
XoASw3BrDU2xnsDxRyDVvUNXrMcNdmx7bBHG69Dcv3g18HCkJuuWs4seOFO+BDbWJS0Pg/Hr99U6
5sULR8a2jYls0NdxgN4QQVVUDi1OplBFbFPSdm7zLYJAXB7OIvXHWnmai19tr0YN4Yoz2KrvBvIn
ZMkoaggLYf5Jx4+tvGmOa7NIr4RzrESZNang1Ne/Xx70Rx1q9Mto85NMWfcnsNbXYtV9QjI+ohC2
sjahh6ADlx5ACLR/Mk8VD9qcS41JqkS/To5fbbcREMNqdf7EWuKT9NRcbBVUfnmTaIvhTppq+oR6
Ivg/SXVwAAw6asZIOgvHztz0ZL34TDDYc9+SDVeQdLU6WmW0ctpdVDQvaLN8/LqjXXPjHkvyze3V
rnFd8POmfEP5/yuSPmzp8E+UgwH77GBQdTrFXVi7j0+wC4Cz3e7pB5MnzM+ENxjLqTMMOSjbEr6V
j6SSRIv4h+djqFZwi4b77hnDDU8uulKtAb97JuIbxYn3mWpPwqDWycLZyFe36t3d9sG5Lrv7UyDZ
DQVN5YV3TGBhvkLsS37hlJtBarBfoj8K/XNEqFmK+PZsNKQP2GKT40fsDTZ0G4FYRYvW/BeaO8rE
6RiVXGY9oNYcyQO8AD/FAi4Y+Ho2jNoFiNHLF+M8cLDGI/MxtUW7bRhtD/cVZt5BUcOyc1wi8WPe
BYK5R0HH0nQIkuIAVb0BTCtbJj6r+ujqvhjFQa2j9tVOYWLXq3qtcNjD4hlUrxhRDlpWXHOA3OfP
3hhV0bOAPFrfR2hLD2CfEXssKoITSa4v2pASro3XIp4tuG481KanL37420HZGuLoReiGw2DZrKNs
UhZCTrade+dSVg7/NwGnLYDDvRWeCpxm+6058FO9WHWH+CTYZMEzXGBDc2jhDTzR6tVY4wJlYTTM
/IrZ21vfA4Wd73H5l6hQg9WvvvPMRluoIRBuFTbUIC9/Ze0BLvA5W3bCJ7xGqQwee0eJkDDWc1j8
k6O8MhRf0vvOsRMNT+TAU7qTUJN1X85T6dkCyOHD9Ia5W3AcIVgLFnlOBzbZbXLsQtj5zP9gEDU4
o5mATkgqhMSOzvXWjmEJGYJ1TSPdgvRbodwLk53s4ix4O6W18fUrOLitIKUNpU4VbonGlSFdvma1
hEDndKajVmq72X2bwn9XUhXrUBqG6Eedx3J2F1ZkvimfqH6eQES0C9Yde9dNwFcCT7CrhGS57QPT
nXOOPM/FXgr22fU8hBu1e3I5kGLREnYQ9bA0ZC4H3ZfUBu2PVV4Xl1xgjiszG6UZ5BFH4pFGU9hC
P23uhon7uxvNRGCYwgyVMMGZt0eIQWIXafZ0A7uqyVeigmDrgj2I72QOLNWZ52B3EBEkvUXwU7hs
l6BrxLevPq9bxG6EZ1PfXcP8hALo79j90lkjpa7xDZuILpVGP7a3Zk0LUU5ahir8PbJ8Lt+1U+/F
wno4YOX1OuG06KXxBYXl2ci0T2flwVJsHJ4gDUOaIr3/lrMuMkSY8oPkkcpZoxoQToc70EBekB4+
qD5nNvJbELAORmIqLmt7hYWqJ1GSMMS4HVDuaHwgKZLdeHEP/1n9owyRsvpSprhk//BYCBVxI8VU
MoEFRp4Ve9cEu0dvXT32uVPHu3dRmKBFOz3BFJgT35APVl7fWsZmYkrYrKie7xKMP4bwEuEi+Gzx
PB+K7QACgSlT8kf5ERnoem94rXpdOmJ0zhaElqLIpVnOuL/pXskt+A7F0YaMitHdXvIqCfZ0lnxG
G/zznhS3SRplJxlC9PZB58MrR8AIrFwEZVeVWWax/95Zjc+tuUyf7/VU3105g9tTdb+S4CNuyZPJ
e86weh1CTiVWmW+5DY9VRjYA5bHsIEfPhBLwkMbCnmaalNuTOzCieK9HhD/9Nrzp9WSuxM9ZI6+G
VWOCFZtl7+KqutVnt+9KX45TIEX6fsETUPhG5SO9hMbyK6E+FLN7YYkzpKZpumioQdip2RlC/nPL
XEq7w0AfrkgqaPhmHu/WhMkQQAGXwmgFNv6XlH+S7kfUb7FASTvT/jniTV1ZRInB0TQ9s96vE/pW
tiQEaTNqF+StlnqkUMITelZOC4BS6oTTd1kZ6i7u35SlVSWWW9w+9VoJ73HjI5WlmbowPvXQKk+g
7WXAOnjLA2XI+aOGEFBo7I4O3XR3Q0gLX87+jecbDKLWGcP15bWSa5CUHmY1HlCFORbi5YrgPWDS
fNHZH1dJt/5aBgBW2lhwGPb0LziMsLRgQfcSY7CuCBO0prssP9pOdlS0HwQIPm/yysqaRLbinFQX
+MA96A9hDd1RoHZ6Xuti4G8+UI/VBbe7XDXg0me1LPn1P76FLOPk8+Je36Dj8bx4Lk8m8C+qJLBV
L9aQaAWE69LupJVPnUCKqTYvEtSdaCDkurZ4rGZQ4ajc3qlU03+m/RcN0h2gMGPARtSClGin90Pb
w0Vphdi6dQc1Ge9pbK3BTeiMl51nYSpmvoBf1q7pQfCXi1F25g5in8vfWda6QtDVLBOdJZ0WaJzw
0OEZEvvMF/NnNfSViDW/WrdWcRswj6229zAzslVXE35lbwvUzAJ6XEllognX37g1Gl9Z5hzYuyyJ
0saChVfiHGFFLh6a/Z442nUP60jX7O2K3GC0rsadbU01xjBg2T35daAn6C4Y6nhXTykDqCeqg6WX
+vr+8PLWKPDvV46kFhiIYyIgmlrAkgU7+cNcoQAcHuLd5ZPJrJP+pFkwEWvBNcmRQqXIOMuGIeE4
lo9vngFvOnKw6hMKr/VYQXANUyHVFI/1XsY8V5r5POZk3CfdBOLFjUsCJWT8VUBuyMvT6NZVV75J
3EOeTXQ2ObRbO2LnLDY6E4CbAOk6ehKvuZC3uUJV9CSB8AnxRGIpub1XmOFGQXcp/1VnBbDl6sgt
5drGYS0n3Rau+kXGQ2aQab1+Gaqme5QqHrvFR1eCusk1u/+JFjjimHcLaiuDMyHyuWgi3j4eqbUr
u1aW8tbXxMH0Riw/vmTQrR/E3tOA08hqWwtGUt4InYlmZJ0/LlDMDqfCL4nRqALzDR5c5forunzJ
7lThcArbJvFiXOZGxMqzk/T2j9TrmTgBJ1X/wPLrA3VslslFIvXats478MEBoQ95Rs/wJNnbyZTd
miV5bux23oiIzlgheqRrhmUNdy5MgySWkCK/JoM84gfdcGrjUdyasNRvIp359qzz5V6uNDwt0rrb
yiVW52kO7fmwO/iuOUYoN/QRTjdXSD31jhVzrP6Ph6svLau4zwYg6xkZTPvGoqa6+eeMsNvHJS3Z
PyZtOEM17TtkeNqWqUCPHQQigPCPoDh0ZxT7L3tSW7dyr2zmAdXdEk62kABB/8+nxNhPVlpLpld8
/LFs4GGnibp/q9tSK5J4S82JWYx3yaVZdwIKJBU/AMMZg8rsetja4d5N5e6OT0/wfIlkcBfkkDF/
KecnMhNM8u4DXuy5wOsa16/mHBOVCpE9L9colNFBK+0DUcRxXPOdnjfCTeTCORc+giGPYvx+iYya
I5AVDlZgEhbKrQyRu53Z8Vq6VROqCr5STNh4hvhE1iAvV4BaNzx1tINWgfuDrL//UZLE3CUDW0UC
GFMmp7mJJCBXfmDfI/5LVf9DMDKPSMUnHSIWM/cexo61Pupb4/JKV3rOqmKuVdgW8NZalAOusHrU
EhU+Sr6FWkcUaD0Gct6FsuWewMtFnXMbmtCl8uKU5xX5rr8xRei+91Sdc+yaY6kFTTT2FRK5Q7TJ
4N7cN8yYfcChuujnF6LEf33WcyxG0vqfjvyjRB2TqsL5Ml/h9AIzFktrm//yH7plE1BmcpjZyYn3
qs+2jp54OapJIU4uKtvKSVawTZwvpGtl9t6C3cyLdO/dh+31PJyNzsJQvYvBzpvk/9MzLeHPmHAD
lNTB7u5Qd6RN5k8v2IUuP7c0+txpzribWx51B8q8gWgTKeid/gWIrgNnfM9IqOxwEEg57FIe6w5q
rY7y+g/vI1WjqML++pMN+8uVOUTXSOkRNqlawp3WWzC6ugP89aIPDboylFJC3/7XJ7f6lDKXHigM
eCMpEhWRE9MPcmIJG2pnz9a8k5EuK4FLzpTBR9a5UbwFgIfC8Ue0seS/hSYJCYeYxH+DlwL1YjFo
Bq5xvVmGXyHtd4t0ypctaqMLZSlLQKKBmcMEAhtbv8/EGC66Y59Vu7lbvUI9p1e2MTEnmUBWOARf
+aP9/7hbbYCWi9ZFGw4Vlv5RD2CIMnWyDPYUN8lg5rvBTC9xOkcqqdomMSA/9ftm30UOTqVP8drj
au1p71Aa6v1AQTT8utbF/YZQkgf4NTQ3lhWisB4vxIXIkGsmQ1ObToCx4uJaZlAeUB3cE8FiQ94z
LQ3vyWbmSnaYr8jEInhL4LR0QU+L1peUczm6J+FQMUXNcMB466lDOq3QCk93cm/4ThaTFfmp71YK
z1A9uSqXAfFL6XAp6eT+5hgMFJEgtBE8x7hCv3m0MwKAf9jTOmxcdAuaJs9X+R1jtqn2DfCgNXMY
T6Q3AHIJqoCcvxlRjM7f2qm+zGt1DeMgVf+yq1SnqbdT++gA0vlDo2RM0i3s54Jkve+a2rL/F5Ho
kYar9ERtvCv5V2U8ntKlE/RlpkUjKiDOdetcoHVqgbI7y0xLNZiccUmDTBL5Ug2JFEbX1xJQeSzX
+aZvKDqAUH5p0LnE1AjHiXWQj/m5ux04cPp+yQq8kYPOHe9ijEETY+9ZsQGZ/GQxgBQFB3Pzh/80
QR9oyurvaTFuyB2T8+omKctIttxn8mySlMX9QR+LCJTu0eFYUFrDXg5kA0MFG5xUUT+brrKUitsw
F4dWcUAsnINO4N/KSkM2wQt96PgX9CNuaUEjnqJcp6JYJWqLoFdaABDhKidjmOZRZmSYvWNxxQCF
wBUnKOqE9Zlp/WVpZQbb8xHiZ6xVJS9kGJxmWCg6yXBv7OF9Z1mls5ySthtypLOo3ubk4zDyMj+q
ywqmESvyUwxH6oLfhnwjMM0d7s1Mhm2ZePS4kjloz3KlbiqTToxs/2oPei/83OPhyGFfFKkJGKP+
fz/Hfei7vGZMQMpk7npfuS2jUwc63uQlFd+K4NDBbihvgw+5TdpIg9SZ6xjjPvr2lpud4aiOXL4f
axEzxz6wZnjcM+DMwm1aWRjJiCWmQTMizUYZBcjTSjD6KsvFWZOABvjiAnPcjE4WjinSURnD59H4
vDpkTTFG0IZq+d+cUgN+nb7G53N3Kyom8GPjCW1wtyCWjCPbPSJ4gkeCSiLbGj0bxAMz0kjOanFC
+udW5evnlT6EtcEhodkNpu+yT6m5KfktszwZ7SLcPdtm/72d1SF2QdOPLi2NESXQ0HXhvr6xpxJy
noJrnOuAf40c8Q/+2hiUR5ybaySdsMbMLZV7TW7XGlQO1gAjIggsLuBeImU0ZYFXgXbKfpNEdXZ6
CL90JW4KH2ABzJIsW2I6BQzsIVAKeT5cmTCxy1/JdwKH2eWsB2eYeJn695axTbexQ40DACM7XCiX
6oXqTjFseTUIM7O+02WNV73TbauRM412Pl23sIzvIzjCf+1yg9t2IB4X4UdLc7Oom7k/PYRascgF
1F4R+E79O7+Sk0+3Eunz43BZZErw7GkoIT5ROt+i9trZzwM+vdnY4OxQgrp0QyGYqt+6Em/7WZEA
e3wPfnpwlOAo05q8IFdDYmvg5Bic8FWYJhC3q/3JW4a0JtYXc0CupGTrJ/qGFlfXIQlSbVAQdTBD
e7wVrJWBri55yxAKIhuVrrgj7IHPk22StEoC4JoumlazRvNlzHZjg0gXjt+s69jdF5JRHUxLBDae
KmViA+8R20JLteS37z3FDtdU2/CMat+3o0Y/1ubUTUTpDHztrA7ICh42dSMP90PqjjaPWGsNyrNh
Js8fYjwRA4phV/0JIallPsF9rkVd75cPKhDbEAzz3f4o3ZhymM2p6GQPelO8iBKjxVj0DE5U/8SD
qyGOR4ZIPLhgCzWz0xjvB2BdmH8O7nUw021rwR4AgVTfNmnTozujA1D+VkeeyFgN7XXDZvmSM1dx
xCDKIQGUK9TM7XHY5CvkCkB+8/3TANoCzRwExIH/6ui9Fbr4T9haJfirwW3h5duwannVrM64GDk4
UXMMsvMQKK13TxA4JzyfBlEfaDSRSk1hHhcIUPXm4woR01Zdf1UQMczxgUKEe6NMQO07piKmhM3l
GR/jwwptFRL22Ho77KZDOy8n3SUPYrhxYeCaPBaiachKxYEObXTtZ+6xuQQrH2kXSXSKYVaRSuP+
+68GecNOYruq9I5U0i/WDP6EKthdSYfuwsQXHTqJ2aoP1USEa2sQj6wSWo7YPeL8T9uF1WgGfmud
mcco3GxUsIMnYhokXscRvzhHh/vZvZK+YI1TcMlcQmD7bCGRr8wL9cOEonDF0MxC9oxpJ+UrLxFY
cK3p8asMazfuyQio9bggSeDymdHvV2iulS1iW7luWebpy2BOnHRKCy7+T6RSWaty/1UBgpH15B7A
TmrvhLIK4tGJZWHA/qUeuuUlcLLnkICqT8GLg3ks3FfwqnJOrFiiYm4kDMkZxfeZa1HtI8vNxvKY
1Evy+RoRN1VknbFgL8iyrututUHXfjJFkZEr+/PGbIqovsMn3R1XMLrHtW4gXIRnvZQEaE3ZQaLA
5jFj+ebgMR2knmYNetF4Td0CURkTaFj59pp6mxjvUErV0aJW6WNL4ra7qoC+BssZjYBlQ23A34Us
EsucxEPUEt3F+joWCyv2YO9/731zRl+p0zbXQjxfBTKBh5jU6MfwSC6ZpJDzoZxqXNBDUFhIJGLy
hjIDHikIkUIpo1i9S79ey7btCdliTldjk2AU9KisFqB9eSoR32Cs0KjEwbQxDcy3AYmWfCE1OJru
rPbl1Dq00hn6I1wlYOOYQbXXCYmqDw8D84dIAenK+CuX4Ptdv/0TbCvU1LY8dsqMcqK3cc7csdfO
ZnpPwx6a+luTcVfkY7QZKs7fpoQffpcqNpXlbXtLB4/prf1Di/1ecrRx31yVcZstDVVJrBS8n9Lh
Cv1AbVFjs4myg4+0iv2F8E/TE6to6tgVHPTOodXhqlwBvI4qZTRlhL/R5YagGYxb0/kur6DqCVFX
3DepV4VljWOUxCTfZwogSL3MEEb9VeCg0nSbLVuadFs8KqUgwS8MrWIrOq5a9aOmcaVVuK3uMRTD
j8jKrP5Q1cg/1aJng2db8+Ksdp5Al3lydIBzy+GaYhJ5tU0vZk6myd9HwHMP5cGNLe8DTjTG9TSP
MGIzeLuFXDxxx0cckvGQJGwbofgxI18+Lun/P4Av92trBq0hZSaVwkJLxkNXmBziHbvSKdquPDuZ
Cn0fJFy1c60ETNqfIl7I65yBLVC+1Nxl7yHJcnODhrtbVBShmk4rqc0fkLjo+goHQNoe/I0p6QBV
0mLAeQYxBUsdKanmj6LzSy0K5QAzb2tFgbF0IF5kh5L9oNcvLe8s8VAa+fjCeDlX+zUtdVNrfxPB
Ukuc1nMn8y9ZUSnCCOfXpKOUG6b4gs1dkBtQoYTBn14ZaV8JOS7VKYqnLHl7hR0BDZriV/ZMhms7
ELPQkqXGFp+nHMl+zpZigRWhuPbETPUlGXXK8c1Rp0MM9TPD42HRSrH8HRN4f0a8mtIzdkm2GxOj
b81y64Sq9M2VvYdWwtiozlKDFozM0/qnjS2xKGAHhU6RrSG8PhKvn5CP1mx4NEBGqaZ8AQwkL3+L
EwocN9b1n90i4R9tEBDkjPMzlfv6lIolUGmixl/lwNjMwdb1DPPUvU3dE2T8tAFGbiqLGbIwF2fr
z/BlCFSf0lITmGA83x+mTX+XTOxJfziIoHLX/p6RSp5LZBQ3EXrTIXmRnxK8LcPbwBrhBiiyfQO9
39O1V136PB4TTrJKcCuj6WvRUf6IwJfK+0ZQ1J2Sx/OMXvke7VfV0Ei44r1UoNCK1XqWQNcxZ2zq
dcf2R5h54IskVKsI7fPo0gSUWqhSwdB4uf0euWiGaGGG79QZ9UOTgWbO47c5Sw1kcGHzMUm+cXGf
lU4luThg1rcQi9aYrpPibLkx3efD+mbwAjfV57lGg7pAWWhAlTGsctpKKjl14mDc7AKSiZRDwbEb
u6VT6s1/K9XT3sWBZqsgPJpmfymYGPqfUz15/tvunrq2MdRm66sC0HptAo2Hoc8NK+DXAbwUcEjq
99Qe37T2vZoK1jEVgVYTga0T31U6wbcAErvEpM5+zqDyuFFZF+ONb48btl4w7BPjI2tl2Tyijauy
q9W+eIdl8uqDTKT2g08B6ab7E6KMwJ3UASJA1o2Y6niNhELdCo1TdniABe4Ogm4LfBgVwL6JFiux
XW9a8qE3knkXF6xOK6RZtseKHkMVH2zj5LZm1OCd9QPNn1CVTs34XEt0bXN0dcmLKLeI0fF9AZ9d
8BMyxPk2ih259lnqImgPOeQ/McwtWQSE7xLDLewvFsijoNu+YmowMX6l5UAnmqNmzS5WfCUhNScA
rOxS9otozA7qbH1jxe12fCd3vJtsTujUwFNJN5jETXuTTCsvLVFa3JT4b519Jsl1WrvUMLAHK+YB
77EpfLXn4KvmKmh/SYBUrVDGJX2xYytU1XfF5RhcysDsy6wOO9qoXRd9gTQmP1sRPCxrV37dbCyH
gogoSC769v1JweyJuPlIfdi9IR/tpkw8aRT56YJMsQ1Xl64DinLuG7NuBE0LE+xAgdgUCjDiDUe4
SCMHhFQ1sC1jy0DpY7PG54cl8AtlfnZXFb6ENkxGIK3XV9fhN9RodSsNp76MNZwJNFQIOBLpfasd
m7rjNaDvrHsr+PTiuxtBvugtBdTiMQDqTRqz5x2m8zA3hraJMxlCkJN/MwM+O8gc84c7IbgRb31a
sB596wMBabglg0bEJ4I1VDA3vitFCRoCTzAqsKcRTctpfoe2CMfVUtoFdUIeptcFjms0ISUgaumA
d6fTUY5g3Cf7B+inMwmyQ2g9yEjfAbr3/6zioo4X/Y+wNpBiSXP0uPFDxrlk7KCj+KXeS6aI2/C2
xRUbL30YrOSBGYlJj2cipf30md6rB+QDrPPTcJASO8/UXuhNvf2rQhUvg8YU1OX+xI4UR7gPcgdt
7sKd9eEfO62eoPYztIRdZRBjZ20RNJiivh72vfprzDjyRi62MlXFEp9GZQ9chXkervBedwkphCIA
AkJqgniR74QKzE9vgOEacq2hb0iLw+5EwyKJJFuNVZuXeO1Z67J1hGx3GTAlSsAncOneWQOSkEUc
pebvnFwQFhtAR7cfeWv/eNUDRn7uICYH0dSGV3t2TMb/DUA8ptdWsogx+EKX0adss0GS1uSkW/a+
17anD+q+CM+yiIqPacMscKvNKQGIoXhI4Q57bgYzJs9dALioS3QzWJfLS4rkAfrb3F/7AwWcILps
h8auivakV7SnyUQVHna7UfkWaVDtSUDj7GYsvHHNlnvXGGiy6oPdDeP9YpC/gRHCvY5bxe9lzRR0
sZBuLvqvvRjPjjNjy0gEIBnBSBbrYe3AMwz+yHYBLbEiwwESKHPw2Nw4ttEG+UeoUluSqIjwJcl9
mbevgoXfjXq/T23hKqxz1L5V61WjVtz5JhmKRY0O2EKoP0pkcccAhr4nfNMRUsj2s8HGQ7v9sW1m
lodHh82jskoXiDe223fksoJwdFFR0G5lvD/TXNXUDvn+hT/3/vrKVobUk7S2pDz8oCWjQHukmFoW
S6AY1cucYv2ynj5dn5o1isdpVE1vWwlfBMygk7peCi8/3hNlaXZxY5VCLddnSBKqVjXeSV3JDwYp
rLEorp+lcYgbx3V6R/6uPe1tymRJRGlBMVWM5nogSN+eck0Ac0Fgbx6qtKEZBpRuPE+p10cy3JxD
lKFMM8eZCqt8mMHBZonga/CiFtnNkFH2fqT0smMgwwCFXJ0AJCcnFzqoPIwUXCPMblWxmrP5kA4p
e6CLA/GxFVBrKon0erq5rMHntGSG2H7nr2/GBTjm0NZxMYJVBG6yrGGH69rfqTHi60C8sdyXNyEs
a+ErDGLojoAZVTCNuSM8h936thhK/6ZTRDqdjpW6UlGYoWMICTu++01JMKBJ7oTdNIxR11d+PfOy
1LSkWYbKas+jubXuxwB4K/pwR62i0D+0mwXKYBYBJJkfhu9AF1rXOZ8xL7xBz+tPTKk2yVIPItFr
5V3OF/WJB7iCfp/OHfN9qBm1xeqfw+VpJLxxDHmvxgnmAPr98Tklh4yHRKDT22wBfFfvGz7OP2+X
0pz5yti6qRe+Fxd8r9Q3S/balqNFu656lq7YqdbTT4Gmfno/HOJZAmmIe4sdKnrRHkesyFHuV/BB
HsKww2yz+86zlb9QcMwVE/p/dFsdSMQ3s0tO0Np4DsD7g6pviQmVvEN35f+C+4tUIiFY7wR3lhjb
6wuM9xpL3ZhH62+udYiBlvGX+fU2XhfQFHf9xCRRLMR12w7Nq7Q4zUVc4UK8WCMDLNGb5eVvppIP
RBgCmvc7aNMqIUqFi2E8fE5eoHF/jPKUlZMBCY6TyVzFq4OM96ef9fow0Tv5P0cBKVvE6MZsj15M
o9Y1+sG9tfSkmO/rB1imLN9YpmSQkHfkJofKZ/rwyGsdts3NDDmAMSu8is3UpAzWrEPFUQ4foLx1
O5htdHiecc6McPHFEKX3ATbcb1CYbxHKCRQhP6r3QXen/bR/4ZaVpEpi2aNDtwfI+q1TwMMHnGpB
SYfZehGDBJfgFsbNX7WWKacbmMXRhKPrgyQyDJ5PL1YmCO8mZNb/Oevho9wyMyDbysbVpWoAQLEH
brKYzYRj1A/O/+yBMbBvw+wUzsv64c88kXRS3NNke+cPnkZp1tdek5nSQAaqD3us7vv1L6Ivd/RY
AVBDnANrdIA5LF69BG1WEUT2pPAnKrxfSIa41N3YovGoz7YIOd6cePEVtLiKKoRuHHwq4pas0OhM
bqMNtOapuLEcou+BffG1c/S817gM7fgOdoW4sva4YcYqv0bpfoKPd8HEWzfwemF7fF07gcI21E92
YLY5flyTzb5CHKQa1llTqL5mzKc/PmycsM2vXBx3spgExuEe4SOQUtXBInvrU925qbw3ysz0f+wp
qFjP5Naiam11vO045+MMRfoIMWfsaOnAZ/oQFTvReO2yofgR6SmsRFwIRlwAFhtFy0FOibYRwF7o
3ZQUpLL98Sy4HEOKWwJNthGBDo8E5qReWCRs3CelE8TO2UWlH36MI3NSs6SNMZhIDc8Du8Ik2wlw
EzoE6PVh8LMG6u8BN5oQDIeOPVaLhsimayDDicdIq5czFHJIM2fPbA2ZsNhx4o/YuJ4opNUvB9Q8
Z/19QhW778czV+kO77PmX3iADhIWrdmLWR3HK6G4M0siUKOK0zOkxol6uKKMzVYGt4z61XjeRm2o
+Ske8cDZqhvXPweEA+LZ3tQi/eMxuBqUjCi0uZsqFckdzkjrI06uCXW+DP04c29T4E9Re5KuJyW4
XXYgzUmVrxskdyhjq9f48aq/OBgubAKWC+k87zBsAiDwTUA6UnraoF/XysJUNW+/Aq/Cu/URMys4
fo6sdyzRzMZoA9nklbCLIpbpg5Gm7m7g7Q5UR+VFXHF0cqwBzyknTNWnWKJCWU0XQlC35R8PMgCT
fsDsPXurgMD8VC9gh7EFejH+EhWsJ3Hx47bSJb05tCSkIRGwFOkBlq3DHFtIMPWyqNaIsj+mpKxY
oyOsgy9r/7rSnR0mCqTMI5sJx4XhnhFADDN9lflgbj4ah/Axf8eeAl1dASKAGyn1PfYbOuxVW09J
PWZR4PHbi4FFrEb6bnnxtJ2NNJqLIaRFEQ51/Q4czngwZepktXOBAX0yLIqfAq4GfKr/QwsiKCxU
Okx8NbHyvNSRobGvk/HeEtsGXqFXQeim0a2xvxa4P2hbmHl41V0vVw2e0tDtI5loJqbMoL9K0wCW
6Ocd5eDm2Ijrroix14xfUQADMpwrN6ySvrRPEEwdE6txUlN1ZLqQIz0ouSMtt4d621C7SgTv9bCg
8UdVfUoaj3qAzkaeCJcXt4WRFe49dpm6pU9ealThVW28bvWqkd10tzQ9kznI8WD1SMM83Ojt0pY+
vxYlfMOxqewRf2Q/iXSysqHlDnbvXRjcm2w8aQAYYdQB6h6xhs/NkBR+3KZMxiA/M5E4upykkbCM
K/uolaNH9obtJjIcU+n1OOlQABYdQmiMwvL8bfUpcLLXM6iqKxS3+/RHaNeSqIgQupAiB2gsSub8
LGnbgRyOxKpNFidteErlo+YEcckzvk5m4WAxM2y/0E2I0IyF2SwlsSdg8M46omMjFVkPunmAND6E
UCk0ehn6n/zZ9/6Vvey2P1Ns70Hc1opXB5dOv2oU49sygtWhtdXoyum4qGwnFeDmamwKbCTa5ORB
HwZalRB11zNQXB5xsBIy3dcyRFjTDuPt52gp6MkBfUrfz6X75O71RAohuuLHz10nKunFTjQVoApr
NzV3IiS8vP+eQsF51bUsvKN7OisTuhu+3NRRN+5zV2X4P4sNCLGkm5Iwzhae59UBkmGNnjKA2tin
Sq/jxsqvlFFthii0UjDhzhc2t0gd2xM2uEhWqJzCNbixLClcvSBjBTZkC6xvJrqvWfLQjLUqpil4
RCptmvZzuZPrN5Q4IYlvqMVsw2wxg2/8oI/TqJJn16iKai+T4lXyo2ba4jLZCIkShORqFuMso+n2
kPokR+pg0ZSSWLwK9zu6Qovca2Krhd7efrhMsWpf1Qim9cImvfngn+go5o0/vTOnuh4B+gRKiuk4
YgacFEg6iJB/2KMK/IMJcl+EmhrcYBQWWkhRQ9RjznX0Yvy9a2j1setUDbNleg2IfZ0y/pL7gYGG
qpW7ApKEc5PyJcULgG5/4iiSIFSzY8wNH8bR3pFTo3MfkW7exJlGMVwqLcLXTpzaMb6obdeik6s4
c+39YKZfue1P8b+mdZiNh4/g9IkTQ6DxF/FoXEsghO1IOfgx1MC12FCL6F3sTSTaF1LlED1iW5ZX
kK259prYMCyOpc/x2TFZEsP6+rZevDPdkIgv0zb0A7gfm2rTXmliLTg7MzG5ffH2eeNJxE/dG/qc
nBceknn2pfH9+oFsfWbjq76qOOLDfy1FGMRyFYYRFXbsB5C84JL0EaM2lVW6m33y5eLVrBYtBUl3
39JqX47o5IaHHDIMaCzqt9z2aLOKecG5lBJHjj+aVYva2EAhBnOg0/q8TItPqKp5WfhN7NOesTwc
tr4w4IzhpPCSxBp/P27STYr209UAqwoAVLszSciI23CS8HZxmLrPrRH0F28jo9D1bjrccRHd6MPi
AF3RA7HDuKuZx2yxnmSCAdS+XQDYyayNS09r6E0t8jvrOG2PIxTNJ2N/eiaLojCA5q2JiKaRCaBd
f0/H4js7j4r0QuQiX6H8kf82aT8S/FTtp2yx4pheUeA4UOleDuOtwaCCBGxpj2oiy5QLFT709myg
pU5LbPVrUEOOLkr5mLqiQsdZ64GyolMEnglXC/+4qb494Iuaq61SMAOONmfI0+MHu2lOF7ty2IG+
PbqzbH82F4qc3u3xUmlMrKBYJfcLoxwOzcQAVq/8sbGOrw8MumNEUJAVV4zhpvlF+MXq4aMB3g3c
QdD72BykCW/TW78jde+kphHceByV3ufPNxG/AYjxp0rZEXPM9Aq4kIXDwXmeqtQqAVRN96G0+JZ2
Nemr/xqYRDYUog7ESwB3uOkV0aFvUTWbviSY5am7VhDhpOpIOgeIR1qqrk1UOUOERkvlD63xDmLn
XLPs7tlfXIqH16Z9x1M1WSvdp1o/4bdgmAYIXlTZaCb3Am9OvM6llq1ExWa2QIzxYrCzrQ03W04k
6MIyqAEvXLO5dv+zK3EH5Zd93WKlsNR2ryFkBoY0k6tVNalkhwpQ46VEEr+ETavu97UZW3TccXqv
sAOJJuTnvt3Ly8Y+BmVcYqufPQETP9uv2JiqNMRdPPzlI1eVRI+Pko5S5iS2ruQJlygC4c0B04Sv
3Hn5cp2VBnF30Jfa7CS6zViehRUrE1vYYaZFfljBOPT+E7jDKTSbA6Ho7Ns1qFr9OJ+IHAuqHgXa
tReK636+HO/vfxpp673o+h9Q2O+EKBEcdLzD3i/rSOIVCQU5wiB6FbEjkGiXr5fPWBkw5fRpU38v
I1InGrBTdOg7soWBk/Qa3NvNfep6EXC0yV1b7I2+YgqgYPPHJdt2/58O6ClB36M1wedslTJlCZYo
ZVLJa5Vzw3NhOvWPoMocZsmSRbdGD6BeleUgiggBKYGBFwyFM4006Kg3XJCcnnxBeWSzIgDkazAa
DdPPIZU+r7DkvYaXoBx8HCGz8k8BKmx8wagg/rXPYHUe7IWcTZD5TzKN3jZ6aPFjzAQXMNzZmgpe
vPNIDK6JBfYoNBS9AG7mBGmVPCUmXc87YVbzDrBhGVSJN/gkkWT6/wYJCWJlCdaT/LU24mdU7Gt6
CLyJlA1/LGPSo9ARVy/KMg3ZuGk4wPJyFi/JxpxF3akgHjc9nZmH5YZwG34ydm95Z9NWbHzpcUgC
GRn1w35GweSnYPiBCYM2NZrYrsdphG5SMEwX2njfAbQ9B/zdpmJ4G571Zdj+pjVK5b6mKMo7aL0h
Wx6IT811pwWWFwzYoeXEEYG9Rn9nrVhmtD/WWGzJxFV6Sa3tUULe6YbbN1OZzDrVQ6LZNyZ7kBvq
FY6mZABqbg4eTXFgYQEYGJEcaGJbeRzqwRsFT0rt2Mc2YHGAQ72Mnjmui80hZjx7Rj5XX2XMY7Bo
V201Ev1jkZjxfxROY3A6r4eMQjRZUuJ7bjTk4lY2vJAhoBP9/DPxq6Yjts3NhCQ7VzjMeOWoDtqX
cYfeyHq3Negh0ljdVCt7J9UnFK8LSLpsnxeq4njHKlBG1zpdUpnGW4eI8kHUJ9t7peCjF4TQNop2
HJiDZ/+bv33ymgUE45Y3qTBMDEWU1fH95gnCWw4FHrvkUbG1HqILYB6xPH+NiDG7uAx3V0j71NyJ
+9N+fwi0J4CP6BTHBYQ+L+zpJhDT+8jKTFvkp9NSSYzX0SOCGtTr0PK61PVexCaE8PT8pE+Jegfq
YEPZAgfzQd4SUl2IuTctwzQB0X1fhgfBqa38PjvE3zC60Ah/80fmPswB1Ajtu7vAK2MCAI0R/GGv
IYpM/PufUTJo9Mx/mw+TN/klqFpw5ecDSXjDlX8rljoXhQe67vW0/5A2LW1JXxzKN0b8qTHFDo4W
2SSRCCLGx3SLH1JpBr2dWQtlNmIXCqArDjFodZZOhO7dGHELXHeB7xbHNIKD96F5+WP5LsRSBEEu
sO6CoGq9cnvWsV2y7e/dKxtAwI2zR74KfwrkuMOvvmj7haGIi/GdSRmnHyUrl1zkfzRqwW7ognKF
tdhiB74NzYxRLvDJecq2OgNsh4Z2127GsT+pLqAZqwFVqXznp8t17+VzNiDh8GlQlmHS7rWjvyjz
NjEIOEes9XWnQoO4lpf5yNzS+Ahr1pong1yHbPFmrS/oLZSi/41ftMyBQksDisBBfZ9zurzdJY8j
Gry6lfgO1EjBknS03ois7k4rA6AGO7x0EzHgj07gobHvd+V5Iaw7x4j5G0BKTH0tPZAZIx1x9WDi
OQNXz2Vym0AQjWMV0kKJpy4XsCrJBhuPIvvCFT1ODRZeP7tO9Bkb4/mtlq+y8B4yrmie/qzyllFB
bM33+UhMniOFI3AXYZJ1WpO11Ox8ElMURlhaZCeJ82v3ibMz1QG+ynJ5OJiBpyw/GPMrgE3x7pH6
77xmp87EGOqnyRU7j2xhmrbwYxL0EEtO/4Pnpvk6Lj4VqLyO5KIIeHhm9hio49AZuGxED/G9ik0b
UKJcZT/5qe8FQti+K9taI5hacnJfjnwLlWxs8KwuRMNC6nUVGG+wE9d9oZgpGzpS9Ui5RjF/9OoZ
nU1o6gdvb/i4wrO1w9Hfd2X2f5NsqGW7fCvrs05t514f/r3uggcZdD6V+AJvMpAZwDlXcTWXhLKf
dRAUOyra+I6s5+HiRWnFAnTb68PS4fq601gS9m2B0rGiOtEIEPBBbm8IPPwi7BJUGrSv1lK1DmVP
xJ0/6G1iOa+9RspjlO3iEu6mJ870aJ8VqY4Km2xKc+PVyoHbilgAI+Hi4mqsVfevX0ZiV1W+ZG4k
kR55lOxCYdSIKBZ15qJjOTz6XQKABi9EVSWttKcdiv4mfv7u3XdLauWqPReXRuzFeG3aViskDJpQ
kjLtWqFycvCIMiAq6/XYkPoOO5V1fXnc6pWUVTlU5b+xuVOMw7jggVemeyk0OqhO9GzbRz05UpBN
zdwVtJDoxua9byXJWSJ7q4shjJsw2DjUS5dQj35TO4uTGrbGFZukYEYllaMxTMvFwXNAGvXF0rjz
ceJHlmYdBJNvZv3fKXR51+hKe4M/oMe0opXkBloQWJ+x6Y60wvP8VpXLZoXVQ0iHBcvDfIvFftR+
+F5rLOA11wv8ctJsATdsMDBv0QMmilpGFdj+nYQuyMuPnYftKNulOb30abPblBhO9rSEDIKQNjE5
1hJ2FmAw+eI7x1dBDD3py8JyWthjmHXRH0psHNkCQr18xb9lVIJJS2pjywBEQ0QGnWTqc9y6EgI8
1DSAjKakG/XWiIc4mkS63QhCH87fP68pr3sCHQMgbDAj2B6gfCPjo83c+w8Q5vnYkqU16eOszO3P
b5GhItPKYu1lyovFrcKKIzFCLq6/XVWPN5tVIPOApLyCIGwKg47dg1/L3Lg63ycbjl3pgJetANP4
364chsvnMnNovnpWquWuDA7WPozfVySQcq2XWKlhHt2mdziY0hDnbOLxenylqbZdsiikfGKhW/3f
6NfDJ7s5h4cb0sBlROJg91uycOoBWdtO7s38BdEWPAw/Gsq1F0w8/BqjT/nmF5QdvLprCia3HySn
SLIPxVZpkXRq7xrhx/SkG2jhyAYujnMT/ap65CEkf+winqfbCtCHe+xn05t2wwzu15hjqNlvxO0w
xlHkwQc5uKIL53VkEI8QaPRC86isfD6Tv5XhaZP3Lpz/EegoTrzqS6gPP0qacBG9pTlDLq1prfct
XOiMcW2BDWnxLxPdWTkFyA/FRFN97RK5+nC9+TdY27incrikjQGuSduoPK6vfbdHJ/IDXNLE8XK5
ygZ1J/9EMLqx4E/orYQH5G1B+CNBXnTRv1JFLyMHNmdQtm9RLPP1OKyrNnWKGZFZcUp2B7UVJUGA
VELEayAtBciDvyqdpMpesFb9OUqZ4E4AzyjDpaeXFt657clm5NvncD8QUZgPtWKdSz6v7NpXt1uz
zp3DYGJ/yPjJIZV+a99toX02ZXTa85gutrjETfCT/xeP9Coa0UrYLwAY8hyc1IMH4t7jKiK++E/4
Qylr3lJC09X4vO5Gn+llwbCRH7kuD6nzQ69rk060Bqo1g8J4qRd58YVGbF8U4Dh2hqrxA5HAbEtZ
PXQnGpGtWh+fr2wCbjUuSZO+fBw1TReK6LslasvPYjRmJZXnFkiv7YI8uwqqjH8Ke6TdJhtcFDjh
awv84MmmHzJBKaemW4+or8dMsNfFH/1rwpZr0mQ2GsrUpx01tCg6wIpPQfKVjkFbzlvP1zxJE6mb
K5dMREeNwPQ1aj4D+Gvt8uco49Haz0mm/i48Kc9WSwHmniy46Ij9P4QuCtsK6nfkh34Quxhbpr/B
Ntjel+447wX8hoJsglvRNuWT2B51aTOeeixeZOCjQiDdQ2eTTTqu6bQ04cR3zt2xSzStcRFmnu8w
xIJv10YUFdU+AyOUCZhXmKIf6q83s9du0PV+skKngNt2ZByQ74/kBDK7jLUXumM2B/nsCqMfWvdt
Hf5marxx3CKPMccNHvoJ9Od0QfXIjMO9TMCVYh1JyLMX/bIEqyoGQBJRxNRpztdINJ7yyxy3P3k5
C7vYWhJaQSRUwmff+LOTeZ2flDYYGrel9G6pdBDK0tRdUbXuvHj2qQybGUbZ7eQm4RJRZ0jGbvUr
oooy7nn1Gkhb/LQ9raUzBD6FSweKFOQ0eLyIPmWdsb1ew3rjv1DDThaBXfiRTTcDpMBuM3XVT9b0
kDXBRsNSn+x+kY3zVQDyxmN0d2PR3Y1796yruSzjyi8BJaqPoaGGnWG8nEBHhFN0dLZM13Zn2DOj
MEiERjcx+TwpTcCz8rB952YQJ+VJwlDK+V2+/YQY4GPL7BNNSI2nb7x0wnbKJld/0wPkNBzhGYvg
GNH2dMEIeG9g3HGwCjicPqhHWiU70fA2zY3zPyT24AkkssNut5P9gA58m/so1w3ErgEYhPDZ3YBa
pgaVxpf1S8bKijSOg7YduWhq2ok4/QwUSbkKAZyn4O9nTEBNP1pLUEpY6YKF83dU5W7mg/kc6aCN
9Fh4+WfRYKGZPVcy3+Ob6/A0kPkt93WWAejSFlnEmnKdWM08XUFjF9v/FbaJpkLUmyZiMAETbGGJ
tiXZyINO0EvmvTPIna35tPI7hXtf8DimoBPDJS/iYc+nNVhSYVkjcAauk40d3iHQQNbCQ0s3vjBx
ShEr5S6AXmvxZf+oAeDvJy3ujyI2cIGWU6+ejNpn3WEleeCNZ3irWoXBViIZfM6awoXm6QpVALHu
s2Czik3y1Bu//W1/0p06BCMghsWO3DO9wihjJ2IcnWL075OevVFHlQR+xnAuf5iXOJyvfvX0j2Bz
xAB2xBLtC3IMuKj4oEfKUFOMEyu/ofg3HEYEfQnaoSx7c9FhLnC1ZtSrFQ7kvkOrO/STGfDhIk2l
yN18Ht5sJva3TKuQME10pTmZXR1ZsErvXpLAwpSjzveSttRtnAKesJ9560vGudx3LbHM7b05psBD
FnV3LwMTYFCkfadpQgYRpiU8t+cNrEocJclYksPnbZBqSR9yUMUu/cprHQLII51JBFP9g2y1Koj9
Kjpk2s+tiQojB3MD5zoLiNC2NON+OW0xNcYCyYvESMKMIQhIEfshDBKcUJBkQTPzrLhXSrZ8Ow5D
kf4r7YnN+57eS+Hnvc74x07e0H8hCgyWEf+BBfvHnKVEcxja+1+RpbZwL0CbSz8McqQzP5PZXnrV
ft/fjqT06yqPw3La9ujOW3airq68cJ4Lc5CmGujpgGEpNycnpFAUbq2vlai4s0kJG5KACCpWNwh/
XX4U+JEyuj97hN0xj3zVBvzuC76tWNSOOeXHeDv+9bFuco6ekJQNQrexRvalKoIiiHBP7poXL9+j
zWGFf0QQH8XvOYCOBHcfKEUnH9b0gqzq3N5NJ5E/7w7oezn7iIGNhvRksaLaXY5aQigFfYJigqPb
cIJYTtOLbkrVJqWw4GQLBc0DMkb438J7wu6K6QfSYxdCHLmtAGCm4g67Su1WCGztZGqyByt49MXD
DFKug2NVnizDheM8y3NJdAuHrW5kUiH2Q2VXP7TqpT41Kd2zcZKx5DW1E2hGmopPvFEdxvuyq8Nr
BZBiiM1GXvLil9tlwDeEsaSawpbvyZna1FY7QnBPos6uKYvp95Jk+Dov/yhLVAh379JP5HviZNb+
mZLygX9Fqx+g/lTLi1OXx8NJjjS/FxbI0MCW+kg7Hl3VWi9sUNWpPkmIwzMr10b7Dbje7HET06dx
ELLE9aqdepwxh/eOBQl29wtZ6jCRKAm5tCeLkXPpD61R5JI28Vx9q/e7BpTkun/9gKEavALWEdvH
nKIwC2iSqWMBVCgrMM0FJqucGoFjsCItcoZJYwaZNfC1q/tsTgOenDapELs84DxfxEu3ZaFY2dB6
vy7pNALZJc+EiHUK2V/4fqjc6AHMGllRL9heMlg9hsCamKsUFX8P8qfA35zlRhN9UyABR+1+kNyU
WHimhRIKP5W3Ic66YFMAd8+ikJIfM2t+tldqV140LgcSlxJCHSTGO6nvVocJtCeWkYP3cOoHL8Js
GqNgG1t3L2PjGGcRwq+SjV//9TG8hOIJgDtcZQIkXt9kXuhHKK/dYvGi14k4/qsqcZMbgvG6atkV
npwSdHbumc6vsLJbGRo16mwc3KKM5OAZduECiLBPO8USAy+y2jNhjBIoycwm0XQAviObyMNVOkRl
4i7VOCYOgMTyUk9Yp1405YiJ1rmOxnfXwR7zYvkBa0rUUp3NKcQL3sNvQM6Ae6N48eDHcrs9HnQZ
ghDu9Myni9MLpj6GeilMpnChXq2vtyIPLysvwGlE1Ax8vrvbI4SXWouNQ3Tb5EcqNxGGgz43vqBt
IT2FIpuLzUXYoOUzcvoSLFXHPxcjdtDDfehjku4dF9Qeq2ltn6iaMoS0jl5DhxlmW9HtnGLMGxt/
0J3NA2jMnaLeb/+jGGDwcHQ02J2RJ9Wp35PwLSDqcYDN4IwOu3GoSi6K1l5N3QuHDFscFfCiVY9x
at3Af5sD7dRHQCN6f6/1gMrRunG2NnW3nM1Ps2nbt1KMzcUK/2GjIZZS3bhdG7jpu7i+DEeMuZwN
oBB6Y6qEvMaupl82lK1gxB8y23L+EJaBzhdaUp5iVVXgiyIpPfOTbUOIqKjXbPrYqf/UsRmoRQOe
l8BQSMDbtiGl9MS/8FoEFp0fX2X0ePYw0sA1JxY1YKgcugQilvBWSnO3FCzGRBFA7IsNgMBoQ708
JJOZ8t2K2ZYHw2PX1iw4RISi/XHbIBE6ld9NRmHojSzfS3nizXDi0oXmCXvhUbbqgZkf08b7hIX2
ohmie82yDcnqNS0rJiE7BQ93F3Lf2DH/nErURC72NspdHayEwVSS5nvWPp80ng/wRnATP40zgc5A
SDf3AFAACphJs9QvFVGdD5MZsw7ViClOaXvLSdxW9/+NXUTyFfhohx0Z3lgwFzHtokJFBCmIUy3G
sp8jbNUMBikSWdWl1X9p8A/WEezbT55r2TNGLeC6V/PvkPebU5jNwE5Urljg32IDsM0AvTjquvC0
ouTPG/3CFxRSDlQ/kCq+8wGgDsub35LvQ9qfTwu/JMWN7FgWT3KcC8RSM85apLwkXXkugWVMwmb6
T21F9Ak0Qhg6Egdl7kOoUwze+JRF7WkiKmsBiijlLBzzfUWrKsBU3kP9ZLg8tuklUS6Mezs9D2WX
H+DpnbLGXj/rHi0knWH1ZfANPxas8+zFIvc7UnOxI4XWy/xfZdwi6J8HvVKvak2QVxkZNwsziWbF
LnufyAX/CTieT6hcVLcUmONkO9+M5wWZ8nSy80hw1eWNUTC8lxxQVhPTZmIqIhdxwsEn0QKKzoKL
RHaUsoigkUOqGeBUTD0E8LPqeeSOlZ+5s9Bf3PlfnGd1oiQNRadIvw4/XjbwsazE6c/Tu/h4cAP3
/mmcWCU7I4iXonEMokfYhlxmJR0ncGVN/4yyMPKc+f7qZdJQT2wSsVpBepOMYVqPwy3RfJuHL1Ed
YF2j1NyCe74VrTRLFLWp/twBWM5gmk/GuLxmgFk1Fgv25+DS0BOeKYit5Vx3W/aHVLUxNpSYNH4N
YaE1CGAkPrq/FMPbjoMMn1iCkAHOlcdHy8NHttJ1UmfxlhHR5V48OoSv1dNjHXuylZo1LFlJCEQ+
Qs7SjBUxD3xs6MmIBnXaRjPYhMVxWpzmsQm6Tjn8xVnicPJeCNQdWz1mb6vMHWaUbaABOUIw4yx4
Q4+x8wBjqR+VEXTnmhqhascaE0RgtUr4iQIs438AWHw0tj3Uix+fnBroYe7sf5zr43jHc/6WpxbE
WadJSJ2P6+a6RpDnUxWMGRKMrs5lNuccCnK71GgHV2uIFuzdZK2WUZj9DUk5xQigrMIQHZnEGj4+
3EOaLslZXKqa+CCs5HSfqRUnslG9MGd0z0ScLBIOjnHkcynBD1bl8Yk6M2qxJ+I7NC+bjpziszaC
Pnlau5Zy2SxYa2TEQ8kjzVkMwI8vgmtk+CzaWotXlvrhpvQW0/oJcaR0uBs5I3gn/ZRWAeIVdEML
3E1ohheRCHeXf4IwFWIfBgZcfrom71BUOV/JLjioQTOQhOYK5pPIqwauodVaOI9rxewDAroNqq2b
iNbBmm/AM8wuJmWNnAQdXEiptrjmodToN5A80ffE2eBvbVg6PJEcWF82M+bkMzo3MckLCSkFq2nv
hrRf5rIgpStqlG8J4Oo9JzKEOqaUU0U9KqSzQGwf7wFT+d3gEVPJaN62zXI6Xsy7UaWfFVPQjB5l
xFtN//D/L1NqbEC0M/hMqVQSmpLCxSGBKg7pIcuoWFjRKLRl/FgCmftPZ/hCg72n4Z5fKoCaQgq1
ECg7H4C2SKi7GexLlB03uDXz5I9qx6GL0b28snMn0E7zhi9mhaS+M3eH0SghEO0AQPOQQ9BM+hxD
RjeJWMTZEjR7HXWwl2QE59ugnyPVmgX3KLgH6tk9jLXt3pZx8TrZfLI2ryH5d+welwZM7wNfuDtb
Jr5tYU3VH57aAnosmPqaZ1q4uXYQTUsDTfHLpXESDty59vRl74neM28nf/rjTPb6+wSE8ue0GIBm
BRKwy6yzhDfkIzmWAPgr7utD1PdJEsxxgg8nhYNvY+b504l6ECtzmWVy1WjEwsKeJjOPtGcVna7h
cc3lrve8Zj3/NRMl0OK0HsO2Ir916Z1mPd706IzZkp6OL80GnBNamFLooZTvlRqGcYqFc4QtYeVm
QD54XuupEmLh28LYpePGRG36sx1jOvlroadL+87JtfbRd+Bs7X1fuZZIhJjgWAWS85dcnO1GbEEZ
hMsC3Ejh/3zzi04Lj+O3blh8o1MAB6fKaGML5osI/AnjLCc3dvw5c3eUKZgM/ndP3wqHMGeM+P0+
rgeCqnitePQ2m7g/MWy4jkAvuTpWRRV3QhZc8XumR0hnahWjLEIJwBCZ37V0LUQcNGz9luXV6chX
oyZJOFliqb92Zyb3Q0V4AeUtXh2XKQ9E9ICZSvZ3rg0EVJKlb4mbgSOUqRSaM6/JeCHiyHyyMGPJ
npROhvnapSJBwvhE9L4w74LyfWbctwS1nClzoxQtD+uVCOiMsrXjfK14zJcVQVKKiBVzesKwBl+C
UsCj/eR7OnD0Vwi3R69nJKviYFNFuRenzGwARoWVdWsm7JZf/LgjmEKi9+7AEqb/pt5oIuKRG8hC
c1zKGyKQBYnZ3r+s3LX/edhrWd33NBHI3uFeA1+dTlx4l8ZQrs8213rhU40ferfzZje4q9+dcq7E
fT5JqeTX8suQbV9ih6OMfcGZYNc/iwY7YluV9IWIjDMc9xDTbM5TQvid2U/0KCW//1K2w/tAojDY
xAGFqJ67iJcHk3hIW1BrWubdAYuj+jIYXaXLWFBt04LqiuBbdMwAFfGZZd3/utxP0J2NPwVnY7Zj
70n1SXVyM4FxZVx2lc6sP87sVtV2EpDofC/iIdOT6Hey6YebYp+/x48tnusJwV/E90+zls3jhrVa
9vsVQbpNPNALKK0rAIvNOwpz5gqVwgpbT+Oi+rro9wTOTfH0g1IUED2IKc0Wdz3cNxXCg+egOpQB
Bi6ZjSQVxR/dvbom9dz6JN2RXIiZGXxfAkd0wSvObXQMBJUALiwfFweJVPLSRfdU4o2Iygf/LfjQ
+R/PyBxP+hErixTwh52p9JmeZyTkOGLD7P7vyf799KY5giHlF8PABJfHKlskd1FpjnazD+XG493m
uj3BB26G/vFGpPP+aPYrn7Xet+TD+1b8ouTd/G8YUHEB4A2VgWLHL84g6p9pv3p3MpSwezO847jj
q0j6IlfoZ6nAMqjkAPxt4CuD9QrFDZkVucQYqLc43XX506ChNL2rhdqz3pWIiQhXPZ41bH57tzpc
nfOibAzANy/LPcZ1xCcyzkdh/EVBFRDU4XTw4I2nZ2YAbQRH5h1znvF6WcDzKl4CxLBBeJtDlSU7
IZN5sEmCPdA5cLJjba1JmMzE+dpGZ/50fi36rgTesFdywhR9NxTCrrSFW2WBc/rD4kXF0y85DqFq
ykhmmhoM37OQZYzSeOdWFTMUX781sxJfUfrq9RdUk/dQXsr/PNTJbwUNVj4wH4airASue9o4uVvk
zTYYBNEaYF9lWuhDts/AWBwBcgNtUpMapj2E28ZanNVmRJar5g8wkFQHohe6d6psGJzduloNN4O5
S2MsoJ/wn4/VKZgObbpYJG0k7NmfjwcGNKB0aK509yEMYz09R09E7CWXdUNPWd+HvFg+aozeGcBz
Ol4QDmIslerQkdqYAcJl6IRi51Zd/IVrzXpIw+uBfP2PXMnGtevpa4aIIMc11XS+FaCxCECOrouz
/zEKbHCBHrPftXLtugxtMAU3PCIej6HytNSJWriwc9XB5GNsPdf+1ap25qWjVHTdfVTGrOzOunsy
oKjEDuPRTObdwQeE9fuZYLIW0bmqfrym+uMrka22Kv2xW9ct1/sgQfxZP00PriXAIFSnSOp0g57F
2454XttJzX8zeGfHqnTO1EhWqgT6g/zIxFDvldY6ZPIvTGf6Uk7qOfbKlmM/Z0t4smYc8NOpiP4r
OLuZSY0I+6prSINPMkX6yGAc4cjHL9cG0V7Zxlc90j328bU9pyvpsHicXwvliDtjWdpRvFSStou+
0h6MZ5F3/DE/PUVSbHGbQaFjhPtgBDKqfFHtaKYYIWUU8WBsW5V9scqbmDyFitnMIm0LWnVYUk/8
7lRipL8WTPXKaWrcQJrqx+70gErRU/x8w9pIXST8jklO/kbGuwh6mWfP2lEckYpmvSTkL6E/I8ho
HK4OlFIMYwZiRoT/vjEuBherQlfggei5PUsfv2o6y/UC5i6HU7GJP09kRodzyrrWswjjpCwXqBVH
mQ7+KO6BVXWG35l6iFwrtgxVbr67ULsQxVDAP8Ef+6DUUvsHa2meFyVMzV5sM4fekfhwf62HCzrW
1vviKeNWlwSDNhQejTWd5BuDZMJdoirHw1JpC0DwEo6NBBDUOREazBIy/JKt3CLRbMEIEjBdwtwx
90kV75M6gE+ben/Y6WcCImYQpS0dlHUW6Zto1NKmYle8hzrIK9kNMmVi4tN7hCBXLhF/KdjWTEpp
t7MCEnsWVcYzC9qbm2VokwXManZ5JTxfEkapyYRq8zOwTl/GRd672Nvg4Mvb8LNHEMZ8txMuW7MO
My09Sp66bQjQUo2/dB90Wj66CaRMmUIwAMzkdoowsrbRHhWqlG6YqMM2Ya7ua9xt4WPSo1z6qZNz
aCIqS6xcPrqgJkC20WJlTnqPQYoxzbLYutNpmWYU6NAJwJb4lrtpbSJgEOWgMJqrbhi9xVg5sBmS
u4tfJ4Rhyry/T+NR1uICDvy0ZwRQMelUqrq+CTKCCCUgK47gktrbhD8tVY3vwPrh91raOvxYV3qh
BY92mInK2ZkvnRpwtc53Q9bngDHZZhePW1mGHv+ZiKsv1vgCou5kqnoU6xkVAkD9ZUrx1GvaSZ2o
lCndC6DYENxigQhfrWbvVz9+7+u8Uu6qeZQ314M8zjs+rGmY+An0tYgjad+V5tCNljsIFYbXctBj
GSndOoTj1Q7f0YGWpwJAPyPyLn7hcuhmgMhJ2rxjw/mddaqFKsyMgKTf138ZbrmZSpYtpr2UadD5
2vGZphS1ZSdd+GyBk4ydywO93d10DVync7254dqUgFkD8YUmDFUKFgE/4X18spZKCnHofLRGgfKk
GG/e3dA2RBiwilMmGMuf8sVM1f61pEu32aFu0s11Sv38wGVJfNvHeu84XQUd/7yuutdN3Mp4fA0P
3nbJHO56KcsWBy7wmYC2ZYLGneV6j7NS/moPQS+yGnds/LYvDzRzBGISMCdSC+ufAITh8OS6+5Ib
s1HdWLP8OA1nD2HVaxfC34YMukgZRrTXbnEQkAn4Ul33Uw6jMY0mygKek/gmuTqPbNzjuBtXVelI
nguj21P4HiRCCl0U0Fvv3yG9y7wg0+zZO/njdSMWOXUg70anhrio+Fd1x8Jz+aqiAq0tMb2bfSB2
v2bwVM9I+MKpz1DgLllsW4NvS7DhqkbOWtFi6k4L9LD4fSXv3vRPiVsIk8iCv5gAn79TXKqJLHta
6JUGs8UgQNQTAR2k6rJ3Ty+xRqCOZ7yESDusMdP2bTMKh5z3ukTGLDcUqcF5X2xIsGgX7+p7fzEe
V3qiPlv4k28yCTzxVPak1f3u79hlTyWFN5VCn4cL4s9wajTqOd3Z4JppZXN3f0OFoG2oFaGjsii9
uMYDKUsE/MIQWqHyLjxgj3X0qi2ITqdcwHjPyibyctSyHH2MNeCZWXdbAg699nrFHw5h/vJTTd9z
FIUZIZgU1dGz2OWbXDW60BrsJ2FRVDGvMf+nVW+skmKAwRx0ZY3Y4gr44y0LZntoDC/zjohMWz0n
eu5uZGOXqEWNL0qATnuv68nLNSmQgS9r0jHzMbP//pUJD+0vj0ooQ6p2KeMl2+B3xdQoDhwblEhT
L4nQOCB8QgZJq/85JwmzM3WLpYTXQnxetuC5PX4f/lyQAywFMvyNt1ToHVIwoVFIyBohHrry0Ypj
WJ4WOFpyRAog1uAeMmkxvxmrsvdVGYPoPLNuuCaWqGYEyQViEVkOvB/Y3HrCkxZXBcRHXtCOPyfH
ZSazYHjqKLgYHRbMdB4RwB+vdSVCO0AcuILFF1rRQsB1ARWIsyv5H2ptvBNC3e9V1T5KoROfUFH7
Ue+MJhMApbBemzkyJ45n1+nFSq2P/mM1Xt9QRSaREPPyRtmnlib+0IEUpzOgh4gUm6sqVgnAUQLY
tH0Cs3ZD/DLyroCZ7UG6MsuxXnN2bz5+Aw1lcrukvXZ0SoyHR9n/dsV9qzeA4+jyF5pVD9n4nVQ8
E+9YaLF5IRE2PxJ17uy1UAy2Xil6U152B3EwOLm7orMlKLxqWIXf8qOXiD7ihIFiGOvxIgSWT8cz
iTYQUUzd70XrL45W/vU4hAiu16JzcuJHR/gNnGih3QecdhSzEONjtzPiErMUwL39++Ed9zSvkXDE
kV/sI0MFqGjpBuoSp+3xjPN1vaLQXd7r6Sde6MRnkBLU8nYj9V/xaPTLP6SpMVkDxXOa7eH29riU
doog5H+ZXZcV706VEhdgLMuJKN7mE0Svk2pIijAxk63y3mC7pDcYQxv1vzYD6qAx73KxgPh2i1UM
NXEBzQ8yNxQpK+OGFWHUPQmxoRdNwfdNPCabnH0GwNZaXMdz90CdZ8r7kew4ds2dVMwcWDzGFQAF
o1LeL4hb94ImTaY3BHk4YaPxkooilCowz9IAIUG4YA0Lovbt84wncGoGGW7pg5EybANPzrJn9vfQ
8ErpBpKKHAQN+coW9tQamInys0/kMaE2xd1VDEeIQKNbsXZCDpDlYj7azxqhDxQICZvrmxh8SkTd
GeKfw2b4suaJ13n9r5cRP6sYVspBUbz3+V46BfHAwXwaDVgZlOcChGJcYPJXBRyGHr4wRDsG8jbG
3uQYANxpVPt9w42h9VZJO8FdftVvNoIvvqHI4Jo1InHSwPpo3l7EZQi+e8gVV8SjcPTVVhWpC9mU
bHbK1yJOV8et9KtSgDq3Odv0yRRFKtgXeSDlD8vQ6HAUIxCVhNxd+5gAkYSK8i2GFX3lcqtCMlY6
yu/M8AMQpToHqMODHKbecO1rl3F3Cf3bfQnz41irI33xyV8iS1VqxYlAd7XFMAN/i//zSd7o9038
wDunehVRofjbqT7GkCi+uYmbZCdoZJY4Ilr3pHvZBo9gaGQtL8JMD1C0Pr+E25cZyB79ePefdJHv
G5NZ/UxFG52XoFPUCGglh+crKZ6O3ywDTEKX8XMAR+pCZOv6TsDDcHKjin8FcGpLtqo/kbHHZ85c
ruKJAqjQHcSmbZvqnHHcRh1qBUy8uheLqd333add//yJ9AZGJdR6dXxb3a9x5lQjylI9LHyXbZKY
F+jXPuqR3OuwQ1fMHEhrjJKzIfnbqVHQqNIgHhdQ8h61/Dib69wHafOaJjojn9sQHLyEl7P/IFkZ
ynkaD2OwybMrPj2XcxDogsmvDNjRd4hqJClK+3uJLhgL5yjRc+EgvrQtEljh0R9iCmHZsw6o2y5a
3QYhgBsbbkQvSD3VSEIgXA5OUVs2zoRAWCpTDCepUPoR62TrJJpnZVAlTuRL/1eXC52npI1T8Prj
HiyikRkzXTTZO/EIDvoVNoWXvcP7XbTO2eXKhIJk85/H7kHn1NpDb0GeTS8wSiF3UyGb/1poxE9h
B1bak6HYnsLH/8I39KaL2+t1luScXJYToNk5jv+VbZIwmXx4q8H4S5TUXJjPMdoByr+Vx9u4uy8e
qHmESnSGrdwieK2hcp8iv5REj4jDhgiatiY3PyTLNslUz1jEhx57gLFKEjhV+3jGVY0g0kr8Uhum
vXoXgZHMmdO20kleYgQOwTB7fzVBO2e/dqwPVW/JjJZMe/xXp28/2UkeM1on0wdz92fNSSU1g+Hq
FSMXlneTF/AXsoulcHP06p80zI6WRzzyvO+NTE2aHTmxaL7fg5eO/OIHBre/j55rIIiaUKYeztrp
7ZNDdc2Ilwop0O21WTm6ZHHt8fXakdqQL7h9t5j08RPvycNwwm0K+tZu7NwktjH4oXTMSLdHYUPq
DJCZccFcZdcs75yHZg//ZBVaRou+TO5zEHNmYlFWzj/0OcRH7TsNcGhKYW7lVbZ0cw0FCP4EbbHZ
5GWGJEpnhm5kc9sQX6j4AkZdjTij4L9m6HTbbBnOEUsmVTydudTnT0UFrZGtuJA4ngjb4HqAYJNn
Mlt6g5Lqf9anH7B3tRpFYZzbYBW88IU25Q4P10TUQaPXdf071QAzcQsXPkZSq5cRJ9d6rq3J1gxT
pkWoXNHRImQezg+du85AYyitQ2zb0V/Qar5P+QBU0f5u9gXFIcbJiqhJaxnV4iHmGxoqju9R10pt
QLUKw88MG4rzY/F1cKEV8q3lXi5fPI+sNTHjf52IfV0B3viQHflH837q5Zlu0o/fF0+pgRmBdtlE
ll3YyajPgYdmtqBceDCijpAA1UEaWNXORh+4Pe3YQPwZye1PuXGqC4JX32G2i+RQ9f7NEFs4SQD1
ShkXMjebV73Nr8K2570lxviUtM7BFjxwFRBBSQiQWgUSYQ9Z2l6vvgy6jpZ37S+c++TJKLePpDNX
EV670qgwC+Zl7o7Hrz5C0txp4F2+2zI+rL8m2Xt+FIeFqFz0IAidEvRjbLmP/BbpUF/NneQsgLQA
bciBZvCEpauDOslydkyaiDDeY5e1nEgNIfAUhIj7PBRq3SjceFsJ4Aa9eq7XaPl1ByKciNlnBDT1
u4PPsMU37PczeGhUMBrxSx0SgDGvtmQmWbsz2vxOEiqNOH2rx7DbaFhmoVb1PscK+fwJjWmMmcRE
/TIG8o8BTMVKlFqWHdTjPrk11qCB7BmYA3igbTIeVWss/TZCnqKs1mU8XJuf4BiE6trftZ5wfRwI
OKaXbsMjHJdBrnFKQRDFAcKpM8SrInO1P+oaVevckxxrZ6+8ORq2NbQmb4FYz9JmZd0LkW0MsOsS
MTHTu3dWBaDtI6SewgL6+wCJYG1f1tGyjWDm7r3BkZYYDa6FyN2ELWATsX8Ev67QpTwQKoZXHy11
oOI2uWrY/4knQjnv4oLnkaX70sSJTtNAes12C7OWLCy0OR+jPjCsVDpA9atCFVGTG/p51cnXRHf9
tR0CAPcPiMF0wBphoSaeYoUC8RMfV8sdOGMlNzYjMsUDXMzmnz9p3CzcfvwiTNMF0ZVFc6YEumO7
g29g6JBryhhueTSnbcITn1sTRV/xql1xHd/QWQ7lAxonNZzEIXI9nzjIMnlfZaCUFnAouisXrJZo
4d6bEKTlz+T8W9ASka9lXCGGveJUW6qzr4xwge2G0/D6zbctUbrEwYX2NU3r4K4UIsvRuXE8SIee
NhOaYcb4JlFwq/tietxUnZILoHah0yXecRLWDDfbJbzH8xlx1GboT20tZ+6PaaPQaozBGlZpNDU9
cjr5KZbqNshtd5EuKITtO7f3M1sGE7txWieeYmZdC/9p3MeWVv4So6pqwPk/fDDPLuxayEoba0s6
xT2wE1oPEsmh9+IpM9UFnrRWfugFIzG2gP6A0sF6uOJogLp0hL66PoERZPOd+B1VS/Y0pColNLZu
EQHYPSfA6ZW5kxcojn08sqpxGMebpF1EWQz2UbFZoRQFZNa9riyZQ5kWaBlEigih782ldD4CIc9w
H7fiNE+cG8s0UR3mt46kCioQeJ3i9PW+vpHbUy3ArKhq93xBJanDx+t/7CVXdYG3qGHUd2+wzE+W
J0nJZ0bd7tuSg8yPwvzsKQmDDdt65h3bQwt6pqwRjnrevS4oMNsY03Ivd2DRSf8qus+jFecq+a8g
joPF2PjXe7AkvXcVFg1BLDOb6B7r1OY0+/ituPtkmQVMJ2Wo5mEcJzSvxGFXx/F58BdiYzVf7h5v
FGZA9s481OzmKZ45ZL823op658otKPFG9DZ5RZebFBgsWscu6kseQRRUr2TC//PyS9io4VnR/XcM
HjxT3uV/IgwSwfZBwxosD/f1LRdhX0PTaXrwdgUfmY7pwej1twSeEwGP2sQag6Ax+/fzM5f+U2ev
42bMjN7kRtSJKX7eyOH036R5mb03NMdwz8FmRT7HjHeMiYwXYKw28wRN5fgpYEBzDFFaMQ8eyXz5
qz0xfFebUpC9Bluj/5nzUbGxAvByyk3jK8hUk+j0HL0i14Gcr/++zRYdf4+r1W6pl60eDK0VQyLB
ncr9MbeGE/KyQKKSy4fRseMFCkLnwRwyvFLCjVfDlF5cevhfE2YRpgtDSx2HmqbzgImETASWrmXl
O/ebZzdMngkcQ1SwziHjSGQFn0WBQcNb9BKe6KQdt15F4r6xu97t1AKxAagGEQrqw/885x+07+fF
2c0OYmXcCZBJcWjAkz7vkD46S5xmLollOTvOZeJjpEgKZCEhlmuOHKQxznj1z2q1BRt+06v3tZ1b
Yx0ufbKDLSFkxYj+QjNAp6alPI7BLRgS1R4Cxmgwc43Vos6YzqgBrC+4HUbOT19BiykuzucGdDAP
waybMRhIqOBPISHsVIBToB8BbSzHtYf6HeFeHl+LaKFsio1j1n+8S3G/CsgrrgjwMWHRKgP3qnyt
SMeFI0MLXatnv2dY9jdQ3/UwS14IaGuILRtmSlf/wgEvmyeWnI1z64KT5pduQgPkmEjdBKMIHqNA
potdexPKEWxx/x1CSvTemWItvyylWrhoMRo7mba0XHWwRA1E9wxsb7Q51SbtsLqrjbIJ7Zq2L02M
M8ekddCcrx8/3cZuCi6KisZWOe4CM+WwgM7+d0sRYOh3EXXTMp+G0r9hE9S+q4muCmHF4nR86fJD
wFDtIND1gQ4wU95Jxv0Cb/HmeFI36Kz1t0VHCGEgKhyKt2BzXrcLTZjhp0CTKdvmkVO5mErEPH3e
75C3pltRVCh5yK83fXhAl9x3qQJRMksvLp6lcIowMPpzM9GdmasPpmcIewjrWH6CfohM3k6lIvkq
XujCrQ1BgjgobWkYIKY2tgiyiMOzKMhBVxYdF6grPTiDEVC9q5Guvf0hTID3SR2dfdLZdxidpbXe
vyJuuyBTTtjW+AdngH2skJgh0bTMIV5ayCywwdgepIfvac1CkqDlkEY0IFyWyAj6GVTfCm43bw/y
Jgq4kYO6rhliDHsaaPTNDikPdTUL2J1FU4VFQUnB1+N5y/+BxtRNRUtM9bgtjE1wVfUKrRBwdrBZ
AiPQLIePa5AdU53ufuwZ75kPOLst8g73H70vV1Sd1BLfc4dgdna/jDNBP+6V12qbHKCMvzdsZooe
f+vsXzCz4M9fq++zq7ylfhgKAsQoL7K99fu5HZtWUZhyorHtftkF8LEaW4AKwReWGWzjVGUHtcQc
F+l6rl4rkZlHiQ2m8o31kLAYvrMKH82YdxC+nA/iLFgbw51Ii0lMX04sUZV0fvk2gAp9QZamYvv4
JDODkoO9mjuEisArNT9rkiDVWeJFSFgCXZLqnYVpxxIblZXU2JU3fJP+Wv3E0yJvJyWYYLWiKU0M
1WngFR9zIMVC4+KWIISXLlyQ+QuKv6jW3jeuLahFZL4g4E6/HLPzZWVprwrgEmD9ltDwv8ZbHUec
pbItr99tYTV//oltYtrXTRxE/FrFmvBfk9/X4545oYg4SRguvQKkhCCXEutEglrcCfwHWQH7zL7J
4Sljom/gAyMwT2EjEuxf24BQB0ISEtyZZJwOowja2JK5ZfAZyV+NQbF3H7tHlGBOR1ACa/jGElnb
UCIWC6AOEbT+hv09k5yqR8l6+bPPi99pHWympGa0E6hvPIeCV8aRhCtsR2O9HutxPxPhiE6Zht5T
cNSCU3YDr5ko6qpgMDQpwWOS16PMWeU5wlIEyIaMmZ1TBaanVB3e6wXaAYEV1ywELNcVaQpSb+/k
Xwmcvzifo4SBPNlcPjbBYirccl940uMJ+GXz4sju3+6KppzyLxqWArrVPPZw429W2YCzoRYCm/Xc
4pExF33CBonxB0iQle5tZ6BC4bZy0YKviI+YDZ7iTUIUYztVbySuwGsGEb5c6aLZbE3SQ7OB1pqo
k/AjeFI1Nq4fTSgdZ0IE1s33v0ldo33FOtrNb3HlyRyzGFTgNWA3VYo+qA/3ih6Hy9mTM9xZhp+f
YvOVZ7KywCka99g9b7P5YfjbjogUr64d8RbF1xASXaAYsqX+YeEtu0LkYXO6kYSTsbiH1EzgTXgT
3VMfzTE24KJcYbylLYjlDE7o6trcyEM9snQDWhzNW1xNdngQmhsefTlChbtp/zxaYsaKgaw6iuiE
DuXAjqn9i0dEdRTmH3YdBLLI32X4hjLCE9qZVS+noIitjG0Vm33xbE7+pMsoWT7aZ+BXQDxmT9jJ
06YtOfxzxHlVfboKRQfq14aZMi3cOjG1qMmDjy/nUkdtTZyaBD+Yr7MK0jZE/5NaLyvb4qiK424y
F611IZu8zFu8nmtMgB35o9uYnJ90fg5gks3xS/4Xlkd7ryVBBvv/MuklTasJ1g9fLdSB6LuPleW+
JqZE8nDP96mHCrIlk7tKUkpGZJ5rg9Iwoo6Bm3pfhLiW0m75vvsk8jaz8BsTvjSLnDfvogPKYG3H
YoVfDfNcVtI5YdD6V34ipBqAafVxKj96eQybc3/keVoAs0wril3lU+4ZsXmjhjcVR9NvaPS2ZAOL
nilXTuIJLZQ9jutyOnM87duwPd3855onTy7+DtNqAsir/yHs4QR3IUAEkMMW3bIOlolLmV+Hfb2L
SGz2oswODTg4O8pDzoKyPVW407N4SmSp9IBdk4dQGyYX9X2ZRobH/mP0f1s+wTgJVZ6Y2a0ezvIB
pEISDV261tZTZvjV/35L1L+p9uCdUD62terF9c0oQjTBqTy7vzBwKQ1rrlzrTMydYfg+ZeYxBeWY
ebGrfdu4FJBi7h/adoOzu1FbrXkvtscFQs6pGFskNpLo/eGRzLa2o0rVhjsE1JF31w7SWkuNjVv9
59kiWUfa5P4adG0w8fp5LCUUD1/H9v+md/g45y6MlG84dLoLMvGnlwWTr7COZplAzJZ8nqMDfnCe
+MZGEwShAUbBWMWw+H0LNhjjkwmBT84niWukVUFmBiGFfQ37t0qNgCx7onEHqAQwDqvzOB4rYTwS
ZVT5sKwc1w31I05mRS+eWm8/a0QbqimzaLaCJsJfJ4Spa1MqC7IPDVAqJYJEghdXW6RJBCI0eGN3
VKUu+YNgF1RFYLAmbnn/kocpHxGANtDoyikv5sNlQA/GSpNWTWBudNyutiI1IDNmuC/YsMNIO1YD
MYHkEgPCyAsO3+Uo6pgT0nRcbGj/L4uKxMMZ9jVZd7LZzfh4urBUnSrDQjW/grXHbSDu9CvhZm1A
TmiIDGkc/9ztgPvQVIRegyC9EvUmpxOpi0toyuxIc5+H7m4ZUJPhDsgHNSKPhtP9uUizXU6TNONg
l5pDV/7HStjdrLF959JHPFKG8CMAuT6DZk0NE8luZuWhZFnoADzNCLK3EdBClVtAKJlvq0NezheO
Okg5ozQ/nLAAC0KGutWPesCcPi1GzRasS1Pg8ose3hY+ezv+mjAbv5b+pqhdZ60LvdQQCEOmc4Wq
2YRwxqPAOFJuPiNgnSIaVDwp6Ohy9tvctIFAA66UVz5yujOW9e2H9kSLnIlQtqniS01DRh8h9rex
InNBfnMMFBUdgc9aBMsxHH9ANL+44K8/ODT4UNwBLHQQ4lih03hOJ9pdEkCCO5mNd7ed9gF5TrFx
kVXmbr2aCop5rYj1prVHTCf8OPMS+B4mQShETWWMB3SvWRywT3GpcP8RvfD1zuWtEdQu+hBXlLVB
afRvmIen5KDBpArpmHkmYYBUlIqdUutuqGd4prTTzSdkfzYADRirXpOmf/0aAEEygD2ARWcfv3om
+I5+MRxu0qpcjmr+aUKN8raEhxuKrXXP2yqQ909T11x17r3Nk+S+vLH/ylEGmr+YopyTKHMBPZ4P
cbn7W/X3fCutAQFtMMzcqzH+cbVJ4m3pnw2yNVlErHok0IeT+Z7gZLjaIkQ6NZWDQjCpPovSLSNI
JoZ2uS3fa6mKeXdthHDl72FQ5suARI2uWejiK4SaEdvP+vlNNu7F9THKik2Ql1RILBGxNAViGsJh
22+/mSzpd+qWm6cdSdIMs3IpVhjPrrlfYv1E7DtgtB1GTbcJUUHMz6l71ZQAlsQgCKJUeAh161n7
NQg/YhizQjJWuHTKlOHWWhXqEJqv6nbIAFUv7OAdEyofMHRVQIyQQnaCwNkvBfAY/CdurxKdFyER
UZWCT9AYvMVZXBGqnjz6VJwW7nTrzopR1gfSZqREM/FInIeVq4DIOKmjLEC23yfcBk2zesiPfFgX
Uh4Cu1FVTn5bgrErj5mIrn5vmfPyYJa7X2Mz2hPhZVrPVLTXtb8PGEN3CVgw9EquW/8JwCIXKZF3
VTEAdJEzbgNjqos1YnaQMEIUyNyh65bNgcPvZWGJsw0UR8WdUtrJKwps39jLHz6grK3Pxv4NO6mE
khDmW6FmMyzJiiWpYbdSYAuyGqwDDw3m0XyZHZ/0LpN1t4LrGXgbUbJKLP/nukK0gHqevs9BOM/I
xCTc+yDBhczU41KQQcdYIIYCfncr62gW35PD+UQtMIQWpN0OhwlUpsOlTMz5XDMvC2+cF5GTkcRx
LZQCdNhnPDtm4PtpIN9Ee5uUk7aCuQ8rnugEswxX35c/Rm9nO64kp8UN2V37e5LlMelas0Qw/ATC
zO1vd8YhdWB0lQHsnjpi4JJT9u/FBWdsBB4TJFIlUXGtnmJoV3XBhDBGXd2hkBYKFJYNBmpQdk9J
FmHM4wK6oXYo941E4UGfNvdrRuNol4Vr/q0+/Hzuy+ZOAGded6t4qAlFJkrpUGy3zGgd2zBAXWDT
aqVBxGFHroisucq4WaXseeRhsddBzUCJk0dGSCmx8eASiPQrQ9T5m6rb91kE/v8QHHR3CWhsBddm
LKTHFBMNuQRLJVuQrkMK+bl27QYKACUcnz29s4v3E+1ZRmFHwo8wrNMMKMwUBx02MtgzDVEImNc1
jZCCJ5DCm1ApP2kD2CLCtAPwLi2yZm9LhaOdENRtusbzqGAgvCj4stXrtNw5VsJu2Oqztui3O7Qa
vMAO8DIMFmCxYD7UZFRWnZanQw1XhNrEnb3ATl2UaSwzdbiiv5FGIb1/ec9AulPsCSUx8i9cexEM
eYCcaQjEN9bX3g1Bz90K4QqVfCvEUJaEhUrmdypdEo8M6ySQGX6v/QHA5ITGyV94EZFkyUu4GvPx
rDK3RvTvh8OWu5eiARptEkDfw1AmB/0lYgDcbmWHuud8Riw2owaU2QNun5lQAc/dTstuaSIw8woL
flRN2WtfHNGL9iXO44SzdQF8BU4WKH7O/wg4OHyFa8/F8Zc0ztMpChSXPb9rwREWhRxynXwaJ+Uf
dAHLNXgXHDEHfxJYESSijODFrLCFSuozajLhSKGCBgFd+gLuX9/gnC5gkTZMhYO+Y/Klr9i6Omic
tMub80xQGBmI7xTWwyZDG+SU7dcemaimV1PKk1NsbbPNsAIGduSzO0QNvN80jjzdjSfdZfNDzi4h
OXERFW/nf5+t3h7FLRhZZKHACWD+KwI0jKW1i/+iZdcCJSzLYLKPUDo9V2t1/gsHu8iIA7dE3spj
7G51gsh6Nc+MyEOO8nyK9pkIgSOgWzd9h9ngefg8RVrD77gyNXIVSeNFi61QfmLXJWgYu2Oa1zsP
11vz6IO88bXKKbRkNFJy6QDa7cQCWR0Y/j7Dg5EXULVYbhPYkI42DzFSvb7j9Ukp5H/5wvPL6uNN
d0RxPxRKJw/tdq5tUbkZIDYN2FD2YcXrIdRRYmrA2VqeX0RIFezjWxvcPx5+Gupjr/NqD8YxXejk
GGdxzHNofKlhNQNEPPhgMW1x5+Pfde0YUSqpzIvhK03vpEQf0jsi4zKzMZAa6ffhukHuVpttF23k
foFxHPl8PiO4ttW4/ckRuUKuhbbr5xp5DMMwv1B9Zrnkv3n+qYH7MnFgkB8c621bcgBpEewt6zVe
qGHN6pHWJdaWHSsj/S+bGNtrNia8cHrAlXi4Ywq8WpW61TMItiNmJwPBXkxuV+mGImCx7wxVEl1f
mGOE7cooSbLq4ThqhS3Scbv0LssBWW8O49id8Oa6+gTAcXJcDsd6gyPB2rDSUTmcQjFjc01s2TtS
xRkTyCi75cCQkpY0tQ46FrF8XuDLKSIJpJ+kK9gK9bYnTTsiih7XXkCBUC231qwiwmZGpKSW4+BR
e+2bpevp3zk8bvMwA42oXn1YFSeivMcVxSgslSqUah5TP6bFU/lrFkomUaRl2+Ii6iT72ejqAcPL
rQSZu81c4A9moQb9YgaZWkXq7avLQpb/0a8lgp3nabWe3R2X22yxvh8FyDafndCAd9UhLMIW/nne
S4xlLL2M2TLVWJgT7IqCB4Hw5zr1ryrCLp7H1lovrTe/Z+T+XWvIjjspS9tL86CCANoLxMH/97Br
+WRlyMO4R2Dxg21myE7ePxIc3ieoPbaFT8pzQt7jjyjFVc7hndL6Cd3TGjokNzB9+GgMgh9s1GUe
ytb7+xkLv749WBjZAFET+7+vPJuMMBscbYELgxiCYouAnTHQtuKKvvY5fCPHktYNpkCmB8Wi/bCS
jALHzGOaCwgtULwHyGi8ZsOQhmD6zdzozYxD6F8j6F5D9bgP++tx++q+1TXSvXiW/NDMV081gcpE
T9AbU3RwV5awfnEa5pjeuaBUQ57sB2dic9bhyyluQnYRJbXqVEJbBUAlVeCtRYGSgFZriuGNFkR1
cNm2/VbOpMQ5H3fMsGO8gM9dhWIDLxwy5KgWr7Hgppic6RCmbq2iTf5blzgxqKUhH02qci2Wv3jy
tHs2JiagHAnOmoKxUNvhAfcnnshSahDDD2/2txVlpJa22zSVJrKSHsGx6u45z9drERVBdFtIhUSD
5a9TrbPxjKOShv/u/SFZr9+amGheksuxp7pgKo12m/Cq0ycRvHWs6xhgoSVnh+x/Pi10L2NJj5Hi
y8bv7eorsG+Sq1tAZ7oEZMqR4/FwGP4oJvJ0VU3M/9Rb2ADCuGz2wa2XyZYrSwwL3xHrtuFLsA1p
iCSINxwsnbK8EdgrT77TBSfjs4Y9e/JfF5b6hF2zN4VrElUx+0fMjdkj5eKEv1cfKSbQewj65eLZ
d8N3+RYC3yNWG32iJjl/kecQdkdxRLARZiEpN++oYSlaGA6vE+EPTRGDzpilitzEvUpsy9qfIJtg
j34U6CpJeOsrCPCAxHIKsWftIylJvTXusXwhqbC3fS/tJTS5N3LlHYsIOnqNvfq9/IjQsLZargTW
bC58v+DP/itEO9JqR60+9Un12kiQovK8YMOHGbWGAbklVl3JiQeL7R5DYDJEWYQF0doxXWMSPj98
ZfLkutaTxj7VIYOwfWvsDbCdFWChzIb3LLXBFErrnq8uKS5NJwdndf7BCDsOM+pmUp60kl15xVYe
kdubDQDg2amu30Q9inSksBeuCNK+3s9K+1zrzKKxLmjCdQNjy+ACLAzSYrdkzDtKcMFA0Jlmo++B
cAkzhI+/6F7SeMXxirTOI/j8Zaqz3GNN+Nld1vKvrZo6/aDD8wY89WuIyWj+Z+tmuwTa1lrERWTk
0+zmxi9MdP3u4YGMErkvSRDT6lq3Lgw9T4DVmEFOV5Xq6YTk/75yeYUZeXrUcltRCzD9HoRjpmFv
ZYe2ozqgjZnm0d5xKhF8vf6/xKyMfv/KiXLGNFI9OI5JP5XU8oTXHRka2/IXkTNUTWq7pQKccEdy
TiYjvMUTO/DWHvMwokejBqMX1uPpa3P5W7ikvop3ey5l9ZqrVvEPkPOpGgaxUQWXsjaHP6uFf+08
TPIdOMEIS0b7nNWtEZBrTi79GBnTHS4gX3auHS/pLOVkkxtQVuS6iv3UnmZhTJwdhz0mtkD/K4Gk
9gT/zoRSrVgv4GVthppz8xrLRrNPSJX3GwqHM0iPGKxmLpgk5znNbZ02jpdKZlYLfMyQ9EiNMSHj
buX3QA3CbIlYnSVJjgsUOOGliPomCalvLXE7adVinJTJ6GPTmljrPTA1ttj73EvtQvhSu2wATGqG
e4UBpgVv5ohXAbS9TQ3asBrXW5hKxp4k1hDpo3HDp0+xH6c74AhlhJla4rThl+Yb1S5Srv2BuOrq
kDxZSK2cnpDgNZRiO7/bts+6MIokFckhx4zCTnhy8LWcHSqs7Qc2y2XJ+J/0jcx+fUhLLFAcaq1y
9Q4tdyky8wOlOeJzpKzRuJOIKnyiCUocO/WjbFlLrE+rj8Gv25zHHWoawDHpkdYhemyyBU+exLGK
rjS/G5lEiEXhA++MWABozvkjwKu/kSbfJiOG/ZdtBWr3zk6auINkar1yLYVq+DxkE60/yHMvxBxR
OjAAJsV4LzTZw8bhumSAUFyKNhxSKx30quilUm2IAYeX96ynNe+AcEMwSAD9NTxk3CXkMl6FCKdd
C1ks4Nj1VcTcgVlwfUrFZywCA49ivIYdFV5zMYkpBVf4Gb9fwiqbA5k58y2ccydi0bij0cmPI/54
2Q6wCPezqlubA9ktAyLYA83N9xYgQDwUwubfytX9rsmLrC2B3GsYDwouLVJbL8XJ0U+kpvJvBLIP
Ez/ViASNvUEjeznDzhTiXb50xildhwF6eNqbzada7WAOICFZiM80EjW4tuE2GT2rR3d+HKJo1OZB
vM3z28sLtx7xeIV+xJ+7/Zmdc05fXAJZTWq6T2TG5f9M5oSS8Y4rwUiR7ccg7+a/k67VoD/w0xz3
5wmiLBaNHuj6IJGmBYxXfb1melHqJrNDuMWznih553b+onJBUFP2uCoXqcjjGg896pWHCw5oJPL1
CU8sZrV2cAeSO5KSotQMp1TBixalTp1i4Fpf5FaP8DKmdUq5twOWDIEW+DB06p1fWyWlEaGsy7ES
rAKWEokmuUgmpXCcjQaDBcBs5YhEVB/k1kI6jFNSavSPrDFNEs+Af5QP7YUeT5VfMzKhvDroR3H6
bievzYix75X+yLSqDC/jbuKJAwOGG1qvIZ0JY3wIG8ueJYZBr8oikyYUl4tZ6Z1xYSvtsVX9nBNl
YMXZu/+7q9kbpOVPEbYqi7us4L/C5N1FKzPYH7yJeIUh2ktb6Ya34fA6MiKbFUhEHuO8/0sJcXEk
dnF41h06Or02jK7UwpiZg3YQbJggkdsBOZIRVn6jat+pwpU+GQFY98jCKSuDeZtbXjccnRMTFFHT
PbG5s2B9VQ/K1f5gJzN57NwB8b8MifHRJek9ur1PoVyC7GMIuSuNlVlA/E4ldGKi9EPuepX+0M8J
jZl1yYiSqYfoxk0RNuwmtaSv3ei19de5fo9Ql3PGwpryrxZ5m9JaTElKi0iFzl+Q2+vHYjPNsPYp
JTJwENr18yYINN/j+r7nczfVfF050Zs/OR2dSqkW1ebs6PqHXeDrFIzpZreGM6VFOvIuPYI3LaZl
pedj/Ymee0KUJ/z4XU6MRvTWI2PTBiyCZd1K+C/MHtgrLeRaiJVQKGlTaKVX1lPnC2xDZlb0pl2V
Y4yRI77haSFnEpIDsF2ujO/ETiUWGSP5XsLn8XS79CO/zS4QGDw4/EyEghIu6LccgJjxOtCDK0SL
kSdWgfWIvTX/3Z26n90QSrnVOgNtQqPajWMnDDZOl2NMUUaDVMklukd3m0HMpV9zolX/vrlf9dQc
eqXutWHtmUA48OQAkFYPM5cPT4D6T1w7SQF8Xj639U94giIkUjoFD/gVxngjqmGRRUoSNLd8ZWyY
AHmjR0e9zbG53sS3wvB1S50fB6pmOBKON9mZxR+4kk8QY2Q8yuW0l2pKzGmABfi+WiU2f8zxdaTS
gcUioKJQUnrCbabiy8MFWI7sU0QfzD359A4SlmhX3h1/WH4I77TQaR9D400MVxMftulXEr6Knqm4
WCZIuXb8YU2QMhk4V5wzAIHJqHazJSJJD+mWf1fOdJZcFvyN/5PxH+8nM5cY7x8qRheOrC4oEKJk
4FVyD4IE1//zG41AONcAsVSOU2QnY9+dQ7K5Flbuq1DOv+QMYKZL2sjxxxNEzgyCkP8Xyr0wvC0m
DXDubb21SSmFUI5HmoBrdebS6210GvoeZ755jyTYtAOC7bqwI33prk9DvFLz8rxRhOyTAqjMpI9c
SLdHCwZIwI2lcpHl0IVKgDv2rLbjrVLlnbumdLbXfBQmRKLBb3z4+R0p8fJCNkmw+sT4SRJ3YryP
t4ARRMa3Sm1vORFtJwcwIRBAk1EhOa22IJIcXU9Syg0zXOYgvJVijjIKxz60Xh2BZYgVCQ2NS3NP
ONvLQ/w2LwoRqv5AaK11z2BkKFdQvfJPtC7xYNINocnqe5jklWiB3P/TN2FLoz3sEFt+XOoivVvw
7oWwL163mPEWqBMApXFLBvNYsVT1YNX4w+UsWhtCQOdabgR/CmpJiGkJ/g9gDkQzXWxr1b2Zr7JZ
vAxld4NPLNedd5cHPat7CFIG7k+YNP11ofuVLnqQAkNmjHY1+XKBh0+r6WXHmQtL2frqTCjxZUmA
of5pQYTFeW9wDwgETlNkImmX4VLRS3fIEEaGZvEGpoq6A9KITlH1kGvtJC5/BA7togFdsxkU3Ek9
vtaxpZki91tF5QRGEKX2JRLPvTspicrXo7XQZLqTh5mCBr7X9B9g/7CQZpMSZCkrj+AQ3KcGO0YB
3BiHC22KxYdFbTJ3o4vU3VaR0tRSATId7cvxMUznXAaO3qkf+K28xa/AVzbprWSuaCz/RbVrl5P6
Cv2ke+A0Im6WzH2RtmLVpycCsugFcLfPZR//T2xczc9MaI+HxItpitraVYnyoLAEEbPwpODiAK+3
Swp7n/nlHeBSZWB4w2W9YwxpBWk1hm+fTk1oUYQMA/YxHgTNUftXg0gpkSmtjN5z6+kJDCScYwa2
j3RPm6oDeMts/sj0AcZVnMaDAYHSP2B86PCG65vSg/0kY1uO9ruWSK4tpJ3YeyyJSLhyHW4FYlWE
GSmfLLCGjRc1n9fIztWyV8mNDRFkuYT72620w+WSrhMLbCgRIoOBnX7f2CDe4HXijN7rECCCMykk
+thHQew9LPA2CCzDwrx7FzkaPWdS0+yYPQ/pxxkC6ZuvIFl2DiMsV7dRWKuzJbByxoUP22KZ+ZUA
LzIDACDclyJpwXzkl1SBseq8EMzvqJNcFlPE0TYykMNTFsYmLLp00m3DJDdMGP6zXhWClUb81Khh
NY4I5KdrZ3bFnNk9H+CCZ9Xu2DK4qsLrG5ERD7lzD2paYJ+0q9Twy2WkW4K8/4Clf0fE4Tuteq4J
C7z51IyhmwIA45r689LLzEHwcPvQGhYPL5aaWU7svntegOW4xINPe03tI595cOlgCWFl9izonH8w
kci+rJPIH7LOG5uJkyR45nQHAe0JkxeZXFjnKj3jlpKT7Zzjz0rxvTQbd2lCpH6d8hKiRirvOUrt
CBZXXVQPVpOzj+EokzlCxqSbSICylmC/DztU1PfKtk0C16I2+EzPe4X5AL3OABwITMePdMhppsul
bjbzEmTNpAxO0H1y5zV5JYPyzGA0gQwzqKz16Cm+CSxKicz8RnioILPcAg1xFZocKHatmv9KNi20
22XPgsSAdv+Vh4rT/KKLYN3qojBTYyaVp3NF/5unlcvbcrkOj6VgjbrrAtAHzbfXlEXReTleawNx
AQynfInQ6X1tXRq8Om/wR0r0MjzTc1mIzUS9L62puJ1c+q5EDD1FfXbDo7q6sl3KHOx31dq5ZfzS
6xsrVfGdMisBAYh4h8sW1fB7ymimiu46S8mXU6SyEsh8LSQbT9pKqIVLK8iNpxcdNCLPFzkgUuLh
Tz16niYWQA7sOpM6ebdPgCC9NslSvjlfLSDjFiSkf1WU9nsP5qz5tFy1XHdbWfkgQJEVydcpZXbB
fq32XY4OhvkBiWkdDmPERedNOPgsa2TeQOsNCHOt1AJMGbptF0DWfRcfqDNjm9WnBQYuZ54xLgtv
K9jDFgGfeMimf3WuS3o1selsIW2qJ3+cqcz4s5OvypJumteSpkMSSi8nQHqZd9wF0UTmOhfovc+C
CGJOYJwBeu8/PX9/2Zm/R4JmYJrJGmfaRNaywoTkeKbWPvseBwCbKgV6IybAeEFXs9oq3NURa7On
DHtLy5SrSlH7mttj3KoNcKo7BigcT4qOz3w4c3P+AomLwupDag6lEiWGxofrjXhq2sPbk8Lqv53t
HEA6Ht6mO8GZN0wPP0VpwuJrUfIU49jkOvbIf0NBEuJhJ1KvcgwYHLJT/JGa1YN0aGb1ESNZ70n/
Ai0eSF2+4YBtpxHfOzx27Lmsrua3/hK1FMmAWaXZe7I8YOsnTHBHpqjKjLFO0dazp52Z2k6rYW9T
HlD6GWe9/IvlKUqa5YoelSCEEMPog9rH5twK4/qB7AtEsOmTCNAbLYXFfK3tAYk2Dos5Vc1ieDhC
ergZad/m84tFLIjuYO2NFFmZl55vYYdqbkSZxBj+25RdECGnQ//PirCwmzQGpuvdfsrkGHoTW6aG
R0NjttJFzQ507Gql+tkSY5g9BjhPEAq7VCP8vzVCYV/BXBP/gNCPGvpBsMUCpCV8V9nMHWVT4i5o
qdj36YYQ0GkxkGEVF7YDJ3HGyLg9ReU8qTlAN1GWqhhkwktvgT6SZCsPyI4LGUPFlZqjL67U4nFe
U1COU/6weRGr7mr5IHg/KzDN4hTu3eGiEjBQ17RY171O1FDJKBS/lqdzaejGIRXty8ewiXn4iF0r
R9+v03hWiQEXhyg0YWG3GJyI60ZEYWvocNLl0JPFkuYMC6nhhOLh1NMiaa1sydkyt3mCd9qKdIO1
qYmRHSSA8C3Udu257he/8TmYM8uUY5BFG6ABSeHR9f0dCghrJnmElfWiEVXOjPDCojTCKJipsFyc
qVvhfvcsBLb9x0r59NnVhxov6ML62hTCWgU30DnCjqeVCBpPnfCxYIBtD+iZNFymaJzj9Vtwr25o
iSEv1LLyIgEHJ6x0F60dLMa+ZD19w37PZTRWT50fHE6koFOWCYvEZ9mzd9JjMO70w24f84RMWiDy
YoEoZBjVFZTFB4N9P0bT/ePTTjyw26RCO4b9gDLe6kUQL4IXVD+eG+u6GeAE8q2pRIkrRT50hAdQ
rHUyYgXiJXjkvoLPT1oNSU9Evc89QcJtmdCR0kf9/l/LguXOe+c//wnCoOznEsroV1iRiwvjwUfi
R1q7C3IbDfdaDqNdZG/MY7088jr9fwC+TiXh+z0z/Pyzo1SeFJp6gFVRFzBxTAi/fFqgCmLtvFRY
O2ef+9tSHokFv8iZMsewb5VeARQybHvE8/r76MP1Vga0ZpT5hfn61HgPoO7HbaFkMslQctOueNWb
3DsjDshyQW2dKuXRJuIfVKNjoaOkh5QrmSCsHOybGJX57//7YFMoxDMmPd4wu9W32dPFdQZBah39
JP7aLuawcxongqaqtqRihlntVAxqPHQ0hOHB6tRQU3r1ED2syOulrvTO+rDvfPH37tp0NeRSBpTx
RFdLeln8qlK4CtHtZH9nOGaP3vFACAzqp7qyWOyuS4vuk25YCdl6nB1vwm1WR0FkIsX3FxzY//mn
TKJLzX4aH5Wv9Zr0C7rZYO2eQpF6QMfL4XTz+pRpKEwQsDCZdsTKr5eD7zHBamUjWIIuYwyz5SR+
cXqAEyZo9Cfy9QfSvQcu6CJow0y7f8FbX0OeCan4J6oz1Mn0XJEWxEipf/eARohY1/GW7btuCExO
lsmnxKa7N2ZAQBylMWGizsejnDuD3dMJlCHjycm8CgIfUWmrUQdG6bWLMvXD/KtnMJp4J8/OwkqA
CtfIJSzMNgVdeGNzQDj4H/vdJiE5kL+VGg/J491tqClJTySimP5ZcvEVRZB8rKAfKKJB5XtEvvjH
Q3gTeNXiYr6tHmqE0ATHeHBhkpxfmUYJCDvqVtQWaachw6+FqkpYmb8nZQUd4TawQKS+SxMQO62q
IvyXxlubOD3Fw9LmRaJwUTl/tBU4up4S4b2THQ9QuTu3dRaA39UmtWIdJYHSZxWj8qil66cY5wUg
4ocZq34rVU1H5D1N0+yWIlddBPUpQiHlKJPuMppyZNpSY3psn3ooWWittiy/JjprMEXpngaXc5ef
/vKVVaosGUkhnC58DghNuFLfMHfnj92Y+sPb+l30lWYQmqoNJOTc0vOiO1jgzU8pDr+9D9HK0IiD
P9QAXF1w0ZQuCIMDF20N79aIImmF68GJzzoKpEzFTNvovLPogiu4DHUIlyamKoTi5G2aIhJjhuo3
bRwxis5dq/LKO/heeD9+CGOvosR6frN9N0M0/mxw+1MPZvyH2RvvIT3Xa0P0B11vgeyZzj2S1HIT
QvNcIZHDRQtCQQAM3uv31WNphB/TuazjX2MnVGx2xAwcrTO5APdJs9SymWqtg80TpDd3xs/KYVQl
Nn/Bi/q59PG4QlhFGGbx7HxnuIv69NtY6EPG3BLqOmGLItHWXIvq5LWvBJyu8dRvMEgO9X0CHg/E
i6HtGZmneGbGpWCttSBQNyjNNTmGhS7LYYbZD5EpLFn5lIVztr2rCNd1NVdCV2+X2c4n10G/GDgA
TolOcMdsvWi5Ay8nooB12SX7n/f8qg8N17ov1vjS0C3bCO2oewgGPbgKJxFK/TvufhcdMVNyQFds
5lhRMNvhk2DycxNIPSoIfY1HPMYl/pPZORyK4uDITUuQayDkU9sqPYzDWk5I8wdd2LpowWekpFj4
NBpXv561It6EXSd8cnduyhhTjOHphLczjoPQ98T6cg0GlrFtIvDZyYEEFVethXnOAxqvs7pxhog4
JnbX4xnQryJ01l4h8r9dfgne0aHODWb9XYF+XZ4iUgJgu5d7W/Pc7PQkpuJ1nOk5aKCvbaX/jS+4
XOEFhOsk93UyPKnUYWmEkNoLiG88l0TMjxqVmqv04Bi1BT/c8v8C0zvygXpAjaMKvlbyOyXrLDNp
U0T29eeOSjnnusjk9o2V+6VoipxF+K6A5YdIjUvMcHd9crrocfizRNJBeqd4z0mwy6Big4DEiHDE
zcJIht1i3e0M17/YgaEnDvNSds8EPFcEnk1cjNd1isHtYdHJyCPw8lCudRcoiQfTOTgO7+jd5PCm
SbIQGrqE5JBJdH9VMiYOGQ/6HqoLUT2bA8AMnKqJBTCmgstjEkHhyL/SOniEJLBo51f0ReIql3CF
RpLXxqmEbl56hELgTgTY30VbJHbWm4tTO5D181s/rXgDUqtH9A/Xp4dpGRs52RzuA06hFHzOK1b4
tM+AXdTZveZ6S6HlTL7H4b8sodDoH4D1F2M+34N3Zzutd25thtLCjZFZRtKQjUbQEy2zMaFtBL3t
8SIpcJJluP42ym8nBrDfm4UYHHan21j8tur/UzKSOEuZGcyCPn0Z7KH/fPtRUYivc/DsVxrmO06r
ruipXIV6c50nlx3oMNzD2pdTKgzlG1yf2lOWH6JPFlLfimuez3mTuJUv7+58J8m8HbatgT40uPJx
GkDVnbZHkFa0w+B+XatNdBOO9HrQ29x5sp+EfIqbzUhbnpoJHXQ6d/UZ6FVJ9FJUSx2zGWxK3SPT
9RjfzA6JO6Fz9J3LduRVf+gT3ATHwPSHYwrOdSXTKnboUS6We9b86tiwgQDGyrEIRFN1xGKjQNTV
1IxOyAG9oWSeYDg+XydKPI3Mn4F1qSvbWOsfAghRNpIbbtnliTzd1wWwAZ1fPPdYevpIjf6+Cai8
DuRcPx9Ux5WstaXIznQXDD3M0iDniMKWwFRln8kVrk8vnKKqch4rZMr0smizl0g0q3dyi4FhNvgB
5P7bx+B8ksgQOap9ZRQhW/GvPWnmF9Vi0TSYSsGZFD6EMRe4byExLzxLrFlfdUQPNVUixXK9Ukh5
kdTwZBEitwjkPtWftUyHeyqEkcRipjc+s0Pxx4bnsgc5pjzfskHjPgsrqndvhd48Xw+1ogu6Z6OR
JucccaQ/tLaE8XB7JloXy6tx0fr5Vzs3uygI1g9UmfyRTG2dG7IubyreSwnHozNiz30uw31+eaEz
5nFWkA5YhX1QtA6mtpVPUEsMMfsPBS8vY5JY4NieionPXOnIfZrM3pGl5hjqHvuyGvKol3qgBzYu
cpPASpKzaiXgljQZWmY6lluYLzOQHOPFGHOEqYT/gdFvCrwFasXlab7R0DcI8IFMtjng6c6y55mC
bXA3E9Fycv+ArHkRd5XpDpuwXcjpBZfigT0TNPIdTVrzeEA7OpXF+GvOnuI0lAdPZj0qXi2mCp1D
/BN8SYGpSaBMwNjs4Gv8YfYzlyJxUci1M8HzHlnJqL3nWvBMbkn4sD7US2IAWBmympQxOrER1rQR
rFgDOF+oB1L3uryg/n9Eam7XDiD+KaUVZTiErSMQ91tB7zrUFO03cAFpzkAo1kSiqlI4egN4CuwW
ulZqUe0v5VwTrBUvsbrEgZX2GYtvn/5quctX2SXLkrihhNk+LA9rI8GKXeEv7t+xRg6QgFsLE1oe
v6AlKFYC43Squ0Rl53nyJ+F9rxtIBcbe+BAu28dUOnbE2DxWU4TC/lW+OL8AKrVJ8ogC3Jhrbofp
EpwBRooyQJQJ4AGaVEvfdoGOkfazD67azOWTw9o951d8GZFPosDHVQW4G0fwG7x4+dRu0bXWiddt
iW9jR3NMHI5GmmzFLFDR/keU7yacOID6c4u1S/UJy7chBjuEbvUT9Y3DaAArCvRG8n+buGVwJ8W6
6w1BzQgVQZVTrPn32Xa1GGOdWO/yjw+Y+c6n0l/iDNTSoTG3LCwT5oYXUR6qtnQhqcQw2vbgJgjc
yGZC5OVNn1lq11sptVd+Pst2ZBFq1Llz/cfaYtV9/l93rbvU1yqqZvBzqnUG8Q7COykd8qqvwK15
atFf1HtllJ5w9mDd61ly++dnaX0xG7PgumfsO2EYzY9el0r3EwafJmtgbMXmxtVads7YNnTpj1no
V2nRQxUf8WwS33+ya1xZxS4p8St/yH/GIbbm91ugiigeYHBCr2vUhicHwNUaKfmcc1a2B/N8dvD1
+GY9eTnnxewot4ivKM9nRlkKcn9xqdJBvpFwfgqvTd2/4N+DVdeAEKvbLbiaNbg04YCWKcYtJUc/
/ANbWskO/VxtTJVMqf/pgGIQ2lpwNy6qiUzyHmm1nil/1gBpADQPYoJTqCK+FztiX9SsFqGj6xs0
ij6cirWfPLTKkdrFLKkEUAqWHCUE5Suy5V/Lsu0Z/EZ0ep4+LsKJYaBrCLBwz0WECpuwW8kRYoxx
DNNimsGFviPXpxMedX9Qd5ViTUoIjrGz0/4WywZ28eob1IeGp28u0ejwg9p5ZNE6YMK+eH+5APgp
eT1yLUxFzcYMMl6aeZ7ffdi8gb12KYjecXnbYSRIQIoJ/X4dixkdiMUvJyJCsDsXYu2/y9zhVfCE
vG7KG/+GcZomh+MGrJiJKZNRXd17B94lHIwmTjBCst+dx8PLfK1Yh4eqEp51EwA9JwPWof7KO3Vu
BvW/6I1gbPA7ylq2SbBoj1B0NHuO1SOtSdaKbCFyuDYWvACLIl/y4IdLxW24f0neVeHRWmpxlX9t
JQQB8m+AkeKbF7jhvVhKprSfjscD8n0FLK5UyT+JzzZ/zSxehfVtMSl1V31AjKcT52KViMxLYYrM
u9SqZPFAj7vxN+YXSzqv/nKezl9AM1qC58J+5ctIc7j0Cn06UOLRGyJLcoUNGJORd27GX2ryTrwv
ao2OPe+aqPChMSczC7u7vLVAMOaGiCAzc3fiofMT+wuBU3nfC5/o8KTrhSJvn/wbGxXBaKV6mJ4f
IFUGpxNKUUAwn4Y6APnHHk8eK11JnnfW+JTZcxy3jCQn+XGgTCjojW8WAvQj/6c2wGhavX7/fxbL
pOEFQIGFTsYY+2VrPXO1Zs+lPt119VTamg4+bhRKS6L0jKdm7r3lxCrsht7luM0iev+Dr6DJJr7G
iEdhC3EN0NxpPm2qa2Qp+GHSS5VnK/Jx6yJuN+Ez2AQmf+LhxoevvCoSVFoL2Bw8Q+QnkN9/eHnS
/PWy6durWNBuNcpcw2qCHJFB/uzz+vQJJsmK+aZYckcb2qqkmjMBEIfmjppw07ZTHnO7/v2LdYn+
Cc25wSDwSTtOmdtsZH+rBPeGIkmoG6kxauDw2y4PIs3NRg6NiXeU/Gc9BDzFZ+rUZwnnKIh3GFJr
YNuU/JC4ZO8z2/L2VphIm/kMJQSSzg3XKLifpNcOXKSfUfiYkNyrpA1UFNlRwlm46bBqFtGtASFZ
jR4Y/3WHVIC0aAvATRhuCbbZg0EVjqyk6fbe62+3VGgx7HWq0AZiW7J54xRrXIHSiwvqQc+I4lYI
ZcelZGH/2Iddh7s1fMJITlOzIiECGlLLca4dnR7OCqnX/fmM35nDyKwzuAGc5xBlQSTZybshKSG4
qpv7BkUnJREpCfIhYsD8SQ2m1dJzMn0zdbVnQbTdPSZn2yzB1d3rLs1bpcIDmvIH7K2uAOyc3yCG
DyBNHLqnddbfdi+coCaOjcGKEQy3CgubWFUMp47O0qp4asBlhk1YaNRhdPf6XMdhakKPUNxFNF/k
86Upfj93noDcppMpn3v6Wv12Ad7rtl1N6DxVLDbmY/T0SgZY2kj+SrINM3z/TLKOWK6cUF94laAg
HBPQCYhXMRIAZoZAPeRx4TOWM1Qv6S8mC44D8Tenq+Y7k43KaijkrHetwQsiQwnHwuIVT4YpszS7
oM7p9KTVbiRfInFQyLwbFlFeFBO1nGd7sXOuAot2DZeoP2Sd1sypllPdzDpccFR+vjUpmcPlBT/m
8vktqRA2yDBOefHps+6MUmOjdLwZuXZiSfOxU/mLGFyF8Bw5F85AGsZ9gijmDeZ00OiN5kBk7SLt
CeUySrpwXqVGONw0kO7NvmZwLWf1IPrHJxqkACj9j6ti3metAJYVYt0P5CLimr0yDVakxeW3/0a3
ENwvDUwXWf0hTYfBfcZvj6t6pcNFMcRre8+hFazSFSPYvRCIbvngL7+y+WTF8NNXK5Is7NftutEW
2dyaHY9bnOSCt744fXTipevWTNoNNmyb0OQuquuCEJrnzVjQA5e+lyn6AX2IY7Ij3AKquc2LktcC
4kAerCpgDG3pJSVC1bdFsAkkhvC85+iNr91pFYuFkwPffzkzZM5VNDuPiA4mRNII9hvVArJ2XMEL
R2tzapPhlFzQZX+ZeFIPDeUrvg8pKcwrPCwWDBbClGg2dOyVeOaeepzvDHQ5Sni9C/1FyaB5TjvN
5PiowQdlFfHQV+gKhfiEci7NdNhX19/TL9FFyfMdgSClWzT4oTUsJ+FJBLRuvny9Fn0tedbkDWxI
1qyRAEuB0+ikHLAYRsSkeMmYMmV1RfSjnYjwkoXyBrChE+v4jmJx2lTDMT97o35KWmy51Z5cP1fw
411b0+fODpM6CumqLk3GEfPYpZVnu7ApnOgcb0jjKZDj9SE9dMsSsiH0zsyjDo3z9L92r0AfGVlY
HrDLKz6mqdh5HExoiCnSKwPUf0Dzx1YSVpXrfzPymkWsL49TAsyfyvJyyGC/wZ6f82Us0pV5HvOW
6wgzFrkPPKb52Pw1l0WG4tXkGjOIgdxwkiahjdY8JLHaRUpmUMo0DYO9PrFAZ7tpSq0RJmm4kML/
2pKuzgKk2rz8YUfgdV4KJcCfMM4zgWF/pi0BGPYYVtYTaSxRUqmhN2WTA3xMqSxhvNkjoRdY6GtV
kvQN+rzL8w2sqy3FsdXuqBRh3gYxYTLKpD2XyFjJwCWmmyLRw80oFFQF5mkZyevYCPncpWJPRY8Q
1W+OWyMgK39F6OFk64Apss/Ubk26AYm04Ow2w3IHe6I3JWk453mb1bdsOrU5aHZ4B9nBL/EuxjTb
HlLjkaCRSv8FwjRrIqRViFpbSU8GdAv40rn/b9SC0ao9nAYsZ/6ypGv0VoukILpY5t+V8kKfP7+p
6usHd2eJZzvBjua8WL//9J5keraSAYH9J008oqeTo8L31MflnLhSSfRnLHl4dwqNg4dFyDk0f09U
YJJykXHFK72q158sMLmR+G+ZO0cAUkv/4UwN/z3dGJ9Quh//zgdZ6aQTq++DH4TzeIp/g8oabPQg
Ge+mSOTGW7azuTpYo5dmp0PiPw1p4u6FeJZ29F0/KEWKHP0yZfko7zpApaYLgChlDtXnSx1gNGtn
6Jgmsp9dLHs6qRTGu3U6pZu2wkILjbqiTl7X98FjsOX2/Dr3EUb7VjezMkd68pGtj+VSm46q9U0v
iBv1w2zrf7mJtqLj1UrvrcHy6FgySUUcOOqZ/Ks1Ww+Kr7/TNsbHHJXXNtn4gQ6yhWKjOxeJfPF3
muSC1nIgFq8J4gSaVIZTIWn5wjrCzQKl2qOqoj1vDjvwD4tzUS6PDLhv+VTMk5mwRvzVCpqjyn69
ALMB6+s7i11ATZgQ3/JucFRJX5gex4hwKw+ytI+kHxOM+aDWaBhzxLld2AQUIhhL7fUXXGL6xbII
guBtygX0dhoF24FKFh5id0Pofs/4so+myMJog9KAMK+U4G+FKUziGJnNNBvSvmY575V+BosZ6t5E
S20KL+gu0riPeScj9CAPe41Bn3htU0mGhwKjRsSBcSL2fwdVJeXK8jv48EyzXtD5KatPEx21W0y1
/QqhzvnCR5anYj7TYdB/w9/MagWq21RDofwQrqjD9gxjeTOJ9diw2vYH6jyEz3m0oAfVRHsrq/KQ
gv+BpvqiGy+madmiKlgUYZiryAU7RIhF3GfbxnGLwY92jaSNsa/nGFobXmf+viWxXPJO+kQ1m0mZ
NA5G15pfN9rqTXMpXvoSZsGwMn8sHe8rXXylNz67CySRynvJj3jyA4o2+dOK/amJVamQgvHMNkvU
hQlE1PB4CZH0ML4FKuyox+EWUY2n7MNJXtSuLgmTHdfwNHTebjHCzMqi6AnjnxiURog2XLlR/bdJ
t9TF4C8hhstZ9NnNuEWdbwJ8IWtwrXc4WsVR9MWDUBarcSyDIp5zZZKmXS6Ieq/8MpwpOG2nJfTj
3+feXVVN+8ELUvqkfaXWnZfXEx8o4HjG1hd5tU54soFPavq3q0VgbyAt98wMwcnnIhTwBduksrK1
ZJ3XVXNq+EKBqOZv1myPu+aySzoD7C0pkkcje10f+piKoTRJ1FOHN/13lHBBZxURQvrZH4Wx7Hc1
SAe4fJwnBSkStqpcZ9NGDNXgZLYunKXqnEe0kiDmObjC7sKrp2HKYQwWIoUzBxqMRNcHkKl8DKu0
Zw4cv2AdAw2Nvcztoec4Xo71j92ayfhPuooL5U3lzjISkMxV4DCyNOKeSiGJjKMjWKS4w55gQVBQ
Vke9fPh5DNw2w2TdDf7jyEvEhWU7BIStA9FtKQSWvJZ+wRfbExEZlUIfmPx0FJgOQYHuXD1zBvV2
yFWiyvhfxILXWeFqaycBxXns5Rbs2faDWERH7hynfSBpuk0nFXXOFdq9vMbTrziG8KxO3eAa+U+T
Bl+sRUHLRjTqhffn8PpjarRcEhD75fqob4ipY+/LLNpbQyC6ItCIqkeH91FtkS60o0gnbSv0OOjt
KQmEuWLai9hTc9JpiaVeN8LRNbwNtmrJOM9b5EgrOiXETD3UEtK7nLmOg781o/GG4M+u9VP/IG0R
mmqivSN8ESKk/SCJSgEcHWHh+EaOEky+2JiwdmZfu4nuGykB95qd1oY0aU7B+siojkKyfLsQjcjA
jtqlbjVgCHHDl0CxekvRUv+aGiN4d/S4L01DEa+S6vUJm0CMfiX+ZN8jwEUXyGlaNCY/Q8zBW0Dw
nWFUGOVuetjVDxYqcvNYsNso+roKLn7BBzTXa62OZGTiJ+kBS5UuyOzmJtjuVLm0WNp1Wmq5s7Lu
R07wMr9OtKk0K67STH08f2zBNVch2CAMulkULvtDtjSChl+y9Kh8e+KwKbfpiSsHRyQz1f66GemV
s9XBjbTlor6ZvSFC10RLGIY9tMUBi/UrEeEkJcc0Sd0P/2qoBWmgW8O9MDZ7pbBzyifUEWyjRohJ
XKoIi/QocnXRjEWooI5jv78Ll/aASZ3fI5J7ynOY37hb908amHcykGJNqTxjDWf+7KWJqAYSybrV
0EUbLxpddzDIutQiGvMy3U1nMizFQFQLP7CIJyed75ODV1Ycd3+fyLUm5fByZXSzMN9ngeah+G6Y
xizJsFlHmdVslMEddvnmJOW6+2kUbNTqufUmTVs9XjWEso4YscUO4Drm8SUs+YLiPS85tXvlMm/G
vCvEOOYkRoz4LhHxsPOa7pUq07r22G36NTKiKZqiGgfxsYA8m6x9Y1di7XJMKWRQKl7x37q3CYJm
YHc+haABNlX/A6Tu3rQAJjCi03nDVpO2Pn601tqsUxKEY8VK+6TswLjMsmbgXPDcIKqVT9g74KRa
SEMIT27xgfQbY+YHtmnyFQMjLjJ7JMFbxulbfUhpYEzHFfj6p5Esp8jw6LFxBKTJUkZPtMLSj61C
7C2icxRMdeDL+Ni4XaezLFhOg5EzVJf9+tVkBYCFAIx/1fuwt+Ofqpi4VnYt0sX6ZpKd/QTcOQQS
jdEGAy/LN5RQFJ2LoOualEFOzpj8JnJbD5N7snEgFayWTOCfqOCxV6/p4RoyetScHZuoJuln3f7W
DRlq6RoB7LDoAYNxr7U4jkiHAqoIwedrzUZzoKOCEFkTtAIEb7jslKGKPAB8kpTbDBzKQmoAgX57
xbzzrwuiiSjAp7usFq4KppcdtO3FrBVRRTgQfCpSow3yvtoDemznaziMAhbyvoPeQP+vOWyp/WUS
Bq66yfnjyPyfmmxOCDhNljJmlcFpoNoBQjmeMDTXzFZDgdUcbPc/LMwGNSDCwCF8ngVHmutaJ4Ru
4vlBh97kcXzIu20rkKcBtAf2XfTniNUKramrTlcWz6Vq0BziLHFmCEDdYp0H3Cjhp802rzxxv8x8
OzIJcZcAYhZdi+vqmIhW2qAHEqe5BNZe6aqZIym4BHNYkDecq8pyd1KSDCxdUI9L9WHz70FRQrVF
WkNtQS58qgN8xjJltkQsbd1mywh6fRSMxfxGvMDnggH+0TOI2Epi7GG4RTsMk7FkScGpr3U+HCSZ
+6iXlnRKOZZ+YPFY9qkjNJ9iR74rGbaJbjaOUqXTvWJYVUNVQ8yf+5GB2xrLl11Juxg4VOC5IKnV
87ZkLz9ga7JMo3v3GgFf6zxpM7g+bpPgSCOVLFNIRylI8rCt3EfvDqaBtJGMbDWyFcO+OxvvdjJf
xFY9L61OQk6KApB/e8KpzYwSRrntHG4/sgaKhSRFdN4kczT+ZIEuCd5aZ3L9XLEFB1kW4x6kvC/V
PekQWZbtlIsZFpSaO1sTM5YfvJZhRE4wFsQCP8MBS7d4YDuapGF8oWO2xwowa1+DudbX/enH83ge
Gk0r8HTsSkX6SMzWNFrm5Qa6Hoe7fb0avKwIa/heAXWYVmEIQY8hcFCraccSfcI1NIJHfLoa0zJi
2WbLtZ3SioIQtx1benP8LKumoXw7CCWTM4LtJJEwIXZeldL/2g1rsyuiXiKRl7+hLweQMCRqv8c+
+ytars2/fu+LadnuQo9EidWfRl3sw1ucRFQnHEIzxKdsxjPW4fSqvnbA6NpPGl8dDzztHwpNeBki
gHxVip0af40pIXFjkJjfBNsm6lkVlg9FQNScD7/kWYLXRvepGxNglBmags/IKlqkQqqhCVRP1S+P
13tvrZ8n/VtFXOU59BTr54JpWBD1R9oNEzGbsJUvOAdbC3FZ12UFfNr2AE4jYGrD8mBBZBdA6W9B
U+o2R659+N58bLhcD1tA8A38IfDoEhLpCO8FAJ//6wtd3bi34a2qlMd5tW12N/1VGJdo3Y05g7xm
k5Zmcc9mwbstOJ9ci3mKUbpD0tY96rKuY56qQr6dzCVLzn/Vir0qvoZuhdhzkI5lbw8ZYKrV+0eA
BLlkRayHusKlxBNlOwBhJbusaFPT6ihAiBkwtniFG+cYG+BgDQA7Tbq7aw/GPAQftQliENH4U1Xq
XIMIws0g9PPuxN1lnNbCZFPb2TOazjzPPLoAJu7tUIkKyFE8ELhS3khOAUBb/6NGJP+64Ngr++oX
sge8KQDYuyq7UO97tbLbfquWFCCSoWFUuWPC2dDGtSdb95E8/aDJeB08Q1B70efLsP766sOaypVl
g43lSkn4HQmdpEC86CCoIAdJToFcq45NyWPB1OB7dcT6hZCEvhHBYl8rG6hp2aniYOlX8zQm8uLg
hCcXyOoki7EqYacCX3W8Frx6XZ+2B/wUxbVE6mffTO5O4AwZNQuiZ3mvJQEA2+flKuJeeSJtZcaH
vs5hq2B46aVcO0iLFPQDUp3lU7Cf4Gs2u/EZg+xQb3dt/gKE7vTFlMfdebJvpU3CJO7fpWldxjN6
b80MFt98cpVwEQlE3gmeB5j6QQJPiAyivYSVWFUB/4HW6UuTPtQ5dLyn1iu+kyrwlMZd6fj6X+HE
yj0MvBMK4W9sdwUWcyXFi4i6qo5ifkTJnnPBs1YtE7V35b/tl7DtVhtx5wIx/SijaBX7pxu2Bub7
WDodXItDTXjUhIY8ZWSHd0B6FmaPRVIVIbIVFqXKAgv6dviqk03m+N0naTpdHo9w0RuuWGc0Ot7u
YGyzqKytbS70ekvKMzfCKygyKleiC71a7vG1YuEJ29pLO3v0z7R+07tVzpS5eil73kUIJ/xuPL2C
PQgf0zh4Glfk///VkyFY20HbvnRK9zjc4uItIFQfVp8VwfcJbWl2xTAlPAOcWGCMk2j8eutI3mdd
cTbqRxAJKIKBECf6S6siy5LPnXBuxBJ6xLMsWtlo6MngcMlI5CBc0Sk05zykjQt82VRF4qJs0fr9
RTSjhB4KTg11scW4OqodZCz0x0Hb2SsF3/ShfKW58qbdA2i/kqMxZWrY+ZmewMODcrpglfOC1MFd
MROOFd9TYBEZKJdVR1a+rb5y+PKDw+9tA8YujWuNvCupXvNwJrOBW9yfzgtQoROqXztnru1K3YsL
r5SkiIcx97Jxhb8oEgdHxdZwxXrkeTbgjXxTVgJX/sct3Kibhg/J5fBF9AhxP6hZRXx/cGI6mGUp
/XeTso5tGJoMQN5xR8O7QXsvxQbVIEpg+xe1J1c06Rt8ggrCOdz6nWHrjW5bMjxeSrOWADW/DOoM
BdYEzFK37KzyIhBYs/EwPdpywpL48jzp9Ai5OzBpXipCvm41F2sa2zkog6EkY/4J5sYjlzQ8GOiF
tGBNJsUiuHKrtT/pEVmm0C0jwZYTD2SwSJiGCiGBhFS3csd9e3RG1hkPioKcadPk+WRhdAm89Odd
6x02roIUh5cGn0YZne7ORszV2gFcr6n7vXXd7nIMi1vb2AW4Lu7mSGJq8vCwJCi+wF7Ij0du0lmZ
Bbnqd19v+1e+EXNv4B5PSxNSaDY0vtwKGy0ib+2R5i+xk8SwZhXY2qQMKjwRAiVR+g/tI2gooFVX
Kru+y6ShH60MirKz8DtF7zNECRli3ETi+vWPousyw8WMM4La69zUsomDbBMXfqwFEIe6JIa1hMPy
UuaH8ZVR6bmiqeSRTu29LpxKqflOyXj5bLIqTmtiyukUB2JF02RnMzxnYJj101Cn1eKld0mo3S2Y
d+lJlKXUz6bKB9Xf2q60/EcvgV9IDgeWzoI31fYflXVSaQJWLm1/sInpYGzEAvlibAyzVd7kduue
VnfpcviOe0JSbGC9rMZidFb4xNOu09A3A6V5l0xPM93hNBByYb+guSoL/0zR/plqMYfP+qYBmBW/
FZJoJZqDUPWLb5+Poh1yRg5USjKPu9hFyTTFuZjwn7+GfCT7tBKTqJe6W1wxDdVsS8d8yUfsKCzb
omqhFctfC+YXcecfcrjygSj+Alwo+DHQOdMTrG8OjNkTBVuovaFKkpzjxfkOKtTVdZq4GhQiuj1D
UQW7HiFpJ0heB8gcmRcdseISzM7HSEziHbUKtLr5+39roN/1gc6UedUWCMxcFvlZsoAtGyAIdbOk
RtDQ/CfPgrMZBoL45krFWEvB31zwSy0olIIrf5+/ZihZm1NkSc4k4+R3XiyhJODcbgaruiY24a1K
maxRdBg5N6wBu7p12fLlnlYK3mJFVcEt8BdpBdrpcYrt3OkIY8jx2jL4zKt/vS3zAd20YYs15N+Q
NVdNvxbj1b8AknSnm8txL8T+Cv65Dc9aunXrFFiDtxYat6x0Xy6PIiLUr0R0skU80CbjUpxRIxvs
YyBaMzYpkr0rRwOxS55NYIQ5EUVe3Z3I6PAisn42tGaL8skUg1n+oPvu1YYkCNVLb85qy4F3pvve
Fk5xL6C1Ariuw98/5RBc3X2ObYx4z/dBoPKMxikCBmVF/AyR0rfNf9osdSXaybyckHH/rFcDPG7N
zGV/iRHUi9lm45dxg7cqc+qc9kBVNR9KPm6nLZ/wBQoe2xV5GyVwXCILz+RCXN80t2Z6CpPDMgEr
DvYJj7mKg/D1TrAgIhqQoR7+oKHBsBzah7e3WKIgrLitszVA2PlyWTxqBMtUjMFPqRQuxbRFcBOl
Uq/a+Xe06qKg5Z9K5odB8a63cY3Lom9SuxKjUQGjUKSZZUFUyLN7aAo/QO1uWTGEXcOKRX3hQGc0
xqwh2i/GhqBk9ELnAKSiL7VV52ZB4lL07pEiPKsGt45RUWsWADOph4CLXqax7Fde3PtWv5K70Yov
94Shnr57KaLU9MCnh9TrIMMT2tsCMr4tNwPxiz3mGsJbUV0oHjl9yLoNjudi28q5QcPHf0CceIBy
GJ0gUzwYt2EM+RPlwytWMoavA/gGcSOCUmWrq8zGx787ehLyoinOlsVDCDQJKPJXpWzl8bK3ylOb
GKjEquEdGxgfoHjPAUnD0t1dqPqoGbCZE4uZ++A0e1clBm1eBFuCATMO6lKrylbedpkJbgZYZRrK
UOROMHl66huS3CrTJWh29Pa6A1coomrkyKPVkSTDPAYW2sOLI1QMGDIvVl53AQnxLbiODwX7S9Eu
X9/iUPpf5VRoMmDVGjB/0uIe/wflsqsk1+LSwYD5yso0zPu5r+9VFYMRekReZNk83PmMWQq9g+Wt
CAw9xqABMkPNoTMwewaJ/HeqwMsdpAn0PR5HsDZLCP/+IRzZwMOYCexCP/5blfi/ISP/D25XNPMr
f+UXKc8dQJ5Q1QpeZwx83/wkiZu2YV6vEehFoSkAPw1x+wTiMGW4bF5ryt/KrAjmnaWO01pjB53D
LlUcMj9ljB8Rjq/EfMjldwpWMMQmVpMcTJlQLchsMuVGzYZXzTSnjrTP1HAK34fmGsakk0G1v6nG
nhuBhKQcdWCRFteJPnDGjsm2KNRillN/fOL27g41om0a4uizzyWEoL40Bs5yZluzmkVcq+lMtlE7
56E6yWJdY8Y3GWy9uWHxIvJxzveDaEYJv9TMFTn7yX5rT/OcRBNlzZ9sbIuBmE5esPOM/fNGQlPh
bV1/Wb1PKIhQR1/1YN8SIBt/aX0fyvPrfJQZd5Hvpnu8e7yJGhvk1GCA82KLRiigPZGob2RdOHG5
31nNYLjpDCQ6s0rIt3sg9v2/50O9+CiYq4FDACHoi5nOPm4NsC0DUKg32ZQgSMnchoapqVDXDgzY
jz7y4q4967HLOaqqOMsWrEVQrY9WjedVsu0w22Lygui9en+JNUmYYZ5FMbKl3LMbe9JEjdg6cEv0
z1FXdx27odMy7nhivRapw8htqLXac9w2M0BXy58mlgRhcO070lwJlpqiR0/i1Dz13lYIHoIkPQRR
woHZVXA9VC4dNLLZLdMa0mRGzZIlpuZdJjmvtZB6rWdmk18jV1rGSAm5ivvnLCxj/Jl93TRUhG11
0i3Y9+SULvMOU49tu9lslPe3YSPzhIHQCg59lygh4JUX69JuKAaO8X7jwYMsls55DDQKIw1gTg2O
O6NZYn0XhWV/kTSoweX1OQho50L158U+A08xXTZQwa17MHoYL+h+l83WKQ0MI7cC2XI7/9iNQZnv
nzq2IpK0DvEgt70shLVGkgw9avvVekTO2ZUvtuih/1SJoPLTCxHIaBLQXg4t0CVCmGSXkn5efDET
sMufNqcH1Vqk50vFNYamhmSTSN6JQjwJvX90p5OHMxzJbWNNgYLpSxyKfhucjeeCf0YKpoqmmiav
mHiTgno8LUk8gMM1nK9JKBiiGqUkxh4u873Yp92OuOy3fs4TuApqaOLMtDEC5Tn1SFElmkN1hUcf
wOA+HjjiwP4PjHFHGf2mkkM0NtpKRF24Q/Q7lObSdXQR91vui5sBhGr+MOKzufxwBmAlPiFIsIvf
uwuaUunouIIYlpPeeiRUqEVhgmCAeC68ibbUU0ObfOsCQZd7s5DSOF3tDO5P8NH0705TdekmBxcy
TA8agzF+eagAGClx60mEaJ6VA1lZJlmWjsa5ZvLBAt0Ygyi+8tbnOVIn071cwy2B7arP1pJOrkTO
/vOR85UGzt/faarfpWtkp2yyVyE6mHa68AZBJ1TB/Svs338Vhfhr+ZPixz7XFuNjoHTAQf1feIUT
+f5KauktCcizch+g0kTbCbNIDf9uj+QmsFaICilUiKZE3Ecfz3HMFUz5sIdCAqGN6T05J+MOdC9T
0o6FLtIdDuM0QNWKXxDNL+g8Z4MhImAnKOL+3UlEBdtxMfZW//Kfvi/+ps/pur4A1i7powdhNiUr
t23wGggBkyGgjKh6Icp9N7IdAtLhWicn9L6hpcFwuQt5C/r2W6S+s6lKG6Cedr01gTeCejsP+OPn
hlqwSohsf+06yBHmEV94JVL9b8h/k/hK/gqYNecraSoFcs1QzThTB5RV3sUnwEYEYH4T1wMryhvp
T1roweehtqrib/kBRKs8eucuPrwwY7AjamMJyVWEXEeWaJsgz3SGxZHGE7kpqH89SS8j0Av42wpe
qE7ntJJs/I3Q5MZt+4KAC1u/IsTnrU1Cw0nzY2a7PL8M8MaqcwfDAFw9Tl3HgWPf1yPW5i4Tc4Gi
ZYK77RcvtikHkCCMPF31ve/GrvR0WdrlbA5RBarnkrsqFxxcHwUTY8XJ3v+RFFsa1qyGxMPaLrDw
j2U644YiGSKrenhQSEziBrsbQs4vHCyI86SPQ0MehQPQHZSJDpZLEhuO9qBNCn7ZqKJxWC4RkyfI
+zrPMauxuL5sHOnvLZSOUHkcYcW+bL8bXzisNoy2/coqJ1vU4l1obB7IV3rP9R6045VXwTPJqp7l
9YUTp5vKrC+3P6m/Zyy92YFKW06kdmnDL/xSUctxdMmnE2S+xJdPnBhpD+sFxO5ATynlu2OkkUx6
8ofTfbq9YsFTS8bQ0OxLPn3YHen/k28a1PxxZirUG3EXLHotio0GyOFsuiLBcGAP1PBpkx8nZz4S
iNqb6lvjzDnDwjvEJ0hPCZSS/4rcDa/Qda4ntpjXA4MnveAPoXNk8hydSA7B9MLPxpNwGEdm4vbR
3lkjRQnpgtMMWPTdhw+wp40NdIJ5hew/bouZ6uW8PJdKKTu2IjVftc0/72ZH2XeuZU4oRqyRVGxj
8em7xfuP0pgUU/1NiHmSgIvUkh+yZgsmc8X8tYdnGyU30LfQsD/2/dRrrl2i7xh/CvAZd6mrtka1
9LWaBRXzMMuNP+VdRsz8Pe0ETRZW7kW/Z2XbOnuJLAwgUuk2cf7OxYKQJv7wsAmg4fU3yak3c6vN
F394DhJneyVqjl5ZRO15erBmYNWdzGfNLqTI2IIZGh+wZGeQKEUHOkvxh9DJgXrk8ZMYIU4RV7Cp
ZnOIqY2Jce+DjCXvr3t35fEICceC5SQeTTXR/7FF51A89Y0rpKhAwuu7hjyGl+bV+mJgU+/VNnj4
A1VZ1n4xQ3+n4vc98/ptRCqnCI3v/BzdmbFREfbw+DcA6nA+JIoFZc3cwyw9qiaw3JtXWIrt0wDO
jfcZcLnU/AM4U9w0VCVlZ74T91cs44mOj20n6y4PTOh662+Sm9XEKmQxS2VMNFEji7zZIQHzZ8j6
JaXPsLd94h/tlpsnFEUNv3EKlebLpv3f4j0tVu6pL5IvqHB8EtrbpLg6p4QsPAFDP0FL+VMn5ulR
jHUZB0y9bUGCdJ2MAA3MEQN6Qh20JjeNUiT040vuKMGztKC9xIQ67U3Zf8UJw82JcnykrEz6g8lf
cBjUSfQdns9lc5qb/LOV3bdjX5eMkEZBxCwim0d05oN/QQZMNkBUvIG+kGJfIaiU6mVqyfa0CdxB
6J411dylHf9HAN32hyfQbV1Rn9A+NsftYM9VMVw7zPoE6Y9uanlrju9TTSFKMfwxhxKQb1gPz+J6
k8ZQOi0Uq2+Dh6q4TuBUFNgSr5poh0rLPUt0VRyX39nkQampTHQMIKAfpSiXTnkSo0bVhQiUrBst
57LvEoHDvFsRCVBrzJ9Y5bQYpBit1MiXpmpjdYzGe0xleN6N31VtoBPqWFJLZHPY6tB1SKRyGAmJ
jkVJUbmNNr5tAd2wUWi1NzKuhTliTFc/dAElVmZQ5n0GyD3AMq9Lk2fXIWMJPDQKiIQYnBAjKdg2
2wyUikgHeKcvGc4UVdNO7jHdXkyIdD9mMY+3Tq6bixHVzojiO8tAW8e/FJHKwazf/g0AT+iJrbFh
9w+JRVZeTt4h/PJrTgNmkiboIkg5l/OBGEeb7wgAIUVCrIr8/vWCaPgm4VAXznMISOz5iAsO0d51
/ZIuQBO5ZQveCV7wYUwEQ/ck7+hEJJaV+1JCIrH/iT7UepdK7Do40P//abLVJMVx0YwXWLZ9DYwi
LLEJpXgXntAdzI90JX7TsjouVInf2+95CFZ7LpUhhwsIWIXXUXVwk5JGaSzJXoxC80D2fL6M8Zb/
3YKanPQ6o0tnKMJs8hSHOfmkvCL6eBHWqMldDT1Nyf83GZr14QZIoctYCyN6JXqI+o7CjwEZY2wN
G2lBVhNrH9Sklqi74jS6QG2Jw4Yl8GznUogzIcn4dPqH0HSKPbAGlOrJDWNE43G/tOMIJidKSKMf
TdsUzujNEiMBFQWjLgpThNibZ5kMSAURbrdILy36AQ5ctyEKW8/ZeEt/H0BBiTBTbB5pXBgLdQ+5
U9uaB2Z/kL4smQCdmtM5vwSXT5+xiKPI3Scp8XRniGEZeXu7fzs7aXnVB5lPao1gP+CKjJ6Ue1Mh
ApEi55qeYgh9Xp1iSddIw/1/Ba/bvbdwchE9kq49Q0NWtrfNF/w9TVCBUAqNPmdECC3X1pe5Dsex
OjnCdH5GaVapJbamynGz53yfk2g3b6lABODkL2CuEUtkRfbvGP/1Trz1eiY1Xf6KFvF/Le7Z120T
5Bp+gLfvQBtJWyHuKV9LQsL+93pYZImg5UMLbmRcGAI/YFPw2073TGuyRog9ey4Hr9r+pZ2jRSfF
MNWCyJAis4tQlr3Uu97nXaVLwha4BnIg9/43fO/DQ6dtwddRJKZYKSog7gvBfm3m/Z7OeEnevjwH
7sdrWKs5o9JGfZJzElWcbjE+eZh7bhsLQCDt4M7X8kgizAnYWoR4UR7shPFOFUBaFRm/AHAuvaoL
rALXXtjX4S3nI07QHiE2Zt5P2vI2fiBhb6ghnFjqGb90WnANgx1ZpRCW/yOCUzqihyu3H5pOwA+h
pxI3elaEeLgfW/qdqL7rOoVaDfICrjSaPxfRI1ESDMvkEuoIEQLxO+zYgaF2X1mTdhK4kSN3yT/j
c98wzUVVEowwhlV7sxgJrwcH3x6CJe/mpUht4U/f7SJcOwIcm4D3tuR9odQzYhjNusYzyzS9mmaZ
p37IqONXfqkmrQs6IxxGEnCCAzv8QuCKtEftsbFzabZb8mQOXcTRM8Q3cqdnGswDfK8D29xXEHnK
zSSC9Ggu5zk0M+jLY3bC3ChQNqfGjJJQfbO9bi/R0WHWpn/weCpYzzKY5gzT1BkIohgCNe8LTV/j
uwDxDlqGAmVvdyOhf+qQOiorfncgtj7PJSJ+AJ/OUoTzrXpphtGSHIy3EZ4ZUZoKMK1oVGxHlAuF
dAw4gUIGISNRihBnZjw8cs/Z4DqM2iAR8k247EHl03mFYynb3hXgF4YqDaO+IigOVySmdjz0DaOw
Jlzk/g0tBtE6EgnLxA8T3sMCVxlSyhggEAZkd6m2zPrImOiNUH/E6onj57VBhLcLHmZlQEvDyugG
iqNsFfNjZ/f4lQeCyLINVHewZ2qfUD0v/tmaMV/jyhDS3VDheYxpnUuYx41E3VhrtBilKrrCB7U2
iW48b1rkyMRZp51YuWygF+k2s8Pb32DEziwxjSEwniHQkncYMcVFSd2U70nxep35/wbKg4HClejA
cJd3GaEUvpXDe7yzsBN0Vo8BsWTr+2p0ijSiN2/PPzqjf3JPafVJrplPRsjSTNhAKNubi0legrlF
5aLJJXutipPz04VSIs9S3mCxNcM0gctWjEnNIxp2EaT6XSxH6OUSY6ogLqd/Zxj9j1iTfVQk8i04
kQSc4FVm+FmcRTbGxa2m3RrotXN9XC1duqQHVbKozYGYGddFf8cXxK+SRqfHqxhJNCBE7+gat6y+
4n2jOOh+H39T7bzPWccFQ+MY1tFfT8cjqAvevk7yxo+u/Tj15oJvHtGz2SYGF+wtGZR0OkrPUDj1
e+6i/gfw+ZwpEO51d95TyaukOc7/jKnLvbyaPbhJJ2TFaHo6nx3as/Q+qPDzhrpCPegwvk8rcBhA
EpqpjspQukXF5wkAhin0NOZO0n0hXp9OyxbWrOrERLd/DBxTTAFXuaM5j9ZPB6+VZ8zIoF6+mIEM
GT3YWtzmgErAq093Vj3schIA3/16ABEgr23FLSVpNMhV/OXCMv1PrZ6lMyvc5V34hiGOu5QKA/Gb
pkGyvnsusLOIXeB1WOpgFovP2cyRCLdjhe2rZnF87nfVZ/cvsDS1JRky6kQ9WyUC7TbSPoRluFkd
ZOeSzH1QFrZBxSJQSkZ5uaIwEXYOzaM3BLeI49d2prKOhTISqS1wVhBZmFKLz3xKPeE0KB4WRkTB
st9I/lyBcGCQs0HKc6GGGtct0IylIe8irbhaeWFtZI72gGFYuTuSixK4BTw17hY8xCpOHpjVh5Mz
97CR57zKmYv4/CI1XHpKcYScIhPRjp5/ChhdrXoc6N8o85fh6w4Q2mIPEglX2/jlQ4qqTEC6sbnQ
YLYpEu5Ru/OK+E39Ap4boCinaQidVSwCL/g0Kixck2Bq6TiPco4Cd3S1NggknySSPJ8onVKc5by9
LoPY6UwM2nFLf7kFCGJ+0KPKd6l/U81nmk3s+tFbqt1vd3UktLg9H4sSssPboeVGSGMSUzBaaxdv
YYtJGHTFinnbw4Q8hgxqlcMGIwZuLxpjRMonGjn2tuB1z2gN5TF4f3f/1UlQrsiYpM9M698q64y5
o8neZVksubx73rQUuppLT5HQtAF5OSAnkC9B8C6/5YP342DJajgxWmv0Xz+gYCswudIPNeSG2X8m
ZK7X0DvCdLyLOz4rwSyqE6j6FakgnN4P99a+syxX5/NHYES5lTmtQXdzamTn2JMUVpzMMlRuy9vb
y8WwUzEu8TQkYiu7T4fbeUCdtp8NzyD285TFHzKw6xyAUXV5QN3ShgqhxHTZtoUNYZMjI5bjw0AW
QTVfu5z/86I8hSD57a7kaQ/QW3/PQbwux28zbpzwTfM0DY9aFGkdDCSTmApCbbdldNi7fQMKan0T
+uQYOE+g8kTlTAp0McEglIS3cELQqz3qm6zVTZEOdvmy+kJxD4tT7NAIqDy5w2kfSB5iI9tkm6Am
hJl8tVM8U2Ro24vVSnUiLBmAugXz2jpL1IS0jQz68Rn+qdhyTFj4NAH921CahcH3H3+L5GKNKNzD
zRx0eijc0nR8zkP8zXPPJlc1nyOX+VTEwGBnI27Si+Lp4jwtsG1gatL8FyL/cOrOpOMLKzo9V2Tu
/ezu+LOE8CL3nb8zj7bp4WF3/CnDc4TgdtQtrJMo2R/PlH2afE/33IfmN8BgBomSRqbbDV+b/Ko4
vYtAnKJ3+t4gIc/QDiBG6+ZR/BDCdDLnC7wr3Cj+ed22L1SFPUHUw+DNOdGh/zVs92j5keZdgsle
+XjvpiR67c7d040y3T+jsDnOWsj3CJT5/MmdzkHH2zsGn7FW8tWf23qzcCeHGa7rUo40LxNAHx6/
wNUdZjdq5buipdgnrTcbAat8CDWbkkuVQeULW+dNoz+P7wljzkP3rCy4q9CcKO0dmVAWTUESecel
ic7q3MNBCKP62V6CmPcvoeyP0rJ3Ikhtkx5dQso+uynOiHW63w2skD7HIn+HCwx+aAw6KuvEVX5T
yVCb98lJ8mv5LQXgfR7m1H5rLxizf9DYX+9DKhn4xwRQKFAho6kYpmfV292yktLWGIkr89u7ifz7
UQVl5HLmjkgeU6H6heF1BdzS01LjjS3hQswYmt0Ud4X3Xu78dTScWiscrWk6UwBw1WlxVZwQAz83
gebTDOJOh9RUo5N+0l5Vw1CmiA4GYj26uu+zSuS3/b5PRKMuCXqXUL/3Y9+3kyDoKopXDSVVmb6d
wpIgbowzlANWuFBKaAcoTv6YKO9jbpq+Pq/8ISUSrD3oeE9JNduqq/M44tdwT3Rla8Z47JDzZqeZ
91GRqeZvqRokAcHLGHKctyLzWm0pFQgUa2x9e/+YGxPbYcCLXDqM4rloYgNB4KFrejMexFMG5nSG
gX/tR7ilVjl7+/8oNqWJ96ETE4+rkgYpxcRHZgJ5JhwWs3Xg4y2yM5B8zAzWUWZbhDAbiJwdZ5DT
DlqBpjK4V47Ow3S0x0eKO07S62KfXo6KN9WJdVGndSpmuGrEEWSRCGZ8uXseeBOkprWHaW9qZudC
MqMxgWZUBz7FWNswJC5CIzIvSV/w+grzebh/EDOcYaRqSnQ993Dyq8nRd8X2yL3OinffPWRpIxp+
/wEYSZlk+L+Ndn0560IiD/FFqwKcKkFkcnhg7TFo4KYCg2nJsjkZgsUp4A8p07TtTG+ONyds2u7M
GDcDGgz1y73IqFRYxsHmH9Hc64Qup8XLuItsNRt1kMob9KUFKBU9S781K+3xYUshdvpXysfbakzQ
LgUYsz4YJd1aTS2bNvlqn+YMtCK24/tBgACXBcz6g6M2FNJK18PFWkEWz0mySxpjqKYrekKruD4v
vb9LoyK13QNdJEGSRmemqUwXXGJux+OJHZ5YwQV48X+Gqz2lAsUIJxzUFivSSWNJAXg0Nm2wfCDH
65Czz6YexKMkOxtJRdk8tKvqfRuPruk74ScvVx22cRcsud943yCBrQVtI1TPI9RMdrCs9EyEcy30
kFnM4lAaCyvgAe7bVHGObiHC7B1EaOupkQxbd6fS9uXnYoiVvSsGsjg+V5ICne9elCWofH9rVICw
ChmerTB0bh5hZhyFYNOYpJLB0PcTHe29uc7w4oVxX0LmD1N2YK1CP0x6gto5z/pg/NgKzVdBgakC
N5gzCT6W08pwmrZIwBxZTzreZ053i3huTKUVehk2AC/ROiUxK/rCROxVtxmt5+L+xfS7XvRoaj9X
RrWZicDP/xuPxJWqcfrE/hIQygTSs8FXWi3SHZiPCgp10d6Vnwq1UexjvQOAR+Et+ThJ8/Fiu5D6
1ml1OqCRDYCeCOCCwsPGnGNoloAI+5JxVO1EJ+YIL2ydcHFMQXbZ1hEhBa307nFdTQe27PXvJ7r4
XLhxsl/EH3hwMckezJtaAfEwViVmkqRcsJ2KwUFRUhHNJ14x/KRBjf2yPjh8KIb7sy9ftHgz73wi
gW2e0hlSRj2vAP5k99pXgbP+fDfjxYT/tALewvoVhidqZYjly/DQoh6CPqHbdoBavLxphfI61JY0
2m0dyOmwBN6NtZoNo8aL/8WzK3Ld/SqsBNyeyRfVwcOoHfhfdvnBPIkhM02mJyidBLIURW90312R
hcly6ym1tux5Kl73Tc0ZHY2e/M8rWIgMwMpWEqVXFNdPyHJ5Bym88T5YHdk98aLZPb1Jx5furg1y
205W0VEen0o7tmpP7ZN+vbV8yl9pD+zPcw8AMYhMB/WpeO5uNJI3sico7AdPO1oLif0K7b0WBFHn
RtCvKGXj6dW8CGbaxVc19XXC0pZP9cZQgFHEltmBjMenvAkuHWPFcoqjgom6XQzL8jSfvx6YIWNX
P4o0Id+rNDEGpLtYfqoOp6jdcJ2LjcHUAopNl5udmS2z7WN2Zdko2J73DCPFEvqbs2CY3jhKydVx
lSTOCbcvBub/ro+4JnITPvGym/yfpWWdUinKLQgaJPyqf0NGn1EUN0BoFBkUnkcCTYjXotVYGeQh
nt3ZYtkE7WEnvSVpQF1RqpeXoyipHLJPlXYC4S9zmT6lBBiiFSlWZKe13TD4DMUDrmfa8U71HrOA
dOcRIdj2y1qpKcZvoYVo2PLUqWmcDWrfAXfZ5w4Kj9s5u/Fqvm+H9JtpCHYQh4/gCrX7Zel4EosL
S2X3PbWaZsNqrbmplM8XDqGdUcNk9IW0YUTX1nw0F47qaPzZI8iivBb2zMjIBaMbs/6u32MuSnxg
jzTiiuGmiPEcA2PNRZSR6OcwA7Wam6WrEKVTWspWA3/9TrfIxIRL+VKYLGUjySShImIX7gzuxoBM
e5e4ojpgrngIxV5O5rnHU7sKPfDZ+o1VsH81W2vzn12uorSTgVXjSKG/T3H/VYA/BlyIDJ7yEkvu
cLm87a2pmSE6jVIS/83sC138LDc6QEpV0hDMSSwJ8YVtQQ5A7nDS41vPMmS/6inaNcaG/8nLLEkn
W0u1fPV1tqKeswaxqKIMGNpDC+Dfjbd1ym4GbyY4ZX5SXBaxNTSEBr5URMBz1Y38JHNyTBcK8606
7e2933A1g5Zs+rO0sBcNO4Yj42VgdaNPsydZLaQImLE0BwNLAnGl0A0NlbC+yASgK+C6+x6f8Rde
oOibo2EA29Q4ApG2toru0ri25kp97bvxUU8UbSNCPCNNhI6ay8npCuWcw5fPO+C93IjHYx7NpSM9
IgwONW/WCpx/juYHELb3uyWHJ4cVHSxn5C+EXACZnhKXtBZU+uQZf+M147fG3XXkE2qOGdA+lX+K
xEjSHJot4DmM6O2Ems0QETmjguLFvmYYYg1Y2s+FsSO4wKeBZZcxpJ6oJ9ZPeqlKWALYqGfgqyPv
AKBxvmK84HZp65cBYTO1C1jUqn5LLVAdosMnxeWPk5dXMESvZRWn81UrEjfb8LHzVWvN3gzXLgIq
7tpcWMl8cJYWr1XYl/07yBMEvALfeRs3zWw+yV1g0NC/ju8otGkSOmz6NB8F57sKbs54FCu3++RF
9SiJ/91TcbRV9m9g3HDiUYJF4+cNZj/dOn3V0EfzNtliIxROayKLM/T+aaSFDQOtqAdWt+qWvpgb
pfDiroI+iPsPW7lkqEKEnlefCa+73AVbIBki0f/097Uj6A2ZFBWw/W9KPmsxyMSkL5Wn3jVnfFLl
/qycWRzi1rZPoRaGaTEJHpv35khO0ZyQ7l+xvPtn7YmZ3o0KwO3IMNz9l6l25ZFGv+Wovzf3ZV/x
chKvPwS2v1YACvafToRkkFfyF+O1nf/+zNUsqS0fkMo+A7tVs4VORMXTrU7LMLkcXgzRDlbUrLRK
1wRxl+6sZ612N1cibIlL6HNGngNukBwKMN6/8RSlFtH8EjtFLbfm31DDjJ0W9jBxtskK3PONnQTR
/hff+TkTeCjjhXytK4dj1VFsOsNxmRudl+6wwyepY4eR5mcEXzlvtH4h5EHH6mX4hln/MUrL0Gtg
H0QD26+4+vXvtId1KD4nWz+6l4ZAFxbbqQjbR13QfkWGXj+ZmPHMHoRPy/w73sYSreAWVK4PDyjh
dgsDTEAl+BqD+E2p8MZNqQ/j5ou0Tp0HsRhv0jiqVMjGWQg5jf13o+5v2WtvOu/gKiPYX6baTfi2
u5NSaOUmbsWzdsEd2IUw+5UL2lWNagUhYB00z7MuhVaYL0IZrJADWpKfxlg0QQOVEWMhGZ/hClyv
riD4i/0KGaaucst3epLNV0HWOrWPhPj+J0l4FYlj2Gdh+foaW8Vga8PwTTdbhy2wsCG6duGCcK9L
09xug1uyTy+B6qXd6sVGJZo9QoDFwLBytS84OohLZ0LOrQNDI1MsqWQNyy0UF/UQ9jmXaptu7ZVl
yetwYTUOOv/J4Kf2LrInkp0x+zzVRHoXx6MI3zBgE1kurWydv3diCYbZs7eonWesFKPglNnVVYvW
Mm6efJ5Ixx7ZxSWqBjuq8fsoNrSh6FBNBdVMMr3OaLjTwGAE1IgZaf1ZZ7M59sBkmvWTucP1y1zL
TLsOLQOgxPwnvrTKjz/bx+QU2cRTPxcJ53Ts4ezOvKuVbDcTH0QmY2pYrGgytHfm1/tLxG0s5CvA
pzVqlxfbR84OUs3QsnpdOjy4EPZYYeSa/hiw1j+IdygN5U2CfeI2GH3TiJB/pYRb04ysFGOzvalu
rXw1VTFNl+5T2YJi+jYByKuqaE6DtrFfw4PBVW22RB5Ll1YAtKKAUMNkOo+hsvWUVdv8c+ACSkx3
JmoZJSpcVXGsC1/22Ksi3t/UvsstozmQ4KTwHP/TCBy3U6GG5PBtfgEkgisx2AOh8/zZVF32OObJ
c66KA1QexKTF6lii+UzH5FY926MQ1HSuZrikJxw1yFN8tWKxvSl9PQcedgZPGhC+A0W7MtbzTpW6
Th+WWp+aWFPzHr1JvoKMLiiZzN4Mo1qO1vDmK4GF1jEklxtcxA0mJIptQyIxLZx/FIY6E9Lsvt3m
fF4GuxFN9PiS4AZiN6lOBzlGAnQe3nJ9mysBmsMJtmDApSS6ZdtuVe6mcK9IlPJWKxEXWU+Mznk6
yo1bCuVCFRieDfOaclEuVrZyJG+TKOlQPODRnGB2L9rcEqIxguDBCWX8Y/d+xMiJwfD6FitHf4Ln
GKLI05rJ7cb73sBOV9RiX80hn2KN8AbUHzCOtSaFLAByS7SmA3CPNd+gclI2eOWo9XPbkHtbOQ5M
2j8/+/VIdEqg1duZJKu0foVqihEQ7OHHZKCBTiOiTbkjE6m/2Ny4dl6AwHiFNoVep+AYGElMQBhD
fnQYAy80XqLm3dlAZz2r2BGlfNrgtcsY73AZIaQMb/ll7mhN7iqB/sPQme5dpDR9uioHJO/GNTRT
YJLFwE7PkEB3ORq121X+a/8HKZrlIhN7El92RCKqWHlNUj44pHEJzIq4aH8iXMvKdoHaNERM7V/5
/43LAOHsIz7r/GLtYTKZvx/4Qp+GuvRjoZZzqO7cXblCUfn2B2EjOB0k55+32X+nBfS3tHGyuCpA
kScAcBG2s8laKlncB/CAqkDlxSdJnzBNpSBgu9TQA1lUJp4U9SQfXmJkXE0Pd06ce5ldTqIvg3cC
ZuKBBSsdilX2IUqo3ydsvfw/2wl8tAAUpwstGWoNIooqei1Q5D4AnlE1hdEJviRA2W87Rxt/K2AQ
t3AjG7dLN/vdkIH34k4eL4MzYmSKhbskT3TJWitQR+RE+INsjNr5+gIszknipIZ2gBlS2ndloo8s
18dZAiF56z5x8pPtP4Pi9H0bOTkGY06RoTD/iAPTWfOVgh00UKxm0vBt1SWLR05HDNKIMiCuVn7i
MpfUoEJXbEV8iQpKVufY9eudTccik8SywF7CBoBCfuMR1WXbexhZ8ho9M6jR5zaWdt9uCfDuwncU
2G5FdoCfuf8oKsjys4xEER9nYv1Vev/lsqxLLkMXSRB3+N/RTvvY3KR578NrPIKK0Mu/FhGn9voG
jnjRZU/z/lGKSh9IThcyBftq2f6Mc25uYpu4F/lSZA5JHPfuwNu8jc4wS/Pe1tckwADhKmjOnvc1
dC8RFJwcVaVpEhxeOsaSGWkGTjtZmdNWNGxMNpTI4Zvf8t/2uiNtzlzveIOC7XgfZXy/KMPH4gKy
CKRMGuKYT+gggZHQN7kyrZJeU+rDXS2687bKCQ0GABmbwZQfFfO2humCTAUIrJV/usH3UmtviDvd
72vOuRc/2hIcueLlc54b6aun/O5wrEmgeTDVoM9q5xc3kHnrOijUaVaL2UA6bPcLgaCd7qGdWbYt
aIOvJoWG2bFi60DvGWaDVBbc9h8tcRMoCqrwr9Ln3hEaTOd8VHXuFkBgE5xvFmgaz78gtSmaSLb7
1sa1nPfpKC/8riaVlWGdcckdBuAlrSKe523dIsKH6Xv+tQ67kjWYXn1JG7UWqqjlqiY5g22p9xR0
oASa6Mpz7uFn7arIYd5WeRd5RoxTUd7VuSzo2BeIYCr34XrIoZlwitrdH/9KGmFqywiNDQNJbPmt
R4qkfIn9Ex8vm4LQhFUeoUXjuH0/U4Wy4X2vZC6MrVKqMOAYe6kGKkgiYOgJJ4W1k3DEpeY6v1Oc
qUfc6g3XulZX1KQc86hfPmfDy52TMZAtysr6FSOmXx90CbypakWgpTVEp8BHThS7TviT8mW1SIge
vukqd6U3DlR8T8PJ0+cXYeIL1KbRx5edK5EmEZboacRYOADCKrV+WpNwtcGdf5DSQ9acTdA+/Ncm
lZZ47TDg4wa3iYUOmQJ+NvUX+aq7jaj9gqbR4mS/bTnbSlYZSc1yvUumXipl2TGe2XcFV5CTBhJ6
mycAKA+0Tm4muI0gNPRQtxy2OK3DHEGq70IQ9xJ/zV/i6G0Xd4FJulQRdisuMMC7aqlNEO6ixLyS
EzOsqOeucNdr/vdAzMxschQb1wSP0nUSjEukdpY84n1DzJ302nAbogW9ztrtt8BqcVn8b213anqJ
WFM4a1qvuwvGArylw41d/XBkvhToV1trCsQkLWgr4Nm2CoCLk9LUw6h6/qpBpXvDDwa3G4E3iTrt
gDnPxFp06MCKMFj24UZ9ZR85HXx77SszxFlEkvPXl2aQWfpHXvHpGQmRc/5E5IeDzXLUl9aWNA0G
XperOw3JTFupO87I227rd6buNTVNpVI5N6oQQ/p/v8rGKLphhriU4F5mESZX6TCWY7SgGtmSzRLe
RteAdMu9DmZRzi9raHvzj9KzLkE3bXIDltLU/F1NrFGZvzd+kkkENMzTlzydPAERUvOZu81kHEiV
6esXqcSfyAoppW26w7h+6Q5A0fsvIKdmIn7DDCORVGauwjVyVnRZihVdAA0kGVDAHbUXVq3U+2ie
NQwvTj6I/JNioL8CcXJ2cCU0nVH2D89roZfdnhk/VqTwhqOFPSkGmkrcopRXgfqdx26ke3rlnolI
m2CoTs3DM+DM9uoex6fjMKYiXbCfcbtUlIa5D/Br0dm08Vu2ZZrzaA8Ln3a8wMBSNHmlJmWXv2En
8YiKpnNgk9p0hBDpnSlCZwMA96CBF5pVk2dnqZQVSbjIkEyrx1mEkeGVMC7I36oPX1IG1cQJWWdO
8e14IX4RZesxmzQLimPavKaG0tQeSJJhW3d/2zMsfd2O3hzJ0Dx1DTP3/+Y7r+tWGv6F58cnkhMr
F6B1pOVAw6Wc2bMoAC1ZMMdeI+B/iRePPUQr2ATBmnWM4wm8awdah+zgfdC56vZX0xkUtceRV3xf
GuzmXi9vqEErDWaVeVtr+R/gyraPsbqOy0ggO+KJu6yB4z1KOxhbCYfJ7EUOPWbaZIbdD++o+IIR
UdjrHpuGM3wm8AdRB4N2PkZKgUQU6HGn3lJ+M6agdIe8uywMaRoz1LP1LjdqUuqChB3kK0no7kZF
M7udoupGl4P8xA4blHFRPFZiDeT1vGHzmX8ML8PuEQuMBXo5GyDeGji5TyhOZWZEpij7HG0Qr6T1
Db3WVMxOYyaBsUErpk4gmnFBaadgNjU4a3KFabJVjdwLltJdyC5DJYvmzFkZSlIo/mUFFJSyQy00
cDgGZedNt2SWl9xuhjf+IgQSvUi02Bzf3h2WtYhq0j2vDuU1Cm6VXJRSqJrxti91MVVGrKUiwTCk
d7rdSfrgrR0KBwqi1D2ZXn893s2PVgT4xXz9PlmNrMbjRPVJ1XZiOkDRHPoaQ76LtBdXMw5ZdQY7
fiTvHr/oFOFwfEoo9Z33HgnD6RHWuMaf0A9qLZnXGOEiCaHNSnVJnqBKOz7CKQ/P/DncqHza+W+o
NIEKdVid1viEL8yFFPpePaOQKoeyrqt2Iba+Id5o4czIAKFZVOtpMlz9m7OgdCbO54uPW1mIDy97
XfXox0M0dfGlYgMoP2O04WZ6HLRjM+McSKreUzl6pz5ZtbGf+39dKfEkR/xJ5Y82s6Ltps6ONyFP
2yxVUElYCe0raDYzTaQfxRjB/jZbWXuf/KCebnKyrrkCoRSIWFZ/jKQ4jhIIznvxQyyDSvcjOKDr
xQIw/CTkw3kb9vreBsiMzqoY+ym9vxN6JZIZg/A+My0F3yQgxhUzLO1pmEhlzQaBBgOlcMa3wwCc
sO7uohUKPEweBLf0T7P7lQF94KLDZuZHWdc+nFSbmKNqSUHQW2GEpzQWuxj33qYYXYsOKyXns9LK
0+0HT9KoBlA/LyUGJBBV2bnqQHQ3h8dwvF5g6RJxUtsTLkFgkkJwRBQL/+fi+QW2pSmHLB89Lft4
TdnyM5Lj28oFPeq0SMlj/6lmIE+BX0eleOMR4XgHswvt9hEpkE60kOjpLnCyjB/dBOjrcfTPB9R1
fQgMl/So+iFfN9DiB0bfJuHxFCegzMdvY1MLOsEGC884tqSzLxYSUivHocE/gaSH8kJ4EesldzoR
B8RG9sLtH65ucgltt68Nrtq3JIkkB2c+B2khsCIKKiGRa6j31mDTGNJr6Ucl6JPxEB92CVsqfPFS
AynP4noEkEt+CzzUvz/I/OHjiEr6tNPw16XbB2g/oFDRb5MABkAZAvr1k1f7SP7rZrzquEmqDxab
JMEKAJGGq1HPQR0UmjBhq2UdqADTnEGLvoJ4gMbiGFL4UiRNfSfzU+i702mqns/N/xeCutvuvLKI
kWGx6EPvTMXOL8S7ektN+7lEfrKNZwdaHuo6Mpg3bBSPSaD2yeGNp6ZwVMjQtx4HjtDjwGDWWJoW
prqO6A9FBtPrPSH+rmXR7xjPRA+gI3UuCITjELlPiAzFWE8rKNW9EC9IzwpiUef10Hgoak76AHnD
UDOyjmfXW5FsT4vv9bjXjEOk7hdd5fr8W+jourbbD1vpnmMgYtb/3K3P/h0jFbaNA/1OF7ZwYP7p
75nK6RDJao8er8MgE/u8iJ5nJ3Dp5RJzS49Q9E4m63878kMWN35yjNGBFmQHyk6yQiYJNeqhk9SC
JKbWXGp0KW7Rz1HiKcT8DpMhDVOK7CTogvSJL7QKWNyKBf+XEvcQ6ysADiksGNvgjXAXNlY9Ovin
C+ZCk//nYTirudGiaRynVZIxUwSdTT0oVe8ipFjtP1ZBv4sIPIqPzSsLA0hAbI/slLGWvrGmMsh+
9d7Z/M3BaHh8jvZ2ObBQD0hSmzfxk87g8Sf/7YqBzLU5qOGrRTdnMH1UydPHLTN1/bf/NAQki+eP
jdsoKmyfMakp4l1PlqbXbyBX/RWHiYJ4tm6Bd/04epQ8/BI3XPU7M8RJsz+emvL0G0e489qL7jXW
YAjg2e8vX9cCgduOBCf6wTXNa2YvUrpicM/zy/24l2vhevHVL3HIDosW7oufdIRvemC4pA6xkfyo
/K3iNo6ggwJ5hyPMkNF8YamaTWpeVufQE9MpDbWY/8fQ0h5LwlTUk1oeFAEPcifa/6U3g5w6WCOn
KUdz3U7At0yde23Tq3eNUsTf6ioaA103aBDQjz3l2w7GBElJSE9/kX0AibwjeyJ3nTxT3ImGUOFg
4mkaf6x/dEsGdTnYdYishYAVrBZWLJJvXTEGG4Fq9jG6NnBQ7dv6FWHXZddSKWTZuQP+rVF572Dh
RkDS9Gf/z3C+rwS5VDJdH/68o7YyhM4i4UBd7CH0BnyT2q9lc/OJAoMlQ9qYH2ju1oi+E5UzseUr
Erhga3c1c6Ejz/QJAAOHqi224iQZ5SH21bsAJ9qAIwho2bcPbYA86GHkXRPViM/dPkHLmExKpWQ0
MaNFNBNMi8OOp0+K2Y34PbMJ+LRSwrJxQfyAv3CVhGeISr7r66zbxin30wUHd6OznjMgSUMoF146
n5rDbx4EPyocuLyI0MY+3fQH67UgluYwMcV8PPHVox7Kii4rLY+lUu/W3ud99m4umTUtOAsDlMnQ
Q5Sc00hqI+Y8evU7vWzUa7cQxlvpNY4YpvlGqaUKiWsUKZmbauQzhL+DXJED8Ec4hF2eIx7/hYQZ
6mJduXGzJ0+5fcnIox73YylnIyQ/+kNMPTm0P/hS1vcOfRe1EThba/z50SgZSvweVfW7lZHORuZc
LMdrNpX2+b7FztG/3kQtjp5tjw5Tps/PMpqYwxrjJwi/A0YWLeX7iH63hB0Hg+mZ9TdOH2hYWMTq
IfGpEzL4T/Npc1lPKnxmsppmW6akFk0IWT46Rhx7curJEG+2JcCubUmumu2gvdiI90SsdTVbGpzT
+W7SbFHJa6G5fBHDn35nJVLIYO1ij3HjvJ5rTpqrARvIrGCSJGUv7yHzqYz43wND6SYTE+zOAsIS
A0JcFilB9x/xiFWCeL6NfpW+3KRzFTquZyIDJsJ2xEh1W6pOghaMEXbjQO78WHPxYG7R78+G+3gs
PvdI9lQbzGh/XXu/TzO7DErJTN/GmW+Rq3UwHxifvjIfmKgfXHuaORzxEEX9kUaNmIJEiQc+Uf3d
LnWpp2K2OwYQ2stu2/GwW9HHOK6mgTGsvm+bBBcPSU2EliEb5TdC0uEp/tdRYj/zLqU3c6U/wdPL
2K3JnP4B9nl1tc8HvLn6WeSXKFaHGpJT6s2lqkPRWOTuhr7XmtRPnZPJ39yCTblr5D+P9ukWrcAn
T0tVnPKg0BtVkI5Ia4Lk6oJE75NKgtbBLCaJHit0FRClherYLjNus9xR0hK0GTcSMTmO2xIYwIIa
mmQOj03Xj55n6n4fSv1XPosHGKJQ/bA+hhF3IZMV+0RaaNv+Iv95SleeLgI2mbMDB74tkIqonrut
ELCrdYg3ypoIePwT1CpvvtWNLKeQ80OWTU5tNyLLM57M64gZPVj4rSt0Ce1UxG71aJqwgmiNC6ms
cu0KPTA8qA7paKzpXONTQxSUzXQMRhCGVis9muCEXqMN+nSBMK9vTDsbe5jaN1QuJj1YOHXbrQ7u
apu3j38bCTaATDSjjnjO7h5lcmIzNxbO1gR+M1pivCYtxokPuYIAMqrugJtlTD2A/lth0tuPtDK+
Zfi7TLJpY0+Z+n/qk9rXZjD6W+YQynm/zh3w1C+7hAGSvsAGgp7AWG0vjhU1p1jHj8R/cNbSM1h8
x47Pi0LuZOX4ni1GLXZlAGXwqDjAJV8F87KD6rq29pt/sQPDnqm1ATPV+o4lLOGBdGhPx1wXIUUO
A7/q9NRSdcOfLo2oq1535+N1+wxUGGaAXab0qoEPt9UykIZKABhxVD26Cp7CWRKNds3+KECEem/t
deQN/UOOrXXVAJnhym/hRfnEmruyfV2i6ZQX1arSWQDPUE7sjAFaHeBi58y+UAu8AflOAIJVADqQ
YfAOv9z5NlWODcTsujz2Le8abN32O9chwt6g65+ZQ4sh0zePQXCEJ4kH8wRIIPElEvvXqNqXR4uU
9t0oJ0FoU+VPZjf/No/XO6oH1o7Aa+vwYzU9kPg74hNQJOkRhNXEIvZwYv9puHCaaKgHDvt+T9rw
A+/B3YPfpXQPlmfH9egCVkGYenUMtKtxyeuAmQTMLQ9+FFouovbNoMRil5825X9Q0+yuFmpziMgx
czyCOLJXHBppgpMJ4bXP6mEruK9gEuR4tnTPqME/39bi74pMSfInPs3QOQ65dHlNlTrbJtj2v/It
5huZXQhloGU1cle9edNhPrDHH4Dsal8arbQM4qfxJ0RFDlhqLe1ZivV9OoHuvMkji2J1DkVpJchQ
c4D3yEh+jnOjCITOHVVNSBSUk3m3hkJbT2KkcE1+sX2rIfzhMNrf05X0C7mdHv8/PfvM8cWkbi26
Qvtpxh6Zd6IUC6trRDOLGYr8+VZk63GqPjV8yZcqhBGxNKYXDb4dXrwPYSGDZg6FotruvVnL/ve8
067c9Ljfjhhol1cQvrY7hRGfhk27loRzS/o8fiRJg/+D1IUX0NJt+785XyO+O/hYGG7GDshhe6Mu
Z11AKuLwXGiXGPLJyzua8tNS3em0Adxw4LXGQ4oIncC2a1S9KufFO89mnWjlSNMgezy1N/E54Fwm
OnJ+EozbIbDYi63zI8TRiDz2ZlURxcsbRTJ+m/4Ofl6xtObK9Lprbw45o5Y27m0jPVgP7wNVKu0G
3y+4KtkdviMvSx6Z/2biE1xKxpscCS0C0lTby2mSbHactxa1Yz9TnJq7sOxpoL20OW00IQAsIKn+
aApqZh7QfptOdVAU18gXVWh9RTXGmjO046C1VgpO7/afkWCpD+5b8V1sFORS8vsFAOzxOCY6JRkF
v/qYW82YagvaJNPVBRB37EUtGhK5W56tF1KR+kyYTZ0CQ9hQcpC8Lt7tjsEgnb9I73ygrj2Y4HPd
q0hog9OCtKmSru6Pn/tPFYntBJ1zT5zyx9z2H+Y75Tut/AkZEHTJa/oQ/SqnzKSB6M9wlNA7VdV4
hxnwavjbF8+sBe0tKKxGllLTCFB2G+3Kd5MmdYpFFTCRyjs6fw7VitW2AaeV/U9xl1s8Ey0Nqlt/
UfCDb6HNkChJG6sDgficyxKDGYKZctLM8xqhHfgEr2pym0rE+YHu0uzmAVyPjGddpq9sBYDSl1S6
eic2qgZ9cdqWZZCgDZFyZc+2Bp24ICViq0Pvf6uCRIUjniE/m7bbHOI5Vy28ym13TmBkrqk/Ozbr
W6xwB8mn/ZUYMkrvXcT6sAp7ox+srdcrJcGh7c/f8YEYXvUdZMJoO/rmAtEx3P61abMJPAnimXMN
1WVxN7ehFQcejYic0nr8UrClXFfVxwe/C4BAa0ntudFFgdn0hrgb9fcZvU0GRaAyRyp7W1p2yHyi
+lGoB2b/LqGcxR2wZ85LgxibFyWpvu8XHkef6pAYp03+1mC/5gp7+IvGNv7v+iDBE84sIUy8it3b
EDzwh9VoImgS5iRomGkh/e2TfTCU9UPV9QjGUuWhn3JrrEP3rScuAgPG4tkL4sChwSA3oHBdQWxL
eSI8bH+l12VdZZw4grt0CueU4TouDFjU969mCipGcMCXRmlcHQMm/zNLDH1usIK9KGcuTuJCQgEE
AA2thvI19U7LnmJ0nQ2LBgJ4LbKxUGAQ8biVxkVwVHL3LdZWpZ8RqImSCKfUYC5FJ/SFS/RVjr6P
RVd/bDVjsLH4hr8dUah2TTAqBfdyYCkTHYkO5TM2MyU/GzhwsTYAVPHMyojnQ/EP5auXRY0LhCb/
IEYezrNNLHFpmrGl/GV16n07IgBXkdYbbllRvaXfIUKPA0ZpgndmJ3hyxJtLDm4BHGzxDmx8xsz0
IhvbbAO/mnqYXl0FJNZXDMsVHPipuIpKB8JHaIiWGvWG81auIXMSNwFfYnyoeW83+mGahqSVCmXv
mG67pFfALUTV2z56BVqDJotnjV9iBH+K4rIkngu5JP6J3Cfa6evAlQ0Reo3KqjAuYas5ivef4jJw
ytSqlyZm6w3p3XcY9K/ULSgeCTS+IM+wR9KrzlrKAArnRdZcysNG6daprNV1sb/xnD5pNlBURx99
NMVfRphHUheNMnYoeVTAFfyjPlyOxcYPbmG8LLW19uSF4IWhbRgoqEAaxZbxGm7dwrqPvf+YUlzk
lDdmPcn/TEwJGyrPqSOVzbQ5Q8jvFrtUhudH1gXAlBFimn52p04G3ntm/HZgNFPKrF6zSH5Zufkm
Vf9aoeXLqvkpnGYEUyTUeaxXzuxHg4l94lPHV2KiHntjhylvz1MhUP3mZqFvNkQXUdlTK0/ezO/e
oJrx+uLims4oYo+3xBo6POAddRoYALVAyJq9Qg/KpXgQzPXzE7Cvin03dnK9tIgLXnFhQZk9NUip
2TQRtCAyYvm/vb7PMHXVt+pyGeGQ9jJ8vwT4UX4mWY1Y5sWbvSFKHgIGlsvVHPuxRy/Ud0+3d1AQ
tuO9WH8Px+Bz2fqsRIowHr0OvZHu+QbACtdJwsNSLnAO37TPGc4iIa8SuGYKeJLzjHEQ+1x41aBm
owNq/PLbsC+4VkBNAVNgjpZJfclgIwFzK9MMR/NLF0ehMcvRetnTzMVvBYsvRnBaCcsOaRm6ObqS
zkrAuSvUVej2JuC2e/PWIgpdQyx+vqovU9qeTAzu/2BGCcx6UEJFWjIN6ZZpMFBdaVVBcDDm13A3
gt7+mg0pT2MwneWdX9jovxvm0lw2mtrY9O4tKbWWii4iTs6VvtsYgo4LxwgMW3ji5g+hDLAgb3/c
KQiMo4oOkrBppBcv0a1pLmo0eJI75mUR76L+wvNQ1VqOlDdJwQ4H597vnJ4ZjR5uLK73leECNKFq
9y2BhiGZHp47bYNBqA5rPlW64k3efqkeKdpEc4W4V8PKzYvLruiiEyeVcEABFgC5flkFmmxj3CY/
8EnGzv/uGGQhhXbCmRHvUpWNLqy1Ij6D2RvrMky8KvPMEfA68bxDwHJbCsW63/JWGjSSJb/vh2HP
/JCuZYAgkdwASCY6nyhBSNQqg60NixG3RhHR0ChqzFimbqnDVU/eaAWzz8dFkCKVDD088MHSgqDr
/jf2z8UkjDo2mvnhhSz0Q00LXTAMSv9S7oM0lbvum9uoq2hTXVdmdQ7tgOkX3yWwJ/TQd/t45K8/
G6zZlTSsA/nhahcamdxkneaVSMZ2WoqrbpCz4cldiVrIuILDM/U++nNGlh6/CHcybtf2+SQva6uy
ABP1TXGH/gGIeNdK6fxGGeI7pI4EuVboKDpRjWORiHK6D+wwblKOMujbzR8bLQA5pLAMkshC6riu
REVnEUu3Lw8okaHazNCe4Q/8TL5Fb1lgw2rWrN3jt81uyQvv04DaweQVzZLLY33xfnyp23WWkigH
1gcJj2OaAMqT+wnQWYGlWeAp/ZPh97C+8PInF6w0hiXAhYoVKzIFn/jZXZyFXfpbsb4ze9iphHcH
y2Du93rC9CZExhCO6I3KLGnMMRTKHyzC6BzMryWTshDTDXnzHoE1Tp0es9FDUIufULGBUFqJQk6K
csuS7FpNj8izhP4erF/7n8OqRT1dIM9X9FoOah4zb4RlTGmqG1+KXY57b4NMGawW0K+jkAy+mrGb
Gt3rkXQDcrXBlpsntnnzPfqr/EL5UYuJwwntHThZUKHJjeC4COuFGUoKCICXxQv05rR0AvXxFTGu
mgieGfNlvTWNnNWZ4+dE4IRPR7f/JUxPhKuLrWRCdn+CyuUbd4pMYP1SQgHMawdFCNA0o2xKbDQS
NeCGIHe/HTPGkWb5HAYtL1uEmqpDnpEgpeI7ZDHVu5B7JmHNHvOELxleeHze6dTyVLcVyhKZRoww
yQD8q8TtwWwhH2AnnzcSV88+i8hUAJm+Pu2GQjJcHbKn+uBzYazE9J+k+AQ6Zr31Gq5/ebUq43e5
yy9T+u03Va+EdEhTEUmwxPX1AKjxXULUTTy3ALsl+MPHcS4RSNYg+510ulQeUxZHxA89YH/R9F8E
C9W/ZlPrHMupPmqdeKvwHoXD05poVwLmNaIGmBh1uMX5fW3suouJr8+qOvL8npj5KAxcVfyCsZfI
5C9ryRCRHWg1Ei8CsMR/IksdzkDrfpZZIqD3BGrrnZmHbkiWq1ZGevj948HOry+Vvj5EBFsX8Nc+
nErq9tIcgl/IhyNDeVxEdll8Reblm9rjuZhjYFtnhh2fZ97EjZLCmtlnD/6epA7qR+qjrfmbwSkS
5477pJAOvgAyZnuSBxKl4xb+B4BPLK3WphYFkWAWyEjgUDsjG/XO4QO1iHCKF6R3CaO2vSZh6UBU
2R0LlmErD1zyBjYhUcsrIFI6AZyZIiZV4FllLrGU6kBaRm8Sf/pL4wPy4b2OWtErHos1OO7JooWR
Y6KvJ39antTYwnEGh63z1yNz8Sk8vYwmdHRfuDc5loVNN088W4FXYLpoD5Wnu5nhHsiHqQ4Yd2Xz
rkmZzrHC4M8Y3bxqnjQUCKZB1BJ0cmLNNwmqgn1pN9Gy/3pPcSkzJJ+IZiZlvxjtwmIccdspjyF0
sQH+UDBiGAkhVqWMni/fnee1BjXfo4Gq0VKJ+Yd2igSfoadRG1ir5tnSTHb8F7mAm+QwJAT2MVbW
nFXFOqKrzJwxD2efRkxN/GWmiPih1Ceuhera9OPiICggaWf7a0QXmQZR9Fj6ibZvZcW+AaKCuqD+
SEc3VrB9Mv6Q2zVIlefo58iQpxFF6kBkJLc7fTEVkTlibcrARMXOjm45C6Q2gebMzGfZEq2E9Jo6
2ZWacGM+5Ueel4SZ9JKI5EMJmZULM/B5wGkbCJHEJ82kQmZYR/EJ/bEtuO6kj4yYCotOX2voB/tX
LeVWBtgYUpZCBu+DIhMF3NMZuuSnOmcrr3aP1fhF0Rv0MKFE1ds7/34NsXwe9QOdeicxFHGemydf
+p776PdpVtTjmH2mZ+CCWwB41VO3RBwXWJm3SnvPG7wCUmWlYtihWHXceWSFJv4QUSOk/75cuLWn
MlMEPgRyELLumxcT8Pe//UZOiid8KDln2wBODq7Oz7Nu8Llh4L8cLbJJycz3oaoMbyMjvoKafMOf
3fstTuzXRnU7BDhIazZUrYPUE0aytWXeg/4Z1qtlTZ5O2Wt4UkcOvT5m/eeTdEKwBsJiNAvf7U5q
zKfooDqAOU/AmOck4TP3EOiaMuMTBa/YYWQRAkywjo2eiMY1X6TFSyHEy6Ud1oVx3c0uaSl0sDJj
vxhmysD8IMhXkYxJ5C0CV00uyBo12RZ6l3cjzweedI/Snc5rNfF7pJPSKnW8Xn2oq/SSzUQ+5S1s
6yI/qZGATFN1ntQ0I1MgLb2nAvmU0WA4xz8wR7g25JSQ2hmdnSvYDHPhLCQEjJl8NsV3ngoX4dPC
/Wuwj1Jnv8E/fYPApfv17DNuL71fHE4zz729Em0xexRlNHWMSiLoYA2Fb3j87TyYTEx6n7q+Ad8A
0js1NtT7HqUdwFhlN9hZ2XlPZl3MUidrjLyYKzqbWvgCRR2syGbDRWRq7imzFC2EK+qaSZptpAD+
wuIhHkYayjJz85v2OlbGZoc6Vbyz3BQhpMF88YWuFFolKJPR9rxr/hb9Vz31eHvcjTrQGdythJ/5
/XtikJ2TREjM/9chTJj2i77nTs5LiTAPCIhdGcz68BUVDyVud+gUQNC3qt+nvyIHxnBPjoBBOBPG
uQQhJ3NFUpLUEh+l4DI4oER94p/akZtYVDm510k0jNWHmqqsFCaB7VliTXvxc4lVwBLctt0mODDW
oUt0giYuHI2d6/m8jd/anU/fmW1iUxcue7K6HKVaKzX+izi3/ebFpJGBTJi5vFoSS0PElD+Xg9xW
FLZDV1hxFI2VQRaZZcpwn4dgVb0aeSydXrgKlM0/P1BLjz+CUmRrcCaeQLqtQmZih0mxoeZY78VJ
c7+587zoW17B0YTTthE6Srk9A0tph2yK0sSVXNsmCSfJTnljV3oS5YMTb6f5RP+GSxB2Pw9Oi1r7
T/AxQv+R4CFXpOieyx9WOH0mvCdDtoL/cpLKSztHJ9I21fK1lZexf1gA+zJ55hQXQIlh/4vFs4Ni
p/kiitMZERKrPRCJhmsKuykOuPbg3RdTqBqPo9fBC6QJAVByfnv3iqt+WMvVNO5h4dS/vArCzVvY
qedS+sHL4N4vZxPfxX7FXjCNQPS1APpZR9ZfG/LMGsRcwxjqIC3C61eDkJxT3wY1EQDp2ENy9DyR
DHn30KLkIQbbpsrvkSR+jBtXcfbXvcU1+Nmf9NzqNlvsgN0nACHS+hPVEuBgzDgAtJhHDkak5kNC
DFCCNJvALYZl8x7tVC8Zn70+HrZjG9qtJHq+PUUmiXN8YEcg9sxdOvDZ45IOUvhvc4RtRltQQC+4
GVarW2La21s4sFX3lfggjMj5hPtsxVl2lTb37r77rjzzs7r27O62k8KPdec7Dyoun91yPK+0CGSK
viBbdttGkXzJKpAbJRnqaJ62z1hpdG10ky3cxQXsBNhZLoYqAliopWTnPuXrZoqo8p74ffSV9Kbt
f5J0nnOVfrCwvhqWRD9roDrE+22XJgxcA39old2+Wpwmsc0d576K+vyOGSbs7Mroj4Uo5VN3aieC
BHATcpFToFpmAuh+JI9/HlWsBzxb7O3lGrUM3D84X8ytAIGRJ/a7/phyElAohaq0fMYi9Qx3n617
TBA+rFx/anyfDX1U75pcdt0AdqqxE0+xYOPvfc4DHGXA4wP5QJcb168h+dtSDV+35f8M9mIl/79U
hwAQ4vQBuoT4SeCNXclEMCvYR+1zDsZ2SQbeTJx4E/tHxItpxIZ12v6EjgBEK2oejwMRM1X/0Azs
kdwIP4oHXcUMVIH1wt7pHZR5y6uKeFzOOzCt/CHPjplR1q+xa2ApsiypiRWDmNNlwckpa0tqwQV9
QqRNajsfXR65tlfDrGUjNrIu3v5yO6p3zsxC6CEj9DKKRC6XYg8jOSlgKjbUngWkbkozg4pxqtu7
qcTKtuJkoGRE4pYThuOHzT9hu63SEk4QSgFkGhT9nfrqbUyC7l4Ufh7mAqfdJQzAmk3Icu39Vc4D
vbqlsqNF5eF7hlprOCfKjuMLFC3EXm+Q5ByKZihI3xHujbCrfd8GSQA32fo1Z/GJCB1BgBOgOtD+
EEzYumrBo7GlOmm2dBIYHllEmnGnWtxUjCOrCmrfqqL76iKoC4+61kDGR9tTzkS4GJSGgcpIZkwn
mRFwZHYjbXc3YxnO14pMiZ/uvQCvhdv+kwdUeCb/mPF28pNsd3DBBovwlDeXoM1a/8yzb2LSPTGQ
NyYI1wZHPkBUB90VUOxPTD//WpEYky3WlSPw64ybRa6oYY+G3sNzKrGnd0E69su2Cai7mapkBe7z
Xz6rk78ki9bn0SPlHjc8LnXgsw2VPr3+BYiyfLJq8v77vs5wJRgi5Rl3HUa1BGukixKHOMf7H5rd
06tWgU1bd26BgKpSvp8VLUvnipPCGbcBnJW+om5H3OSuuboOnfMNhqK3IJXO5mcUDT0/iAJRSyw1
QyfYtpzlRzrCvvg0lsDFVfJ0lKAaUwAqoIGbfmB+q49LU1m1kH0tiEjbtceriPe61PZAyLY28z8H
CNY/VDoTfPzUuwmFXSxwh68XaqEu4cAAugC50sGOBYXp/IjOrFnv24He01pvkjZbwXZTjc+ikZ63
Cht2JXe2SfvpwKRViiESSxErdBFTHZLCAvTAFNheeMkCgYELfksawSZO75uAhfp6VcutBdwkTahx
ARaQwOQRYX72xkYVHs0P7fbU5LZ79OJ41wwe2SVZ1HoyYE0tl9/eLB8zNrS5EpJQNQBgqC2WnmPR
a+elA/sWAsKZ3dOnYixlQcD2RnjIxX8ZD2BouDpTS+SS7TBh6fWl5SWlG6EnwI3DJx3h/sjrhwIb
lsjjMSO+PHx0ka1oo2quh/cEv9kUN0Fz8wxfw62DIT9NpOClakv9HjNylIYHjQP7Cln5/7hHlcRx
PdYI1fpRq0Du89fdQEYPsGfYJT2FA5Mf1lEQYA26LFqA9rP88GP1uLd4M2ZBTVlxsceW3BM/NB/T
oLGkJhFrvay6dU6HLn/hQc8ntvlNFODNwID3ksmsX5o1+2Z3nFoc5kcwC4d98BX5L7QK2Ef3Rflh
cMNo8oTXbzu2hwNLWEyiX2LzgfRbxHuDxe4RJFBwlve2RHdvJDVXfxtQBT3HvrErCwiuS8h/NxXD
0jMR8AJc8ZZRM+BqsQIhwAZlIEdJa5G71aEf3kafNhyz/H8ZxSksjN/FtsVYX21MPn5s3ajO5Bta
JlLnc9A7zTkb08wPj3VbFHlFDL1mZuzZ+Z2wfuHYF+Krx6MYoWi8VgYY6rpb5tZJIHHznrDgijbi
ns4OX/7t1QXezQ54AmvsyVnsM8x48EJlGXZEkkuVpdr9sGVKuQ67SmH9Er4VMePhgMVK170wbonT
H1ARVEHqsY09nVnvrosMftN3DObYrZmIHuWZqcIZuIMuelWlATUqRhxpu7gzdQUEJpAPtEFTDmCp
KHqDes7PntLohMBdJBlIwhLrVFv1ctymj4mXVYb5FlyNTYngmYCwCDalzf6J+gdbcUhnVzX55W7J
OxN62FK1rOmrdllBDxTJeg5jfg14IfY3k5mpdeztz8XF2PiCXLYRqUQN8aRijNbbRJtLivxPR6QK
DxqOy2s7JzSuOlWoXIN9Oc1wh/WmPCgV0DqaPYgVmHg3tGXy3hvGt6p619eDVdTWIgrLo+TcOnII
qXZaDmeFeExyNllonPyu+txvVvB/J52tQOOGlwvOJhsFkYAMna8UPQbacWxPbnhZwG9+e/ualOql
Uq6afej9cqRJKvxeuyCN4w2Rqn0APho0jdirxhXZK1bOITg5dhDsSaNI69KNvgXfhLfbJwH/CmkS
OtmcjaVTfXjqTYErP9aok7R6CQWphTVMFFoAr4qT4z+PDThb0luhI3jtKPzXgM+cfR2G9dc5Dg39
zpabQHOE6rRoZ/31J0+ejhmeYzuuErfdN2YfTaydEXpz2J6VhqaCM1+BZZynA8IlFAGbZGHZqJaq
VSebmRXwbKeG0NQVCLFxulhNypxKdrt1Kqzv5/WBs+quXVNBAdGhSBH/Gf/dCspie7Ti9v22bjtR
zhXNMw9AFyjqpDgiK1Ub8Q+2+qnebJjoROdPQ97AT4ovkbQmI9EUiMH0+wRaGkKHHWDYm/+pI4pc
jEAmxJozXKqtyDT2sicqnARCMZ3SMx+PEDY8q80ve6Nx24L9nIPxUM0SC1/Gp/ENRtn0yQp8r62V
YYpsw0QHB0Cdex/julAtR9ZOu1jy3AbS66i4caD7RYrvli63msimAf1blAebhE/eNUETrUvWhm9S
g3foHrKewk8RWta9eZtT/5SVP6eqvadeXgxRjVeeqsWYGzzN57CseWHgnQOgPw94/MKxlbNWlde3
7Rp/bLidWwRReN1LAS1FQ90t1u/kXmsSCjoSakMSuMfhwYYZV5t2hil2CAwXx9E/5NfxpMIockq1
4YbNM/lnM0V2jZZA7CPLTtz42ZEFB2J6fRbuWIkdnGN1x0cVH4r5b+vpJp9z7zYo4y2RsE5ToxlZ
aFU0V9i2nk0S21KxGqZEbty8PJplgMkaJMsEOjWuVl5uBkZJJ3342hZgS7LiaxcGK4vfNQSYJFgf
lsBkIfXPyxurhBle75iRwQ+zlUy89beztLH/dTrsRmGV/SaIw9EyrNsg4Aw9xybVlVUbiSIHWqAX
q7uIojmIG4TI5PFlb/j9iSYeq55Gz7QXsbHHZB1ZbpANWmOxQZfS/YSbhdKSihsASTvGd5nttg+y
duxK0W7K4MMjh4gdkp9PCfXt/EPPZaa6zrlDk4K0uBnZh0pWLTu+gJIsnKRCdp0yxrUODiArp24p
IyswkipRk2odkPpxfM/BhWRMqSuAMmacMXC9SB0X+OsAwjXb6eblp8pqeAiouYv551FMOs+K+LFH
Uq/IoQiY3xAJg9Bld7c0H/hMEzrWbuobB7oAmNPIazBW37tRDrEmp0FIjsbZx/3RUVVHqbRGpzDS
DGlIpN8uM+1DpkwghShF4cQfZ2PlKTKi1Bp1NHuE1ExOaZAvm6QKL6CkujW6y67lKwhxs/UeJDUZ
HAgDwvM133tmlt+M2PyyAr3bNgU4F2MvjPZAAYn4Fwfi/IhwwdTsBMg0ywj63Y8bKkRBBz7lCBai
JSWXmeriKqWL7e8AuQ/PFDgQNphX3bqiGABIgrUyQAr3UBqMCeZK+vIh/1W/y1Uv7v+fepVx2ppH
FTv1jHWUWjm8VBA4+4r7vY69ict8mpN1qggITjGX0luwzXiblbZpnqBpp+DpB+65ztsmvVtyCILo
EuAdMopgKXfNc0Umzm3OQ7ubis0dTnlw6HHAenVagcV/XOlZJONAghzQFuIsNdykQ9HZYRQ5MsLw
lHK3f4rUJOxYqWxwkwtopII2dNfmCxy4sIejVRP7k/OBIHyQ9B/ei7ag34xZ90IYareLFm7QQa9A
bhTHpteoObY2QMxH81wuJGy9oJaHxA8fomA3znRmWlaK4yxYznusViH0B4vY1nr1xa9HX9OSHkhM
coASowRA4GkCAUAGjC6VYw6MVlEBEqEUKNi8cXTWUW8txkSxuhTByUU8DeB7Se5pkpTWDvpMfj1D
Zh/VpvJBBZi38a0uPbOFkt0Qy4H9+BDW5hLe5W9vgZ3uE0Ihhd4H1MFSY3hEJ2osUqvVfnNnJiwu
0V9O1RHIEVMgc87+agk4GV9VhO0bvS6TAwY4nBJLxqYIP3qk2Pn9BQLdD0t0+Na4xxhtuBn8TbpE
lfWc7Sk2kTgjqcfnOjEoO1gSdc9sMDPOABPp2dMlPbGlH+m3KQasFiRQvuM9CWIGDYlDiyjSr5Yv
mqsJnfa6/CpUrhPL7H4iGzi4RQXMyWGG41iPLWWkCAEONVlC5rVT1bkIfOjFy+F9lq90F0DNfJD2
uF8UQT2+PP1OssVKNfM3FhybbARBedVxWGim1ZU5qHH4vKowH4j0MWx6Do9mmkIYLzFivkhXsEpU
CDNv+13LuKBJajRUdxeRJdbi1MbO20OGEzdSlILCgUp66kfCRKtbHrdBx0/oqnJ6dm6qEooPFfSE
rGdb/OcE3tT1nco5XI28vu5avd3gpojNh6Mci+U+B2GgOCiDBDIlZuNp3hvc7OthHlpKkS1CBGQ9
NAOd9NAL4HnW4ow/6fFXIK2PPKjHbBLa/ptdhlDzCnTv+/GeBKzmtr+9J0qF4igoP6z1cF0kavoo
B4KXKEE6V4KKNUwI7AqmLptu8Ep26Py45L76Lpht7px93oHIJ/cWQuTJ4de5LaeRyjnRLqD+PG+Z
y6eP6OAB+4lLaTbQW4Mm7c6OBGnk+ECKhhPjo1W2oZx6rn32y9eJudN4u+5izRwZ7u3lpr+63EvI
ulE9Uwuk+3+M1cjkTfYGKY0EvTf57PcFw1DfrTfCped5xhuWsBN0nz4wd3PNbL1xHnpFx1LHYGCt
+4O4EB79himSciZ2hKE5e0X1gmtEtAs7kpweDJm1iDqR9QJ9b6990nU3wUY+jCymyIbK+auD9DBb
BEIKjjjGV7mCmSOoPuOstL4N8KRz6OKlZE4tiLJyeUIAymK2kN8SXAgL9I1kO8xMUtpIHoNrj7lf
dMTWPomKVdG+TTofH0DIkCBTo7f/ORF1wl1ky2iu0fB3JTiPIMEWyjPrJjgXHjstJXi5rqOP/7bM
gwjxj6dHs+NU3bPIKf4VOzfpf8fHYIep+oYfj14FQTYTt6UuWuO3W3lVIpySbXOq1gJ7sczLKhn8
Z/+k7dciu1xWTPcG49cM9pIKjP/ZZVTbVFGi1ItvUYHEq0SJT16ZYXDXYjprfNjw+DV4kqci41bA
hrtOQVvKbM/DTY8offgHF0NNOrbJClI2EaEhY9sfFCWqWEUZJhVwNZpoM5hU7lyilJhvSWafI6++
GTh+72AZFAsfGy/lHTdF1nioC3Bey3lpGHz9R1JTcklpVWxDEyuz51ogyxlnMt1LBqV5l7w14oXi
aydeVxsASnL7hIxZgjMW73U4tdDNuciuOCcCIOp1/Oot7CszvOx9l4O69tmlow0DhmcqzXvTRbhQ
NPX+L4ka76DwWDP/G5eZ15e+QnIjfpZhDb174tjdOdb5//ESXOEtpC5FH7VaoEewxxdazBQf2t9k
bBwSEc8J7vZzRU/Dj0b65idIXDKqGNu9EKdWElEvVUj9uky7N3oBMKcf8vNRWX2DYmwD6qjEJdZ3
MSzvp3wvfpWOBiWMmHvb5UK2QUa35TR2JL3A9Y/sueMditH0hdVadesN3+oXDsBeWFi8fD8bTHbR
E2vp52xMXJa3I/HB4uxr3CHDmU+HkveEldPRhx8ddIKbUGBgz7uXXB6uyIuElf48DSKwH5lXnxt2
P0wVXaV3r6N4Am0N0OQUnbSRKZsMbskhmiegWhxeF08TPH17KO9lfyMeOa5Vk4tF4G7/FwoKPZqo
TyZhdCbSg2wvuvyTOvuZAP6SyMchztu0xWfXEBoDRLiJ4GNrR7rfK4o51w0qT3x4NUAyHzRyXEi/
2lcNLjnc+5Eypma0KcLrkbBPF2KqC4rzLEAdmyMYu+gtHX1AMfEEVYcUgOfwyONbkBBghLfoZrc8
oFFLAU9g/LSvhnH7an7268TWPPd64dcZlRJHX8h/ORswvB2n4t7XauKsZlFJcRjEyzGLzcapk5rm
SsmRkuZ/zsueJsOeyyk0czPxBUbxkNJ+U8VzNtYrKASJGMPVhvsEr0/P35vcGKMJd7tDEd/keK4g
9Yc5nNkx96er5R7D+Bxb80g/EEUzkp8A3n3apLgnURgrsegumo+oJjtK611A2HNg3KPrlMJbJyzg
YAdN/Jr9x91fnVtyiWzTTg4ai57sWb5/l8NwMBX/X842GDyWCCUG7JdvT0w3ILNkGdr6qs6jeOkE
J2bVdiFfQKq1rO7L+cKaAQubZDVJ+RChrU3WRowpKQwNZq1AiQH0kpeQ9C2Qny9opDLH6S6oxVxX
rzOFJz0u90OQozrSfVT9rXO+0u/4hPs49ib9Jc1S5/QsT2r1sW+R+PY38e5bYW0CsBruU3E/IsQT
Ps9lLG9gjsShWSof27oiYdVtv4LeVEJp7gLG/Jpnr3BGDJUkrf+yVamMU/4M/YIvJeWexMePpj+O
DnIG4mO3IFr47ftHkuXJxpRK1X7h5HvMq+DAOBVsIYvXLt7ohbSgp3kGnhAK5HoyLtJN2ROCpd/q
iFHd/IKByfzpww14Bo2qZjaMKkFlBdkf3tmTJiU5dLwW+fEigecO0wz8Nt+yE+KoeSg+8RQfAtR7
GhwgN3mGFkEPac4EkLxpJsCd82tv+C61tzhOK8WwvrpG1aBAR3aDaaBncCV7qlpZQfTPpfOUnrfp
GAoo2k/K/Fqfe1mFZrZ9MXir0az8VDKeMaWV/6txfLD6WimXpdYFKdm0N5Zw00/eE3qMZ27Zl78T
4OPevEWw7xaL7yQK53hFnEnhnhT0GBn+TJftEKFNEuhigpj64T5b7i+s3lWWMkboDqnkeqal11uy
TEQhkO64edzTxPNpsHLnXlabuqClUmNS6i8De3/252Wkmi13MvC+Lq/+zNAna39EuZK5Yf37cHBH
Oq4GIU1sJy6mL5003UG8bzwCBUkqR+nguHAJOE/ZnW7n2ggGsvdxf3zzWf9SW1TSnDNmwFNQLHQo
7W+PPnwCFVxQGCqTrsSPvDg4iv7vj520WArdgG8Mh+oeASJkFnzugbvtoR7QQ1zuqDOLtaFpAJEx
P08QXODfLI+aNbuPe74oWGPTgcrm+okwtlBOy9MgcNlPEl+bWkD+QZK25hNmxqNjEmrs2Q7zSje9
UN2wlxeg78nv1kiZ2S618hGwLU/0LRjYa+g5nNEXmqQ0p/l6yuyHEVbuYndjtKsCz5Fzp44ECs6t
yfU9CLMwBVibG+iYSyi0hACEXoepO71rWVI6ljbnmHxRb+pmVE7akjIVZeKbuwwHMpCBgTFn5lSY
VQG/CCPMEU5jqZYljjz/lcWdlwlHuwhK4cXMscgq+2e3jkQB1XMj/HWUZBbNzhC9SZ83VMTSa9zn
SYnRTKTfzFrqsbtN/L39oIz5h/43MwJ7zrlx1LvR2h5LdSFK3U5g4zmf6CjWrAMEu5pYBgOwj/zX
fNxxgrruZDsWfSomRFOEG+U+wxe0lLDIsqu6yrh+umDgei3wfJa3CGI5bwjshlBI0jZ9S0EPZBJp
rlmAtKRZULi2iIliCOGlcm+by4vo8C2xH+l+auH6AmCnS0RW+uymn4Uk/+BR5KKW4GQFzVGcFdq0
Q97OEhuyG02KDa1tLKod/FYg4pxYS9EIBH1yt9+P5wHQchYBiPIdM+XFE5OAIDCtEq5QJ0UFddZh
IrfkCeBQEteYs3Oj/Qct5K2c7y290pxvM6Zmcoy35FdFly6g2YrGmWJJ7vlsTGFhTKapyZKeHh/N
/rnApVmEHU566cYp6hwoM02gN8stgj/Bx6CoX8vfU13DyyggsmKTF2Ms0JmBN1zAiyc4Euo2otHV
yzeNkDDAwFQKB5oFsZRw8ADLImQnLttGnQgFF02emCtP+h6aub5ZQmT+9S6GQMXNbLv+/n5C+9WZ
bxs+Fkd7ydjdfKgAVeEy1lpJSXpKczcjeqj8pQnHYJXl1phAKjpczDZJU9Xh/Y5v/GohlNuFrPjT
wfXiH5cZJiUIsnPmGlMh5cagde+Yo9jwb1ezs/pYDDQYjSU+mai8TfT1j08FHAWq3YC4gf9TAokW
zo789uFcBqF5kZ6GX0U3ak9xBDjMP4OPYMBkRpXplmH7VvUm9lLhcunua2xLxX/aMmHFwXH8krqE
5SZ4mbMftE77rsd9Ud9UubzHpwc5sXFjqBpZcwc/zaLSKhJY5Vw4sD/p8Aem80cmMFZGLFCv0x5m
NTYZF1mKPAA1N9G6XjRdx+/02IizkOu25onAeHFfD5Y5HnFy6Si7R0uKVlZtNxqTHLKJRLPqSunq
BSI9SYAoYE5afKSsBXxSOo0YSArEslhmZPoevor4Arl2S5/H+CkOTget/vqDd+kM+O3lEwqz4iRF
SIZJhVstfw8LKk6+eBeV4jlCKocq0QM85XwUUPr73zTZM9ipoGfgg5KuLPk//vhtaWor+/ScCcWi
px+AhNNj/vcBhGF0z+lxEWGMXzdkFJHNz+08Rr1OQ2tfeSvSF9LY10yXDSj5jaUfe2isN0SiUblj
sxZPlmEkQ8yULp4e/TiXcdRDd62A0H5m6ncSqBorw43EtIEItDl1GTFPOW2MxoAgfXkScB/SQ/xc
ls3xymG8mTiQFDgM+lteE3GLtfTkOhJVh/t7/7bLZoC0bwXst4ZUi9mlSEozTdFvUl3IY0LAeYlR
fptEzIFalhiiKWy+XoVk12VRf7KH5236dS7jRtcaie02/W/FUU/a5cqicouRy/1JmPw2SGmiAjCa
otGGjlggYF3mKT5IrnyUZv+ByKeyVzyewwDf7uGnFhnmkobFrM9K5MoS0jrN66ZxOCef6MGLG9sR
7y6z+CZYdkEuGg57yuhW6Buo8a8Iwrs3MzH8fUnPHWqWGL6zAJQeeWxw2aEBlwV5XaBQCEdX546/
68nBHKQKY+no2APDcows6msHHVb4BYe620oAEV4cEoZPOVKSLWbNkStNWrSHeOfT6I/n7ogQfafi
DEvh8i0FmS1BU20KrsPWSEJNyPnN4wf27+MdEk0rGdxkEEizq+a39H8dqDGlu+PmFjObzG1sbO9S
hxNdGP4kuOgFFSs2dZya2IVPEQxum8xAyn0djmQNuGWFISQahggocqdES132eTHw0u6FUGArV+k7
wzAZgNg+qqMLGqtoJMcatPiNM0exjNP484mgHv07c9q44p0pHcQyHeS1LFUWiV2HHoqeXJg9S3d5
hKoUSRFea23KQdbyy2jvSvHlRRx59agwgFAPVDK4iTQd3J3pPrE4qW3p4ogPuq/XruLHKiqM1i+Q
kNffkYKBji5+9WFnGv1GJQRvkeXtj/JTGywcVJiw9nEVgcKYpwh+sXDE7sFLGQRJRCYP5PxTC6iM
QkZ7d+Tn7yJXOdmR/9aBtzNwSFkHdkT3MDGpUF7yNCfmcOYURzoG+dUAmCfBkwoTO7KmDXpXjuw3
Wc+3DQn5eAoK8mNuu3o0kheIXpq3MWXu8L2tV9cylNREMs0JYRazbrixQJ0BLzshHMfv6IbfF+rk
2xXKZEIJjZgEIlTQOTLAwj4uD1xhce2UtDuv3rS8/hmHZoaGOdJB9Nk/hoMmafiAdVYoOQIWBD+Y
OP0sAOPSxGyBo/PjrRV9adI2oqREJI65+RL4JM6efjla4ueR5IgkkrQVo4J+ZanHT/bB9qU6h445
gFoEsrq6LQQMVI9vUXItMhk8Qaqwbgcel2+NrIEZ43klhhvlxJGzpzhoCMnUuhtG0cL09BHopvh0
QznDuIMWnTK/ftzoznMNF9RrVrfbvQbuXZaEs/0LmqW0lGUyx4iJLgvCdml13Gchp3LiysgIOoiA
1HfDFLZmjTM9S7nSynV7DtcV4EWNSNmgd19L0mAmXrrGNrsa8tCIuIHW+DaeM0pShJyIlQXykf8D
ScyNTQeNcsxmpeXrJxguheQpuRFRgnSRfm3x6HCVOBNSrKCnKg6NUPYa3aL+SOwZrhvRjm6DP5Ps
CmxkRGFX0D2ysbPtFpuaugGBm5A2ftR2G6RzdGldxS1NOFY/NWJs31i/pPcJz3FbN4F4mSB7stCB
qsbyvIBk55DTSz/bXy79O1UkBXvNGOxl0mrHY9SV3EQ9G7J3QwgcDuLlY327WP1IUo/DAONzbveQ
R6nLccbeJ5WBGCZAZrTgyOxv7BCXgfgZ5racNRPvPmm+Z+3NMs3zuwh/XH9p3Mh3/lIxLTgceDO9
2DsUsyPt7iqMbPj3cEelkTTO0ZbFHmcjX2+mxGP/ENkEYF1dy5anddDFjHkthPr3ynaMgPLpyrWJ
K9f7HBtH1TZOh0sx+H8v6hMNijCpXQHLVnIvTtpifn4o6cnYhUzsuUo3JZyE2zutKstEgKhZ/F8c
TxuZl661IbedI5NB6k0sXGdMrfWn7cveSx+exc8EtcEfwf5WirkSKNu5Hfbn7XvoXZZOUIjE+YMN
cUkmN4mhLZElff6T3a6OvYz72P/syoeIdoTMVGmPb+lmAnv2uljjVWBVxfE8EQhrD5M21/3LkcA0
G9tm5wv1tsa8b6uzpf91e4nPlDhKe7yM/rXPpMTq8RINXNlMrMCC6f0uy8pGpCztUfk0B3uT0VUV
bNAxebfQz4asVbHB0J0jt70+TmfWMZqUueA9h7Jdt4knYJrAN2WRD4igTI0W1tAnLetZHaEJXDYp
4TBq27QkPrtFg4HxiIZH3W6S6ACVO9UxYCpor911x+OsxOK9Mz0xmMvdYibqGXWJrh1eprzyxz66
6c2iLwA1JfEPwnw2ZrQXFQ4vGrovx+aNjD6rVpg5+uEdcIiA2MtPgM7/am2jh6xh+uvqEdZaC5RL
rltKvs52kkc789d6VCEsXH/b5q2ugWvDDswcT06efc0uzq9ZkQnXBybXQ6t7JAH1AcXStLD2sifM
oQHYga5vQFArLBxhwwUj5uDqZ5vFmHVpUkH1uvWH6Jipa5VTz3DTwMmgV1fu/sLz+AN/16D7iLCs
wUHdJ9uNtEq/xk7Tr4hqGQEdxe9y9+ibXyJiCEeNT6D8vLyH056Ky4i7Ka+e0Qhff+b7f/nyn8L6
J8EUQ6Gm1QhTjrwnIP09GCyPtskv30uOxDchjsD2z2aslQaF2Zsc6eWIsJs2wkcb3gUHgZ9NeAqu
Cd20ztUWwADvwf1PmEzDEQKOap5Gczr0xPT3aPjn2+LRyab6vdzMdam7+EXFOaxoG1t0Xp8GdqGa
kac7JwaEaPKqd0/fnJi2T7f51WPhgzDHSWDfKsEF+tU6X68UmG3s+Cc93hkqH3/pdCGDDXA+Yyoc
yhH+TXUBqxU70cGxIEyWbhh2LOWwsR3nk/PYK6NuVHJ0axk8wNZy9+HlWXvFKQ/69NPOedPvJ4xU
LLYOvCdOh6zVimy2kwAJuMcyOHIgMcdRiCYmJEQuJwC3dJNhUwtH8nLiMwtgE1Vj0Jf1RkHjEBSC
hkM6BUedf8heHZYophM4LrzzAA7zLGhQLEZlwK8Diuhzmve3EMNNU4J0/mcs2GYiyen3Lwq7Qf6+
hcsVzuZjp5jY5qvNTTMaO4+Qh0u3VVY6tjS3r1HRdT8fBsgMVKvUsrk4K8LUoNbnyP2Y9UsNAlPa
6tI7d9QIvE7NP0fKrf3eSqQfaaldtUbdIZEwknMe8kQ2DZV87B7xZjazALo3m8ZYRRskx5/A4qqi
qv2ghhd3D7cB/JzsqBqxtMnVbJfP4WSW9EHKe6FHIrhMyZu8MJ5/xr8NcCz0Vdv9vr1RoFg8EnhR
6epWP8Oxkf8nVAcNu+xWMib+DlOKKpBlwqbdG8l99xabrkCRvjtNmN0QJu6Y7ANtW3j6ZJe/VlCa
+SrOdImFqQ/GYVF/4q2InDVmceYmK4mudCFqJnjI/CHug6O9s/tQtlGblSJX6MMYiN2Q8bSID7fk
XWCN+2RTjd4RT3RA4jmt71A2Al12+ljf2eUnGl+S+QM13rXdSZEjgZPgYKHGXkX9605M3xVNDB9H
ji8IpO25L0A/mS5Ef+vx/5wlhRmVzjlwZU3T6ru/dRhVJNyMOqHushJOCrO7yjPgCHrmdvyC/cKW
bT5WCm5UVghrH7cgJwBjKRwjQpUlPk2HR8Zg0eaMVgm9jRnP6iej9VFkc2EDgd5rer5ZPrcIjvgX
6QKgp4KmyvPQws807GwCKBTCyiCW7J8aK4+6SOdPkqebDw/4ZvmUVjCqATyNFhhTo964MipdZgvm
/wSPeQyWsLKIl8fJWK33qwKvT1pNuny+n03uklkqZlon0oGiYvA856aHpmpZr/x+G6F+wgG0W5Yw
JS4+ym9Sqsilr9uKWuau2RJSZsCoQcOipKZhSWZS7lbrr0ddSdOierDoFZKC86RGpJ4fUmzFdsVb
rdaAV0RAMv3syv9E5AhxyWBYqTFUeBC3hi4wVPQH1T20j9xuVqzrxThJWY0vz8Lu7E0fmTzfagaZ
JsnsZLAg7ms1MxHz/4V5SRvd1J2bwo0SRHNk+wCdIj/cr2p5RFxXuvRUOwRsAsPI5lZoOfMJufFt
v4UDBQCQEYnyHBzRVdAgSIJgEW4fj1AdSikKCE/ACVfP+341MrfuNhZ2sSr6v3vhBjaZRZeJxh3Z
gZoIxFEr6TaB3Q0XFKGY0VxarZ+ArlP/FMDBGI4EviE0cMLFN9njun7c6waDFoyjHd3hDdASnkmA
2J5e/XY4XrigLDWUs9h1PNNbM2GM8QLyyKXx2RFCfajHGa8kBRHYN9ZL5IekQzRSWETmgayEJxz9
BNeNNTycxkDWotahwATaLGzUJt+oFZFqygsvabErBDTQ3G3rY1GYf9PZNE4iRIz5BLDMP7mQkjEg
mMR9NCXhwnFKPmrQaQSIKawmS2RjgtCd3J5E7qJJH2WWrxFQQx+6ThMLYd0jQXszRQfBz9/x0jzr
AlFx5FIR/qIq5FqyXJyMTpDwvc/dnh6SFXIpoZsZJhl8VHZ5J0mD8j4gZcQ9COA6G79NMYSYjFsk
cHjUSmG97EA7PQtEIc2Hq5eQ/5ZG6N7E73nlJC7Iz7w8PgRn7R/nOc3r5LDBqalGy/xPViqpHwaZ
A6lQ9wpQd9uXlU6mvQAnj1SIMaE0P7aJvYBksYjyrOND+4mYJSXaOJnStLQPB6QCFSzrRoV7Qscq
k9iHLHQdLGAaATcrIihGJISzfA7KYMn++svpWKKQP1h/66N3wLgLbF9Iy7+Hz2exWiqzSuvCREH/
UyT/9Xm/YLd6i2xnPpjpxKn1wZ6ryiu7UgwpPw3xwbWUw5S6rxe5le5gnJlZZWqnHPkwzItEB/HS
bNge/HoOFMEVfzdyLQiu07U6NGRcRsaOFsS/ElgstTqZJi+DbnZAyfzFXdlgcp0eF3jdKTF2m4+w
nJDt+GxlNhp9GQ7llxMrYpvVS6NXCxneyLre4tnJ30wx88FTN512DaJC4pmG1hZte3CL+kMXUk6t
igQQ601cMW4Ffac/nc7VMPOgRqjdsoJ6tqcFDgGN25UyolWdn+VhHFzYIGjwx8OqxGRygZ0QkIxA
4rxLa5t3dNpN3NXps8nDGnLII/IA2bERt/jClUSythPTgPiLmtVpO30RuRFAvk6Vu+/OQ3nU7JDk
mlmpPZ8SghuDneY7zFoV0PwHB8lsYjp1XEwrOM1ESbWf497lcSjcc2mRKqr8KAyFf1A3Zl116B8I
V1WKubwT966PkA/UWwzrr7nPOwLS3cIMWQpz1Zv1MSIt8FxzDqqvcVL4s3Ef7nKtNF/8iMwiOrRB
sjdPQvwg+JTPhMvDMzoZGF4hCApKpbc0kYzukRsFIrLlN5RU7x62X5jDl17uhIg3EXvq8MIjW30U
3HEjkhCuUDC0kx5OGh0lOhOh2U+5j3ncYDKsys3GSlHu0qc2T5OQ7Teg2tKIOGvdie/9cr/fyj18
GS0/hShAbpx25h78jMV+kC75UfNAkqtm0px8bFAjlpieJbnGohvasxhZIPKsZELuCWKIHjNkYbt/
WbRaINO8O8TO2asThJ+c0h6CSQ0mL2cknQ+wr9o7JFheoOJcqwb1j8kUsrZc9dJq+BeKR94ST3p2
HYFE6AXv4RVXcGpvYfD+x31kmASijNwTFuzdyxUK03kG+9OD4654tMGVQT/HSoZekHEUj7jmIE1r
l3aH86nAH1Y296iKr8N2qxBVLLnv0MP5cTfRjXSseyE/KsGolA6L/X13/+0jgMW3Lqoop7NOs3EM
UuCIRU+leM1kQhXUPXLgTuDXjQcop49ZMWxxRIXweV+7gdc9tHuWBQqnVYsspNl5iNDslIbEepdQ
79jrY8YzK9BT75H4hHTM5NHE7UsJpEDTq4mKa1FRTGADlmHZW2o4qgyYrUQf8aG9Mi1W96XzyRkO
3/84KbaYPlGWaO2/UfhN2befJZi9SUdEij04+bSM7qu9VW1bDVOqi5vSKWv/ZxWUSybdkq9ktCyC
OZIcCNxi/0l16YeF7oqI8sEZ5QHeB0145ZiMnH/tjZp+Wl7s2v499mQXKokUNXjpM/c/8Qu98CP+
spAH5ze0H4EbfeL5cIjn0QdeiWw4pTrzPrERcIVin7XGJByxd7jKjWR9duF94NpehOKBHI0ToI2C
OS5OBJdkAPGH1K8mr351Ml+kPune580b9Tlqx3VgSW59ebbdXpZUXuj5sbNLNIlRhyqophDNeI+S
qIAMMKI+TIe/QvGWe+XKD1ntOWc/Oxe3H4vFZMfcyOJPuuwb1QFIiNb0UcnZGEJjJn13slxWz/Jv
8Laj66fsdT/p6qJpxqjX8COTT8oncCw0swUlveDxSsCovwU2WzXBm/QRqHfEk4l+G5otbPzOtKUy
n01rHDve2ugLXB52Wn8xYe4U9ecpREbpEI3cab4wkjd/ZpMqxwjsCoDG6uOCAbCvZjtPCMGoVc29
rx0UTpbfydBiRlCAXIW7gUCBRH8+ZxSEdZnmsz2979PpNq0+8Ld94vrGgrTSucnZiim/j3zgK8/5
tZKIKaAM4Cnb8qrXzgz64f7d1C1VQ4YrpgkK90GwDziseR1MiZac6qvfWF//iauUa81fbyAtkZd9
eirrp+3IMrUg8lEkxq6birj6uEZkm46sa2WiDb1OqOnmEkV7gBa6VQBkgDm0JHVyBHqxOTwzMttf
lZb/ZPGof2ACj4tvkVRhpEeAu9HT+ekBhZnL3/tSWYYL/uiHrvj4pNtWS6sRqIWt/0jJS7XTCDRB
Eb2CAQXO23JZTPrEbsNq1JsoYn+8CUZTjL3sBgHru7W2zN9x2FS5TdzYgPve9YQOZfWJLRy7gh6j
RHL0u8olWPnWaUsXLlO77jXjHJkycWSYk02Pdxmb4Cz48l50cYt9+Jv5b3H8FyJonLqSTqATXdd5
8mjIGyNLlVpz2mtPUlsoUd8jP2Q+Oob7H+uXu4xR9mITjUK0rAx3eWn3nn9PItuNSGIxLRFQAncm
8UZN2AVGvQgTNdQVgEpuizMfgn8zzSxMn9JhQnGARjE69cbSaP+xi70Btf4833t4nVMM4PnaWxAB
3sx5N6JdmzWo5HxhdfNf6lqDZO6U2P3rfYSycJByO8D4i3CYSPgICTjjoI2nixMnhUfeRq1NH+Sh
G/IJP14mTQOeOPpq+esfVCcJJSWuPMLbqQX334kEhj+HeWUiZ/FhFbpui+1oiwiXy3CO5CoDtAGb
UEdK7ZeA4lUXtP0zJx6NBHEG3rFTtJOgHb4bmaaOTzzVp3niU0PVPMeSfkKda+AnRFGsB38X7ySK
m8hm8Bz0lyLrjNHKeSLL9vI5CcTk2GJDfsL5t5/OSd+jygu+z8b3TkGcZ4zLDTc4XGWmrC78FDON
NQyoIXpnZGLRHKLsxsSAGFZR8hlWcHEDJlTJvsUPM3Bbtx3tVP7ViAjSH7FeleUpmRYzHX0GsgDC
fgZsX0ON+/D0SV3kNVoCnTF7cozj7m0YnEtDXXn/VECSFYBdP0T/utPjCb0C/y6wjAjWOqEQxL58
IpT2yI24Ksz5Wjbfzhw5A2XooHHx2NHDNJSAq9NXBEOgsbKNYKSrNulFBaxhJIz+9sYaP/rKclLg
Wfg3VJVvRMx1PMWpGKKjbyQj0r+mJEPcPB/IFj/6onipm4yVRYJF1NuRhJe7vuIKBLzHkHXOXDzf
r+1kn6tpcnCY/V42MSB8TehGAA62IrMUpirutUPEQsH+TvJgTFHzeVYV73ykV35rkCkyo4mcNsAf
aMdjfzE6SzHTZJxORyAZCmdyCfp3LeL9ju4+ufVxCLvY6AozPmnP68CZDo3uMEDR6/mj60gLy8Zl
SR7LOrWKoyOtdG9/sPL3BxGllWdWsRJV66j5xjQ7ohrx7S8nJtWMsCE3/nY8v3Ag+kr6ZKr8kluq
eBJcSOky/cbdug6W1mXQl4fbEVcf2GRRj/gRXtZeHT+ZSV+1bQlVC7LHXCnr29b3OHHSvtXnaTr9
ODAKSY2b2/ccZtzwHw/1sW6gtnYr9GFE+c9AMj3xOYPRNa0jkrfiTKM38fC4T0uzsmW7p5zdhkrU
ZqE3v3q7gg5VhvZEIimMmZ5gDYVPDOCzjiWk15C/v3mO81SXaeAEjZaDwZCfzUjgmQg9q9D+XRna
LIG2WVDlHDAKiROuw+ilXtUq9fvfB5ZFsVp/c8+CqpQnc5x/P7iLtNr4sXrDclLyS1FxKJ9Tu6BI
8e32W/UNa7BVaduL6rrWL+JbYL81l6BlFs4+/eWdFc6TqAaGHJjHSp8lsT8DobWkjBSjx+5lGZ2B
vn1PasAdVrKJRbnO/7eyMtB+a8q6wjEcbeh7E5NzZpubIlLTlHahrViQLJtKsPzYGJ7xdo27vdly
Dl11O7Xr+TG8ilyD52QV1dJpyz7kLLMLAxutSQkdSojIQk2gmhK3upO+OlZfIZhmMGLuTy69WaNh
HzT8sGQf9kedC+xQ28/BDE9fv+aDiTV20Gobd1QnTTy0yuHE9/cNTpTNnNpEiKeW7tt4npL/+io1
dgLI2HFwYZw4pDjGBI9kjpvg7YYPne6gYV2VZk5r0thAjPT/7bdMvpjQSaj7gfl4tsKCPZRrQxGi
2H+eNfKF22qgAHsz99ZzFR8XvluqXbzZ86NY0d0P+Sh9fm2xO9os/boQU+mrdN/2vw8LPFjTjbHV
rJF0PrzOwdr+h6ALDRfzaXmRHCufEqvzp0EnxcZVKZ5nnbOLy2Qsi1y3x09/MrAvHOnArCAqvaeX
sU3IXsIQulQJZFMrUx9+QAYnn7LDaeZ9usxbILOZe9xsXeKPMMlXAdjvNpZsdX24pH0vV5oNnNGO
OGYj2OA8brLRFbIewOAW6A9lqp44wrb3cwqz+WljCyiIemW0ElE0hAvolqH10ytw639IdfxPQ2BU
7dOmbxfCu6fXvwgVe72cbg0gL8MCpZ4oE+3lfA1rRZDo1cj88IRs2oPZilmqsejjADcGMDiqKfRL
fcM6W6bIMiSSPEMX0LlcBCvhRCNzr1ZnkcNfYXOWC5rCThw9eQmxhzqmlFA76X0vfjxyERpIGB2s
Kbj8RwzCamh0k9BRN4fyteSrMgRhZ0cOHI8a8D7bJq5fdvTn/OFqsIqlBH+54gfzVZAGnTwYy1ff
/Fh+nBrvcCN3S/WC9foRocYUYmo73wBULJ0bxecoO/BvxjEDA4+Jn09is8pbclZWEMeDcVg+VJM8
AJ89TSMXKk+mhCbVF7BEKOGvOax2ViicSlVASTonGhAf7LubTxfqw6g/AOlGAl2ga/vl6ZALoI9Q
zTQpUrv9ncxZcftsLZ5jTQOWs5DtKCUnB08UOph90XltaD/t/TqFI3q9QdHmTGfXtPwIvQauRyAR
13tlcylu1kFlaewKIoUTf/qKfg8SsuEKnLcm+KOz6+sJ5usW4Oqde79UycMJPLUk/GCUBOZq0Sjh
Qz8msQPJBpo0BUPs6ooP9zBeOaITGhJtgNNYGo2Th/C35171LpeU9Yh7vkQy56ISEJc7UCyKrViQ
Z01rL20TkE6hTaCwvPjZDyNuYsISAkbmHgxbai0ZkE24/xLMeqW2VM64OtTPFF6hWXCK3gNxDZUT
bh0bhwiamt71oWmlmUgDKZ7H++h3uiN4JFkihELXvooSRGaDXbt15a40bZk4czIoS3/IiODp84YA
QXjMjzkvmFWj1aT6kvEOsaOgbcy8NaZfZclynvyxPDsNDlVBaLToknFXHAxN6hdXiZgYUNpLBy49
ylGcGj6CjwMGGuqS0cSYGQP9ex79EDGeDBcvie2+IimtCKy3qoEPiX2Mqv4BtpBrXMgQiN+dfdQ8
biej6rF4n4X+unqWqbsI2oxHgXaTq6zEGT4a+cypKBEndt1ZERRxCWCQhyl0RpVfIJE5v7muylUe
yTXx1gsNEZpaE4gNvVDbr0yICJ+XPNi1QWxTStX9xJlqvTahqwRU1usjXK4ePQdg/4x23RbHu6Rd
ED2+f7U1uTUFQvwVTnJ7tU6JqDxykVdAfqzSSNJ+4+pHLwWpH1HaON3y5Za93/XDgqjDeFijyGGK
KPqT4XhRKI1agLAh+oYNYXZAMXgaCPmajDk9yXlbfilCalo0FEQuTUrPKRP3ZWJsHtz7EVVzSDLb
5kW4h7udRwtgaURrKIITXea4lT/qCm1qvPOsG0vTLvDITTubI5yJm08vYnYsowEvcV0iSipZAIma
b2aHzRqTI3okG5D9TUBbR1wtKCEEzeAUZOpWfhHWfoe40kK5aQivrPr89meycBxIP3OIp9Ctbove
T/uk72JxC93ppze/9CG6w6/hnSHFWBBovzZlkyK5JWi9b5zZ5am3U3hpIKrBrG4hmau+ONpSyQWL
XXFYS4fQ6zdlDhBwKHsBMoayVTZaHYMITZeU33DD208zW90aB0kMVbAB/TvGHh6E4a6awhd2YaB2
VUw5EDSDDlmNGeN/tiZwnYjFQDz7YzW9YaHkDBxq6Miyq7OYbYmHarJryPls9Fg1s+JB4PHB77rw
MKGYRRBJKkiTuTnEfQVFLuoWbUFzAJ+JGGnxHJSfhcRI9Ht9WqnpR9uGOFWghfqIF3dXQRHu6BId
miqskdR5xzq6Nu2CaDSeAo9Sl6NcB1MFO5iAyoiXPwqbLYzLycRvPsWkb/yisYftAuVgIlRXRrIR
WDsCtWIjcDKhl88cHpLaj75kIRKVCLlLDMqrA+ilubXla8Kfg6EIOTMCqR1jg3pKr4Gav/flDzDN
c6dkk4jhiPmeWjCXWsks0zNTuhryuCTjtuRagaXjs2nkMBrsETz0e+YGPoMPlj/DjGjCpRI1r41g
ZXDat2RWvvEZ8zj3NZbj+TH4OOOGWYSNF3HfI/JMUbtmjRjMJ30uA8bkTtdE6AUuw+lMknX/hvKF
r0eWLu+omYOz6YNVbZ8frK11Qo6PZoN7rfEos1HUaPMBNXpUOBXjgbRN2UyXQSbq+VU2YGk6CBEC
4qqR0kjrjDzncf+05tod5m4xuhM/Uf4ssEOZvv6J87lryTrrfogfdzlLv+JaTGwPP2Z7Cs0uwFxA
PKY//Va3DlKCvLcDP1LyEDM1RO8g4rRzTdx+8Ha/NcKsCV6pC6AjTEu2J5MkrVgDPGd5+FqFA9mG
+wLJfLELInr8TMyLyNyf5yw+ZeMZIk60k++ZWCG19z3lLNgRZQ83YOhQ5rHfjWxt9lh1uHwxknhv
9ZY2pJ8e62G3p5nZw15i9a+pDJfBqzF14qV2fFYMMIZ79vxFzNfQDYYNSHCPxxrR7Opm5XTMjFR/
9hzY5baXMhMe+BO5OswBRVgvAqhTV4cNQmJWI7zFklCMG8exdDnd3MX6LOdp8qs8RY9eAl0sLskA
NuMtisMZzOqtabTX/622GICdnl5jbSzqMruAH32OoERjNweh9zsslIzy+aovIfLLUKpEWwk0D1fd
8lTfpWZ18gKKrN9WDGtqC2eZraRCzDxv9fvz6vogRN22If8KzaqrgWjiEGdFVdm+Joce4XVcbPm4
KjYVzhhhdQn9HjQSo+6wMss4DBOPuxuICcLdF6+GiyBrt2X0di2ZMPXGfkJVwHH3rx4M4Igmf+yS
NpacuiRmTt7v0npKguA/H1/u86D860JnjLRx/mu/RI2KgN9w2Ic3PQKlYpT8QHeGrsAbj+oc3KDs
mYrTCPo263EPRlwvaUWHcux/W4fk9qyjqzK/z+/Dt7EvSGkZiAj9in3LN+dAPseRd1cCMU2TNdzv
jm4Xk5owa/ZKs4Oe4v1KFxzogPsMvHDKKP2E/+dy6Mi3rjRp0uSGhVkkcTc20HRF7ncgTe9ylSzp
y3taIzWUuvbhbx1ysFpt/Rgl0Srp7stq8GchlZ2ZVgYCE9XSBAJ8ja6tx4h7Q75X0qqweBnisVHt
In4cNSk5C8abvqxD5cvxTAV+cWa5dn1T2lzEjnZVIAIs5wi87J7HLq47fqM9QtKZfWwZnmX6bjfy
ObtiJuiFL8ooLAN1J25bXgfIPopNcSu1pdTZpQ7ZDucU7maA7VGHqArhQ4KC9n2ri7E4iBjTldPl
62Q7qfCYQjVRQjXNtloYq5J4mYztY3a4jWOdjHLWbO//B6FIgnsJOMPLc2jweiXOo+RiK4DukouD
GUFymxOmIo7am439pYYie+yp4UYpSdFpxBE9eLeqHu5gXUA3755FZfjKpftr/fAAgWMziJN1gtPf
48QtQ9EqduM5jlmgBctponOQvoEX19zFx9sXacQyzW+dA2SF+E0aXgg3dYnLaiKi7BW9MJoxMCcR
kC9Xq2FgCfMEbSWUqxGk8h7oYz84ggEcDbR//t9DmGbtiHIOQrP1kx6uGoE5Fx5d79ro+jj/YvA0
9obcuqQ21igvmm+gWmolj0PyLAJRr3HwPog83vecHq2k4MXiR8etCnPF+s36XeDkZ8fKtG6LZhm9
kUkLNu9inENwVe60uXLyMUQF9C81CI2SCT+iB+ThktHAQDaMJdmTL+nz/UY9ZUVP+KduIFPbGEzI
AIFcJdA7BMdGQKC2oqXavmEgZUN/YDkFmrIvDi8zAvx/IXt4s9nrssS6rDTxiioC+emScOVUT1PF
Cnpfs9fjT9xZIIpj2mmkMThtB9r4N5UJWvnW6Y44N4290leMmXk8PllVByjhnb1qC1w6JLL4wsGv
J3WeXGrHMYSve0iAGfTOZeYd5R2Ty0ZbWXl2AND0Ym3/hTW06oNntD8zzmvTBoXsKU0zVSDR2cFy
5oI1j+jpwPAYjl7NrF+hinNVt/1x3oDnLPEP49CKCEgrht16fitFbO8FoBHuirM84XyPvLynbkpa
7fuSdLlOQ7wZgCY83xRCasnN2kQZwEVf4V95Mk8X/VgWUtjf+Q/bTEkUHK8DHuk88lP6oQQ1laYH
v9OZau7Av2Gd7R3aWIPPHLGD0ZfEGruIhJ5VoKW9YIMvKhHWZFAvzLLcxGnQAuV+OQ88vekSeOBh
pk5N5Nr3fsK1xsSPsMeLWgGinQdJBoLqsNXKyYhloEa1S4iLjvg6//aRMK2h8s/s8+ZAo9ltmfN4
BFWy8Vx3w2MA8lMjS5Nw/0kna7u53pgDdx+3eRE0e1cWkHd9KIrSnkjFqEpvXfWSQCIPEWkWeDEc
37MQvw932WrBI7wpCK1S3VOviv+/d2ujEJDXtpcdg3UaHYP7OI8woPCdDUgslwmNioYle/pz/07/
b4YYv4qUQv76K5EzFyeq0GD3ASHwksMluFokIfIRRj+VMLclD1bTUtlF6X26v8q+BS9EsozG9XAn
tcbF66voZwIHc87216oTbt/Aq+Cx9xVAnTxOQkj19yiGEYy9EI+omUNGVNzHUqVXjGOMafUVwW2V
VuK7bLIQm190OoHonknHX3tbA0tawrzjnDxemCqw9PK4dCvHjrKACjHJvJDqs9EbTNAl76julAFF
R6SKxf1lqi9S6MpXaNaTCYALnhUJGU0+gIJUPVcpyWoIqABLwyMgJQgcX6e1sCNeqLxRa8gaLwZ8
KEeVTdn6ZJkou8AzofJb955CuzGp9ZQmjtxsrb0/+hKZCZj34+cTNccOae5L/fx/QEDMHsvlVWf6
H6AgzQVtVJfs9IHvASRQGH86pWdsiUlzpJRUCIWszZHIZyT5+N29dOlm5Dp+h0lJ6g6DbjWOQ/dE
hqX+fKc6GaAAFaT03lbxwo8L/OBfZt/p6HWUeeR5JvBgjj7kFPvfZzA4CxDmIemF3823tEA6j2eM
gx/aMg2JBNfCkW9Ao3nFs5UXbhVRM1Lfe/yPGRkHizlCNaJrt/vpmJ3t4BFaVr8pSh53DkKdqFWs
ryreeDUiMZJqYS4ZvoFhzKqsJGaZ3y31vRsxwo0Uc5r/vmyIgXm6wAd8IdB4REjd3Pxm13509FMS
sXFcMsdt8ACDKdqjsgknvbCX5hE/oAkFX0VrJqIuHhj5YgShFJvpK6HCpo/0CAwY+ajCiPnkN+51
a+nF1ri8pDyqfuq4mfNsYS0/0tAcX/201Zou9lSf10xPcWJvxp9AeQqvXpWceECXboMByLNVpl2N
ImZqH7gBDwHVUVQ+BFNHUm6WEOfnl8zvnXMlvYJ7d+TvhIHV95d5iUzMeqqUsWyesnbRfgWtGWaG
xWkYbZbtgOGzvmZkDv0ux5uEaQOUMfAly5AaQcWF1Cjw+gx83y/ADQbjOvVDv/S1wYzz5sPXx29f
L8oaakbAqHAdY/wW7MO1R8R4YfBiJl/rlhCbvf/OC2hzAhbt+rHQI2M3fwqzGwgG1GGZwljkxU06
M1+xd0Gr9IvdW8UOsEXgO3GWibFTzViMnX/XEBlJuAYshRJGSgyAT+e0DYDFikZSMY4c4qLiwSbr
+d6hGsjj4tGVyUlsl+uPsg3ViWT0U+WUe91oMdhKxHSzkbWSs6ChwDndU7AMiP2Lnz58aMsl1Yvm
XCcQgnYUMn5YSXwN4SXZYp1Yp64RoV4/WArVpBnPsvO0NoFhBppf4CCmtrokTkTQfTQe9AjepGbo
q1BLHeSt1AEbw0jNESVBk7gmarXRF04lnxMycHrdEieWYR/KTxg9iH0JXtEPxTugQM3XA/jVOnWv
U98jVtLP67zq0uQqielzZZZMy0y12JU0vKLruyEsw1aaWLnct0JUQu7CQHXJkZny4034uPHvSfnu
1ZqNvZcZ4WohIghmd5cqbFEkW8gOAoDIDD3jw8nTZHsMQrsbBK0CrmJdHfFXP29l1QJijoOODNVp
n/Xkf1cyewVjsh5im94YOwUJCg6bOZGklRldh8xTwlhPz81+lkJU42IEhUZe3UZuIeXQznO9uTu5
I1S8awanWpfgIQgyi6ZFXSr9ez/Ti47f8eYmbyyWsR9RVGiach1ulLJ6P2d/JNndLBV45wkQ0q5a
G9y/dsrDlunGohFk5Qsk3AfmuZrKrwAeh89r/QjQoqFS2D0kEtRADO/EsoHii0YXbNLjWuKHkPzO
bsCsgrAt4kVeeJvaecmypa/+ZyDnxlRkQXoznj6yjkMRKpjDx1DdBOhaeto12YVah2RUq68omGxh
+LE2OUdMbPR2G4xzK7/WktRm+zUTh1a4bQpT9SyctQ0ARVP4lFjxDWzaNkJ1TVYmzCbhczZ5I4NC
q69q35j5Ko9WJiu4GW1/9Fj4o9g1EfpYIaluAIS4bSWOPfx+cmkgWu2+J8hhWCUPMS+PQ0o0A4y9
O0GbqzmXa2ZBxHnXOM7fKtmkViDGQKybDalmqqxOBMt0qtPTKxg7hEZd17KG5Cvp5xSotSXT3mJM
JhdJ1tiF9IGsjzx7hM6xz7C1jV5lw92qg9+t9gAi34BEFQ4Tt/3rUhSj+RErKe3Nmhiw9g3zOhph
DOdgQZ9zSY2Jh5ixjjItULNbVq5VZlnKYwp/5bU4HLDNSuuHqTKakrvhmbvEE23OE6j7v8JEni11
/1smM9pzJck2Le5P8JKvV85geVlDP75gXl/arAmDervYslYl4PpmiXzgZYVkqFVU9vflJ6Xeac9Y
l9i5FHmTVv2jilIpRw8TVC82pMhSyfhVlVTmS6KQwtOV3gSbKEBLD+UpLlBsn766T3UMjOED3wva
P5cICAFxrj0xZ1RTPwcwmtErVMv1dZ9bc+ykT4EJPnw9a30UEsP81fEee8cPi/2xGHgzhTuLbxZK
4nClg19O+BHN6brrNDWAy7J4xUOBvLrN6GpzLVtp0OWbk/nyvO9IldJ8MHLhRoV6tPj3rVM8HPII
NF9bm1jnYDAIHo8swLefdmes8PvF4BQ6sgSRO5ba7rsEdgDfcSrTV4NF0rHLX+1k/lhFIRGcOFeo
S6R2m3Tp7AEANkW9PgkXT6vQLNRRZ7UmAiJUnsF113W+gQ+ORaLO/tYOOVeztvzGKRHZO9lJtmkX
yx3vzcsVghEc7C0Am1wuqGApK/I6RoxniKKWUFil5G9Ph3zTWBTnNDzbFIV4SSNS3GMUM3VWU9Od
wvIzWB5DyUiWk9/lxsExZyH9y4wOlWV6QKiMCISVCCoDwjPMjHCtiUWRJZ8bXB64roE/3WG9/PCz
TgfUvCI2oAppzt95Tj1dDh2JXTO/4cWgYd+jLvDolkDN85L8vefJ1nqXezamYyixccm/fcEBJwe7
YSGUEsPmsZHAzj/mXJNitjysUjM7YlLP8vBr7YKpKA3gKbMcoF4mWV9LmZIvoWhRpK0xuImf3rdq
iWtG87sA8gOCVugljzpuWa5NzjxYMSyJUV2UOgnAT1Bd+3zDxXxtEHag0oRfsTvWbIMAznFZrXKR
f+C1zW3oc1zVz1gxabg1a1+O8R9m6lDMuBVzrdng2jwryARtBeGKvIRi+DmB/JcVOrEv3A3uUbYW
wpPdWS2+aTprz5rCZRHmhf5x5uFloE1SUra7qQYYcw0X1r8fTWJl2R2uKdF+rphhzxTpRM2utlvp
LUs3ZaWWv6DW9n48kDuiKqTY56SGO0v3G2l1+8y5o+Qn3IA/2ve0BwWeDzvNaLHvr0wcsMLNfvdQ
tfTPa7mdQxYKSbnD9Tlz3Quz2Mi+r6R3qo23V9VF1g/aOAH34IScuI3+pJm28jqcXOZsnC/ubc5w
9ftWwKiCZnInDtHqEZnVXoPCZrVYWEzZ7+jTOcYGVYMj7CK4RW0vNpsMajD3KIBDRuLL0hzVsgAy
ZPKfm6Xndvk9IDmSN6NKWYETivHruPhLNNZtWWFw6xdrDL9hpDyP/igL3L9UdkA/oJjqStjXQsmB
OHGolH6/UeJQn/lj1yTkDULmM9BzmsG0yo+HbgNAMkOlE8c63nca55djRjyfkk9zUY83SwUQqcLm
60/8jLA0zPP53wUd5eYaYAZzGNbiANkj9/nk+cGsC/NH5Fawg/BrTm1CDgyBqOjS8sI7HUznOFla
+32tfpBs7f/Fg9ZPkUiWYYmAz2vUG7TpoyVQ/Z1GpEgM+J2nn/RSDK6WnpIow0aPQx86CADBKTJ/
l6n1tcUCNMrp7v/UXSrzTz9AbkVdM4fPXt0fKxZ0/QiAQEyf+w4podWRV2faH1n+02asGufR3Qci
y5le0mFc2XMdjbsblQjHthSIOD8nMVAZZXhorqYrcDuBl0BLN2KlH4YmF2PMaz10Y6+UlXBvmsKb
AgQ0jZ4WlnTxaDetT/LvLD3EOoo/uuBql8ToLeRSTGIyc+eAlsjcXNXs6Siz6iEUNnty6H7/rlVI
/VlJaR/kE3Jc+LEB2RlAv1ll5u4bs9Cm67xVAzxG0V09kDf9R1f0pNx3DtIAa3Fd6NPV6NbBRsbl
buzbAJcVJ1h3noKGYgbIup9egEbyWCznX7MGBrvZfBFcPXX+p5wFpUwINvb0H1x8cMPb09iZIcC2
85C9LIyFQ0zvmxFnSvDpOZnRqT5TVBWltYS4UwEgsw0Tn0RC39F1mpc2VYwiX8htQ+1Kq1wUSemX
ENq2fQPBqmud28fo+xD37jZbkI/cbfx72NgtfQjYJHl1T4dk9idYeD82IKVpK2sTE8G3XQRmFF47
8qDuN84hBOdxZovr+vnH7Ug/D4q1OnWpkozJ/aTupOtm33NTIeX60AbOAbIQrGCdmZq385CgqoWJ
YzZ95DH6k8AkDGqSO/GimRFyF6SG/IieJ25+BbmSQdX8emHrLtxU8cuYZkM53OsLZXLowGMz1oAd
EvKDvPDh4i4syw+LE0a+i5ZBJD1+qNXS05lZw6Cqnc0TChwyVtNzj/3DibyQPgOghbcLAn5s2p9c
4xoTu0BSXwP51VrN1YdRGMi7GdS6X9azHW1/0fxpx1xntTUM3Xisk1t1E0uA2K4M6B7LrbZVm6GD
yWgYyPSzckU4RxnW+B7sCdzUsIIV8EDsT2pJ6vdawSQs+izsrVIWXsqSZsq82BEyQUIec1was2Sk
2iepMiSToXreAVsmnqVdWCQuwyw1ohzTBbHmev5etcANwCN42OCrc6O//XHdIN3h32AJd4TTpB/t
9ihrczNYWfR4jm5fcxNNYRoVvxFpGugdN/Xj7A313roIBYzCp32x0utILNJ2Kh0DUg1cbaJENNwi
1pDdI0+InwuIquuke4fXyemsj3VMcCHuB5ZMQMHQMHn3ofptt68EVre8RkRuQ88UonUXORX3DMcM
anJT3QphyKVRX5Q/ySJ6laBLxFAD0wMpc4lMJgPDHQPfHOnxdWo8kVbUSJ0E2wPPF5lpm3jI4VQ8
prOhbLeEnw3f4rBsoezMQa1S3Qh3ldyzvIJ9dEZkqlsFeAs5D3M10UUSAW73LIRP+lT6hsb5QM3q
8JhpUMd7MqINuS24TS4eInlEv525aKRh0R/pH2U+geAtlShM06nVcZjyQ6HwdXvHNgN23zuSS2h2
DIVjY1u9QxlWwL/jzcA31bPeDF32kDw+RJYQWe8DKkXHQYGAAjbdr/25U7EXPMfMUko98/K87yga
ie+mlcBYVUJkHeHIS7ZVwuWMZylKddERl3AmNghkrhZc9zf+h2vm0XhTx35KQCg9bYplT3ZyKRgZ
CGisGmBfu7Ba1tQy4qKMq6UdyakyL31cSPkdiun1F0jMCCtOsiHh9ogAx6E/K7Ei/M0768OwO9eW
FSj07N5rtMrRGH4Stz+KevD1VTAcJN4zT1CTGm9MvXKZV6+YZ75D3UZBZ9SOUTGBc8dC4lVq1A/y
ARfrm9T406T5BgGkGUa1sMWNqWCLBvg/BksrSFeNUZ7QV0Fd+rc57V2r1eCckXHQNOFEC22JRvtt
F2zZEAhFdcPaIjMT108KkhMDo2j9tK2IDa3jyU+yk+uHHFzHj9Rldw3/9It83AB/nLhKRWEMLGNy
7vhYHsYPrR992nKaL9XRahLLVClnsccT0O/rQtXYX+AzBc11U43ducS83klxprDF6ea1ML2Sl8pU
//2Fjyr9rerGR/2ThiCadxrF17al3PWuXP/un9aq93WrI0G/K6uMVC6xWGqMfcCnhHdSDDpaxkMz
lAXxC0p66u22/LxEMDoQNTKKY8v/o/4tqS/k00HBzxfX5mJDeXLyMY+rCkzZc7DRh1CtAbmHOKKO
Rh7yWetW6owP7FTO1IevdDBJi64TYJjyRlmudN5eiIkdnx+5nE/Ypkbe67sxH9z7loJPSPzG1VhE
CWkdV60OCCj3CHn+T0tajv90ql1LfEZby7mlAFfCJnvvMb4L7/lUkT6KgBaMBHEAkCMg71ildvAa
qlYk/FqkdnzZxRA6b5qUBc8QJ5R6NDIobhcJtEod02qd5r8t4gMNYifXTrIF6Qob1giSVJH/N+HB
kIesMK3tBnVvXXY2xk5GOio0QuxCfOqQyI5TXHpdwvi5rUEgYkuK8pNnoqWE5f1ud9ysPPn6DQcn
+crhwoXsTuu/0m226tTdYQCXAlpe66kYXsAw4ZUTfkP0PKHoCDTTEOo/VoDs2l1T5rBe9lPKBbSF
vIPTa7mbhetVF91L34J9L8vJCXPxm0d/KG7qRBbcOkgpmmelpZmM4AkSPRbt/XYCCyyKCaj2eMYN
AmEGeJxJe6+APzP9zUSDwftmfyRalDC9Zjat14Nhp+UFVvXoOZ666eqkJKoBk8A1qNndXFSyVHC6
9OoM5wrLV+9TKV5We4WKCXXFTEI/9X6guPHWKPeRkKHBXLPrLQBzS+/0F0zASgZxaQHcwD+F8yX/
BZwOlH/5K4l2jn64WKcqG6bvZsyBI9hzou+kTzFgVpLBZlFQDqIX478LkY5+j3IcjnMKX4kLr8Bt
tKwl40FTmJQe8Yudkas1mGUGqpE0n8BrYO4UkJ093wuSxSOlBCywnM+hmUM0oGRTQUWfreO0nSS6
mj/yi985fp2xlLWleeiiEnU5j2x3VqnwXhNSV3tttP3PYmktv/vws/fG7q40zKoAuhIF8x9OI0M5
nlaKZbxkRxoqi0rPDbq3kBPgghlS7u4MMpDD1Jtzvrxd0qrFX8mF+V33kpj2SLJiVXKazCO9W8zT
Y80020XgbGM6+xHAAq8qtDmsh4faOUvt3paAyQq5CbDB7ds+SRwCUf049SQlSQayl183qFg2hiFL
Q3lWBD16ornSfO38n/wKLF643EcE9CoRJ8ixUY8sYiCzskJo6SfglstN02H7fFFfH3HOOPZeohs6
ySupFxWVPC2bSxnry8Ggo+7TbAAu0X3uT4/zC/q0wIMN2pl1jiwwIR+a6NWOF3ghG3Bx8mzpSVGl
jab4O/4wLVhjuOzK5tfUN1z/U7eJD9bxsdEArBZCXiOBtEv5YelqOZ2udaqTItbHUQ2gUiIJeyZF
zMqBrlcTfgs4ziiMJPdq878koruOjYYrv3e1mtAJReRbr8IfkrlBO7O9adhsxEhiQs7OzAdrlMAT
UuyrueNQQ+jwVarmLZ4AfsynN+p0T4ezitxzOz6gJUsspbzAnnfSv+M34yCFxm/946CRtiMNdv5/
G/qh++jcjTuCBgsul8sSo2Jcf/cRMVJCtv/aMbUdtA0pvjsCOIa4EwMC2uBHgnvpWi0NtB8EAgPy
nyyF9Vqby3yVon+7DoH9vpw7SJqM7hiMr7xruwqVDjHQsTVLrNjJ9DAV+l/mFogi99UhHPt3NILu
RCSZublJAKCDYycJdluRT6p8MS9hSgrOaWoLTzOz48meQB5RPQ1gdSnWPQ3yKnW66cZ4UNN6496f
QmPIQiRjenSsrWj+x6WjdZyv/KgJ2SMOB4vgAKsc6NFvx8Wa3NPzpUw3it5QyVfyi2cWaEKaOA0/
zGA5geaJ8HA06q9GUi0lYy6XkAyflF7lsjnA7VyCwZtaToYvrApWGeNV4jw6sUfQpibfuLPKw2UT
Al0jFGx4hVWvUSOdMQ57ThjQgnYhdWCnqMHBgsjRyhPONQELYbvn8NXVygi2HMaNqAoFz4TIipT8
xcgBInEviEWWQS8a0/D3Yr0tQW9gk1zGQViZjv4CoSJsFztHohcY2fy0/BQlysrnq87dEG3Hf/EC
VLYlG64QCaWKGBUXhQt/kIULycDUePWLh+L09bnpphmKYBKxsVUfQRALPtdbKydzFXt8CW05Bask
n4hbzCK+uOJ6cwBl3zuagipq9+dclTTYBliaN2eW8gLgnmwLe0jOSrrCID49uNmLKHzPQGGPB/We
du4Ih/5kOATVM0RIkGO0CrMy7DNwHqKpOoM1qHoxPBR/U7/tDvIR7DACwcqCMhP9jAtXh87GlXqb
qmUsA/2ZwhvMdkgR2Y1XYV8b06vm3rnJDtI8u2/bsDTOiD7N/+/eLTC11NsKPACyqkchYNpxTRHs
F+Bsojx+ZfD+xABaotox/4Zy41T9NC0xF/+GVPiRF0cXjdVpPpXLvRjPKfDzZ4ttRMV2dfY7qBrM
p5h0m7LScJa5Gf0ayyxHnxNygcogbDT7Fzng8eH8don9MDK4V2lhBwRBLZn4hBcHApx4+J+zwG+o
KqJvB1zdkVIqw+xSDLOk613/u/iwJPmyafn4qdKwzl+WOEuI2BnxSqN0E3GN8Boaj7o/vVMb+d1w
Bhi3WfGVq/ci22a2tj8BKyWahfkZBaUsuVPW1aXdG/fbOzBhXUn9QaIsWs6xSK4ANw1Wae7qXCGo
hoRvQ9rZlOApm0oheOE8G8HDsRwcWPTtdjrugREnO9UiKzlPzAGs5B8SWXz+KEpRHIvuBLw16JaB
ss0hGIVwAj9CWk1bTSE/QwAheiFkE0Ye/ykp3cZB82jxfEqjRSlaTefR0S2IY1/gDdgC0tWoF2qS
iBz27sH5AbGuHYDDvw6+tll7J9NvnEkUlLXs3jiJN30j232WcDy6x0fyBkcjE4nTn0PbdrR9dMjM
rqzVsphdVq9Dr/892UDLBPeZXonRJj6j/h8TftCL73KlJx2y+SIH1RFxGpWFcgyKiG9M1knLG/Ac
waFfPOtjrMUPLzU4mYb2/R2tlGHZ8q8SfEh7Zrc+VYnUnsfn9IKO7yPyXQpjwozyGoX9WQ6h78Ig
T/u84hY8ngOGtMbvLqF6FoyulO3ZuOJKqGEJXnYOP3TkLOIro0kA2XERHwOdxANoBhURDuW0JVBc
nfxi+oJ56h9O/qFhjmWC7gaAunQA1Jqrh9Ndt5gRQk0iotdWDTsXNwu0aFAHCspKodEcf//LhjGU
2LhEY081Y8+HhRB2lb54BCtDtllKew5n1ZB8tw/7H7X19R78ktjo7tTjHt4ViHz00v5Pnx/Bn/O0
rYamYY1Ozvtc6ULdK3Zdqb9mVQL43xB6VEe63mlbiJufuGWw8weKeG28nSNjaecarF6DYGM1m3bf
aJa5C5s44SI20faT5ML+wX2Dbdn8MJW27//sEg6Q2ANWz91+rSo7Pa0EfaAOgnllsc/a1Dp30lJC
2vbKtAsJY9Dhtlyacu1tAb58iJKNzFj5dN0pI09ozFcIBPzorqX/GyQIAUSWrzv4DcRIcQ8c4Icn
+MgKzJ23xjI2YPtcc+vXFfxvlm6l619JCGAYfVbp0yVml9X8EJODfDLlV8UKtBoynHSkuawsHfAH
UgwvXFVKdI4eTGKg+nGvQKF8sg9ZH8EpdVvWokaUDJcIRiSI7bUf79BBWDxGQT09QmP0h6vk1sUC
U65fOxw5ojMEfIOlHT9A3MhnwO6JIBfhlHISEO3432ngfaX95v1ZZcmjaA4ILo3rA7JApIKTeANz
Fl+fLDsvXLFu078ppUpIglVIFPvI8UkevuwtUpyVkVEMr6aJbkOgaqYgDaiJHD/LMOEB0UxTPxc5
cvN76/x10rgj5Tb9OF/t9Oz0vZ5t7iZ2Qa3ufZR557NUycaMNOHCO5WR3lvPaRvJ9A177osTKdSZ
r6HiExubCe4rV9iSTOTbd+WeljXubUILR4SlPRFNLZT6ZWFrPpk342KSK3RnO3+8JM3g9/mdKDaX
6u1vSXrY+eTGOhwLI3Ae1Hg3/7Ga2zPOa1dTbejQUNgQ4EyTL1+/1sYJI0DezSoDdmyrZnaYcH2/
yrjEY8NLhumCZLyBJrv3gE+2EfNwQwG1+MbPO7y75Ti/TeasaCw/HDEsvyDclNED6mdjhnigTEiT
XGzCSHRsFhYOkURKag5j6pMs85bAr+nNMrliZy/bSrAhszn1iSyLUr56601/lM+/yEQr+Z4Tng+j
hu2W6lBFA4R2ffnlOirOj5fwydbtDStWrKL2Pd5vvjYw6+20iRvhl/cqvQe4WxGSBXRIxyCiAA0E
S+FUY4fbR3nxW/NFy06qmOh8X80Ep5Y1+GJ6DcSoGZeEwvKuIZKdK1pZRzjDsvzyUT7Gh/s4skXG
WMdadWQ3i54vA9y364d07gcEca3Pg2fMHww2Wq3INybDKFZ+O/zSf9zqt+D00r/inGzvl4E+jlHo
Q7+1+YeeM7wDDzneL5V2AHqdRPbrDwOPzUqgXGbg+2UCA3g/uE9ELyx5L9u1PFFRC/HnLHjyskUn
ucdEzJUbzlbx+Rk6yCRFwZu5L0NYALbAxuDacHgTk659C77137uDBAP/dpAXQkbQ7GF6kNPsoClj
He48bGbCdKY6rnAGqfet9dcuLXk6f4tjdo1yp+3eTDQmNjbW/Ze8oiAsq3MuzKvlyaeLph9pOej/
NhQwhrdczvvYkTvVxT9oyT0Zc0q6AV43/kKvPk6x25n3mDAR3dRX5KteMqRyEaW5VvRhln23Pek0
ZWet0Op1t23C/vrTetj3QzbFx22/qEWu+9CCwveiuNX8SxXwYEd4vvrxqpFEbOygo/M8cQsvsgMm
ZE3Qqqs4lW79743jFuhBZFkHx7ebhyjyDbxyfauoPwLODiMnhunsTpk+rjHxcpT7DeZxXjnhc1gf
ebOytvGS0CTbsEC6zEdoMW909+wOCVfJ4Rx9p5rue7jISjnP6lHLsJiQnGKWkNd1qD3gPxCHuleH
JpgvEM04lGTNpcqsH9r7WEYgHAMfDS+JdzKe2h9ChU/dDUSOOSfj9KsUKPkzPrGHs8gT+LsbY/5v
IvKC/LjlvImrH88kjmeB02LcB7rB45JEuBmUvIrGhIHepAdHTOw1Yq9r4+76ondpuAnnxnihfEOJ
OGKsE8Q2iwiq+2ndpjr+7m+kO3PYE6odMm1fszSO4HqBdgonmWLmacpv7xjZ9YG572ZdjIuHx7OZ
en2J0e/cH6E+T9IevP5INmBfSvkxatzxM70MCFB7UORLC1zHDZyOK/wHE3fEOCuAtJRiOAvyiDpk
/m0LeuB3uLUg2NB0vcQNhNX1+wMXwQ/4ABkeDA5Nm0lyHEGl0zWkEhx8kRpNmjqJm5iMiDtYZFAJ
2hhZKTW8qOaruwohcl9JoEoc/20MteQ0aZrej+FzD5TdkjyHGpN+ZNqWLKNOPZ4ep8dOLxNTUy1G
zsqg3WLRRPwccgnRV/RTs5aIi91wEEnJz3XLkB1VHkO44SnQn7T3qCQEAaZGxcpIVXuvUvJCzg/4
+smtMQEpuyqX2jR48qcSFC55vt0PA3aYOEduBXTqXz+3ZsN2SqODiGQOKlVtRPCQKp1Oyn38tjs8
oQFLxSZzKyz9IcmOvpZHy/kEiNeFZYnfev3yxReL+bOkH30Ed29qGoQiROltJ9PMyOlWyqoR3Oy3
vKwOUzXwtc/hwBO3kl4AcaE/g5qD4JnPsWVuc4pxZVlZXDjtMGcotHBqmfHxflfOW7mQ6UbyqR2G
2fsuAW0kFbDtg3t0vuwuqf3mueSV9sCMd9bgUgZRFwvwNLFY+hsyBOUxWmIyT6y2f+daTbHAtMa7
+x/S3jdENfJ8N+XaD0O1UKSXreSo0sK3IkHl1SVAwHMPkJW1TNXdbKNNj352mFU0+szm3cqGRdvD
xdFU5yNXG2Hbd0f7jTmZo8CRcmkX2pKU57pvOfTURTJDXYVS+EcBsDnnM6AOkMWtJQnM0np9qfGf
CUigzj/Ilh6Ronsp7BkCCgRWFFbfp23dPVKKJbP3ZyAqIIDMTdBYlVqCI7LIwysiIRcJgHi+amf2
uHExV8i5yvj/Ud6+tC//znvfgPoBwMGxmIJJD1LXmWFtzfn3SspnUZ5nZKEvrl3U8HOnQWDrCRAt
S9ZP3uizlIqEw8FiHY6eXAZvFrJwp2l8S9VNngxyuv0H5P3Y7hmocpsE/6SayUMCIiQb0IkZyKVo
f+8mOOIf/Is2tYpr29cSPyzfXEuvBB+7A3nsohkHGvJYeKe4eB4+UtBCMj75nbk+T/2T7QNc7cLu
YmDZqOczB6RyiFPr2w8/q9HJYoJqR8bVP0VHBHI3/KV6SyQhvuaJDWa3IEnuWQkp/0+l+xS7VB1q
vL1nqYUbSbDJzSDzwjKzHiWaaVIAdPEZRrUxVTP6Y0qZqhZesNVG7fQtRrKu8xG4hIz3zgfw4oZG
1JZmeNV9pwoArYFiuGTAcjlP7ECzd2ZB0ibJU8pQqCq6tfXhxnaebbbVPjTM7Qipr/choswBog0F
CjrDIK2PNc1U9GTJqiKuHrvZoUMUf1rWDMTLYMSj+JRvXQhygjfR++NCyixJfYtnfIHoPB52Y33B
P5jXDjc3MwiOam6Q9hFLacj2vONvFLkHC3x+BKdDV6OIlpmMt0V5ER31ea1iezhwvCbAkEsl3V6h
aG32pRhQr1neced0iOdVKiiT8nGqRnhh8nuEY/Nr2f/yFRHaVznuHkyqPRDm0bofno7mkdvCn1YV
FN3gVcIq35nTgllZjlTrrR68nb+RvHmz2Je0J87/OChAeeFzcCBojQViNpc4LSxY94GBDIJ0zrAD
19cDW5FMh7P51Sva86QoWELGBTljOSyrpwuAvJVS8oTQR4FH9mbQaakC1HoYaUFPhp4mFmRlmvSF
0HyRFGoFxQRz9FVmeVdFwjYZ9DM3sZqbLIG/uWKcIoQd5hEb4Gh4ry/1/Bb/uXMWZT57sU7hVDoa
HI6q6VEWRxrOwhIu7v5RBSCtGsv8HozkcNyFpwNa+j3xHAWzJ3ZAusHd4sepk+SiUWLdV4pXPdyS
YmnG1XCvnCZiuIj7RcEDJ+w8ILE2PwNNvLy2AKNWEuRx9moAaePTFgl8NEtckKOJ9HgT3g8lrgSa
gnSTZiAqLgCt5/FFm9c7i22xA96vDqWip3dEUCvx4RnUlHuqwJeALHQiNAZt/E30cvAHrA+P4g5o
ycty3j3qGsqqlm6QgpycnghsayqQYrDABsNT68UyRBpc1Mom/8BmEoxtOOJn736SoWOvQQUSfrFF
apD1BAeVhoCV2G8EBIprFegC44vUmDvR3M/7HLcTAE3IUfdTuARTQSLaRVtkn7xxswmq3YTg/VPl
nxRQ8frzRRwEKgphwf/QoROblLTDb/j0/IFfPIyc/nwgD8pvW1rmi+AexC0Vrj3Tj4xDzFkgBxq2
OHlwBU/tLb3lxC+HwLpKuCPbGdNr0Ok/+kYZW2+YHIJghi2VLHMZjwoiNj0IuNg8ivAFV74HmrRt
VEBJYtdfWhJDkL/3RBzIdnqZ6RBZIL99Pv1bKD1VEdK/I++UXC2i/2AM6Q9IXw0XDO6pGK26MsT5
XDRRWHziX8YC/j4MaSuXpb+YbKDPlxueVJpA1bdrTR89UDShtyV5pQlyAYizHy9aW9whAClRN9WQ
N4w+ZTzeP7nCOr6J8fiYCGiYqX3HgZ5/jptP2fXM+88c9pUb7HC2IQjUP2cH8MyYl9GcNf0O4P1R
9XcimNVoJPJ3Q6zu5gHsy4k+mUWXg3VJjjhSYuAaxdQ2DvbhIXFDgZY4/6bnpGbMslV3bWONA73K
UKEiDB4MDUvtf1LS98GPHT6lPcoRtJ1Ov6yuPVhgtcXMZRaKPuSuNzEBUBaoZ6a9Vp5CU3Pu1Vae
mKLBbtOTrr8dqmhfTV6EV2LM24Ru3thFz818m9CElPKdrhCBSJHRiYiblzyUMSKfGxfWhHeuDIA1
EvI30Wz9i2srX/sWzTVkso+SCY37Zy3EO4mY9NhUDKKSmKmuQqwUuozPN+a1C16SVikCWEAhaxw7
E5pOMDrZK8ntnEo+0RRge3iBG1jvSWJzPfaiO2GS4+1JcE/4j1/ZSrN+LVRi8kgBGn9/CAuTHB++
nVC/KUMB1JDlvcEX1H92dRe1aWia/cV+SP65flMohf/+rBp9DrxVb4YP4JXpjJJppi6WrpgcQC0F
3lrTavHX43HQfpFMNbru6pzwBigRVHVql8rXHmzydMLmgxNRSnKi4BQHYvtAact8LUs6dQcebSGo
6qCs92yZaFGEp+bZuv3OU+Jih22gWFijOlFNkLoXbZ0ZqKoOTGuKf2LBXcO+1VvHqYEDyUMsYNe6
G6hbJQQDbE/WEkXjSxY72Ynmk09q0614eeliCvuO0Z0sJbjCdLqBoou7Szx7+adoHXHnoIfhDa0d
zhA6S/yaVN1q3svSVavt90liM6pis+MFFv9Kg0b6DMGOelDsqaMMuFLirgMfZltVXlgkjNe7tmtS
wTAn2n/b3ug6sYC99zu9qJ2Cw+3JkyMqqsZwPSlhpQE3yR39fUk69fx5EwSQfx+fg0BLiPM7Cbgu
v7DzPGF/n6XG72bQKDnSBskfHLR92RW+JVdYVE6uo+95x8+AdS8l067KjYI5G59JRjwFk7eVmZ1C
0LfEyTmagtohTdk2Mf8RBJmMMAHiZJnmj7tSn+ZQbyInsaEVxps5boxIsQTXbA5jqwBT46GVJAHg
sj6F/7HRc9TBkFsB5u4/W2eq0+oSy4LuneBCngg2ZzqozddtqiPKiN6d+y52yd/AChyf9Wty56z7
jg8YdR+6XeGVP5UE+0eJkO35/jERazRErjTtjMifiGpWnajKrPHeqf1CCCkWw4/R/7z/p+XXGAOA
QbjpHm6qSO7wkN9LZ5nzvYCzldKxJhgGz8caIwtIsPV1SpxwKK+1HvLht9OaP4D0PaF1hfV29qtQ
6+KHM8yUc8YEZADGDEow9EX8CX28Kb0acHW5aCkwV9NMLZT9kAMqnVLgDgPHdLMxE52zRLhV7b7R
hcuyfBbIDbmK2e109NSTPfEQ+JURJEffBU9aZ7zP0jaQdti3BYTvsI2ME/dXomjbqmI2O2+r7BqE
3jy1E/2GWGi0bKYKZaNGAdWXKt+N1Zx5YijI7//ugG3KHtMwPtZCjJyMNoqXlcXNrtGh5fCV7X8q
Acmg30TZLP7hdiN0kk3gbc3OM1M28RelT9/frXqlz63B9efoS21JOteueTO8RwRTkyLSipQAF7Ge
LGTxjmV2aFV0R1ssl5kIJ+z0AaHVNWhMeYTkofx0y73T9U6S+LEIkHgbsronOUuxF4HnmkziFUxu
lCd8+Ex8Nk+jZBAvWJuc3AVTvFV67hC2LgWtnVw0P6JRvp6IFb8ewbLcce0iQKvT2js4N7XJXwDp
TbRs9whGgqeZVh46bDZ1lkj5aS1rfx8Hu+3JwtuxgHNy+klfTLk1pzo7RyDltxr0y0BEDlZYb1kb
DCNvcsoJFjnA/bUxV3pRQsZ5akHBgCDA0sHpapOQ0A/lm0qsCT73tojmClNzBzPwMjqfzfQqS9N5
cVcUMPiNVhXXV3g92Tt5igXtdzEPhC4RpomkEIl23NbhfqZEamu5EtIqxJqEq7o5EM56kyUuItqi
NW1gmvcSMVNNeLMIKXTxal8uZ3co+xARwf0WiQsEnZdRK8Mqdlk24Ed8zuJe0axVO2mQ5etK8+9z
c1Xiidst6tmVxkNhlkOKNNExR1e271dbQzw43oIhs9p1BC5YNroEIHU38gIba5BgMYsEY0mjOMBU
bKvDB3M2QcYNVf2jcbZn9xJUreZirvSPYA6Zw/fqPFY8ixsrzZn+YGASUKXxmMdw6RX5nFNZ81EI
WE2JZBpykFD91USyD1UGn+/l/6qFlm10E2B0tAioWU6vP/mVsSfS0RDjbufeVEenmFf30h/lfBRZ
ntAf8k547Q0GHarg2Ga7P029K1Wz1Gn5pvLJ++F6b3vZu3Wv+X3+/7G9kFdDUeWTmQKHy8KKeduB
8vJdgqWB8QkgEDKw+qd41gOegXfBe4tqrBaZ6RRQvm2KVyGXv9Iq8jUaUH4dy4apg5DI1JKvMg6H
bDK+Zgmxu07t4z0ZibnfR8Nz+by6ssBfYCcc11K1B8fCzOy7iUp4LtMTXLBIbIGsXsr2gzjPMtCg
AZ+O7Pa8DM33UJmLRZTueck4mUQK9RtvmW81vzS0M4rHfvE4Y7WxDveUIPo4yum85u63dUMWSzLU
utnzHRFZ5gy2hYcF34JXdx4bABmSy1L1ndOjlLaubvMAPj7Urt3WahsvdaSCMArrhLBpHU7SJXPC
53zb0eMUkDrHF5SVrCNbO4h8y2HL/dkl4ewsmmBC6j4TUvA13FeUAnH+XzmHKuAneorHpFOvNJhF
mKIpTQVFTq/mKQqMRH3NdHeg5jgMpnuVqMIFIQYKF7pcY0N25yivaKLbAl7pRHaCnYrV49q+AZ1/
t33kUlM1dlGZYROlixKaWuazKQV2/BBmaB3y4Fi5xRgZ5OovsNpgbabnXhQ9cPKXbLDOhBdJTdDf
XRu+9qsYMIyLZ0p3AHH4s0fUwys4acPNh0VSLdtMX2Ko5R63iR2Z7h843ODk6G+njPSnNH2PZi77
QxgD4vdlUwp28X4sF3GDtdRAP0B7QjTXg212vRs+Wuvtp8LbgO6Avi1QUgfEC1zJUmBxLv0xdjhv
J8EFiNWfj8Pxc03SzCfgAnMJzPW/q2fN6ecdhtQxaRi4pSp4HGl9ymSu8ujMfITvDokcFvHoRHey
/hkqDlXH+nk9INT13vI82eaIfNrfmD2XP2mmkP7U0XepquG2iYQcAbpGxs+cXYCfPWc5yRKkfsPv
h3bSyDkkTEzp28BbFXAQXHGcrRhbkNDDArADQMLkjoQskXMDXwp/edjdpXltF94cVqT32QsGWVHy
p5pUAVvsb7cQSLuWZ+ceX//t4gdmABuhzM3HZ4TUqu8PkpMgaksgsNmGv91rXL21DfVoT908XaHa
yCObXTU+lr/WcAGAPwbTu5nCQNfY8GSV/RRrKAzZOMkBDuVXdceAOw8QANT2H+KibY/6ZlFALxR8
jJ0EMSuy0yeX5AZNVomhWv1Qv9jXHrzJ4Dg2Jeo90LDLBHSgwMJJCw/hjq2owF2Mtt1wD/330m+E
OiEuPNVqY89IBRY3xBM7HTUW4l3kZMoRiL2gOuAQOkrTu03gy/JQgwJAh2m18jDmictcQxFYLG6Y
LlJhirMZjWVnZK/3T6KofwPtwiVBuQt2DrxzS/TPWI2hFmt8/UvPQS1fea3cddpwBSExPoUb3FTW
H3AbhTo5o7HmEhNk/fvMDCfoOLzyOpzQ4YzK3YChdLX227FaKfqC4dhw9K7oD5K3VJ2DaPpzroLz
eokrUp0vkicyhSrYyDltTe+XO7mf3onwWddvtIyMomMXy+8pG9AIDOEzl/n/oLZsdwVmYkM4hKr2
MQ6y+Bhc0Bx0YNIhiSfhYw8nsqPQ2Ze912dkp4pP4WS5RjOMtKgMV0PMLMRfHAhUKb0NzotwV0JA
2pXrO5RXby3k/4Uax5NzxRrxUItSEHJnsWkZRmuZY1pSVeMFkDO8ubZL0GC5hqu/d31YZc2ERtgb
pkB7IGF5bd9q0YX2d/BmheqeQUXtc5Rtppn716z8Y6ApI5w5uNWuqPyC8/sMhcnG9Q8mfH0/+2AC
Dcr5tS5UXeLhau6mXnBSlgGqQAIC4INxxemc9a+cD8mc1b6KoD5/nZBo9/lm2JiuNx2OYyN8iCYU
+s4gesKGO4iiHDOnrm5sKJIytctMVhQbic78EflStZg+jgCoPZNAAFucGrsewNkZTQF6rFT1AS1R
iZqgWwnpSiA2azmm7nUBtJgnlAXqrkBQLLFDY7SAj9+LoCKHNZ0sUnDKLBlJpKZrO76l2uP8vSzQ
ZQ7bpvvayPFYEyFmS0R/SXiZrEjjsMyLJtwZjWRhAOljc7xHR9cPsZKhqXO37eNxh8uO1KJUtu/O
pfacmHolhIgMi77qBowT1aoFgxH1mmB44rz0E4dT3dcHcwSHzz2DAC/Z3Y5fbk6NsCStP8gdW2X6
uQC288nE5JSOUsRuNA39J/S4PlXnRoWdUWV2SbbYZoRkTgnQuno8y4EHbz/6KBAkifWlGYeKggjV
Yl6vi3oZ97hGzlCh/k9HiuPZ+E8WOBJDIOLkn2S4X6xAtmBUycSHE9ucBumAbARFBL8idm482+YZ
u0WTiw72dAeEEoyZ0pJ3SPxXFaxYyycE/71O5ceo1IcuwWCVYYQXmAJx2QedMGdX6PIhe6mSM86m
yGiuHwFGaU1LWd3vlfs/S6nfcTKXRy6/plYxZxWmMb//sVQq56XMpg6DuHr7PgVOwP8+6MqJSg6i
of8WRfl9TId+7LcEvpTkEM5a4tDfVL5ZxffFPUbBLpNOJWNCFs16ua7XmhdkTKo2A/CzZ0foWmCk
epp9Geg+lQ4KSm3gyXbnxAVdE1by729HAfOd/NExRtFspVH6Pv3hGPLoRKU491sQgokW1uHkELes
5IK4+SyUz6CB9uRebk1ztfGn6VdEE28Mf6v00PojmFJhhJGOj9kHZQHQqtypmq3CKjWenzCciLNR
vVfgpoo+hYVgvHdDJlcu1HQov8xXBcSrTzI79XMUSrFYhXfsLOHtC+cGlQ4nkc0bZHkLjokFA5sp
84Hz57fYk1NF2L2mx8Ksm0MDdR2vVLAaKgVhfTUDAbQh4ITmwxSlddu1pZFoPP0t4VnIAYzPvzcW
TBrbmwlZi1yuNwsDHkdoaO7ceMiXPRX74MA27z1+EkrUZYEps3jcOnV/Xv3LXiieoIrhNitI1XAU
1nJbqTr5E99Z5rva4zjO8IPdxCEioZhDSPqueICx3+6vybd7y1w/OvisnK2VwrtbNGLqP3E1X6D+
JOFA0Cte7xWketGnCn9VHfX6xVOMpTLxHll60k5YNKKs8CPI+hLFcW++PjhdZwwEmBzSoVxSDWT6
D8c2bFkBGSNWRcIC8idRFWc9mdWzGgZpzTmEqbjUbaHwu/xVkRnZ1zKQoPlDg1F02AkGNxwqm5km
xE/2IlmXvD5ypkFBzGKOYc4dJ2q6L+W/JXwg99PaWJw6L0Sior48VdChalXmfYu2eAY3tkIUH9GN
TWVtMt1wep+W2dOwogdJjXh2LqMR131UGja8DnWVr3ciRLd4r0VrronArJidXTAHo0eodSMO4jmh
aWZSDsHeozFu3QfJMP9DECmmNM8v6/NVyGEXr0OBckz0vAFaY/NplveGtEwpQbNIg0oPBns5qMe5
7xy3nR+/h+hooP/5CQAwBENShICgbxwGopokhDGsaGptUBE38txy8+UkkLpyQlFJ1mdNAouxy17c
2zvM7UhgKntF8KG85PfyINECbmjQzzbvpxKsVUsGjBosIFMCuUhKqu5KvfaE9fwODFWa8IIyzOvi
CW5DiegJeJUBWnZ7PJeGcC9ueRTx1Wko3VyLIxONUtmKlH7aa4j0Fis1rb6WX1Vkyzqp34tXxFQx
Nucv1kUsmJVmIyWuvkKYOASW+w8MjkYxMlxX7IOdyNg5PZ9U6DcGrWUz5bsx7QMBZwG+kukGqVXx
8CihbOAw3F8pMhLDVaSw2EoBViy9uFMfSL3pWIYlTAQNMo7o9LXqu6hyEK8WihyE1+nuV/qMNcZO
kJP78Xb94IlutW0xWu8PEdCU9YNkd31qL/ALLsxIlotqhfQgi4LVzppVkqXcIm3RALZ94Y2+7CNI
K+Q8jHzdVWXlI1fDJkgo2IwVbRN5vT4iztQZjFin6+6UC8ipFpTd5R+KfpUGM2WdnGosv57InjQD
PViJN2acII1EPW5+y5gi9EZW5jBegFAA+9MJQ60x7tqzDJSyzZ1qlmATiMrRdy4Vk2LTL+l8agjx
Ewpa8DWDDF+zpM+h1/I74sXWTaDeo+zU3DY0pk8x12Yd+/ErWd3QhhcApJ5CBV24DOpl1szY3RPt
uVMMm8nkY9piC6lJdgRn7QCNQzUiot1wWZkHBOhRJHv48I6oCY5fDQUCz4bcv3uMyN8IhkDMvHVK
FtR8tXrVHtFAqCWCxDK6dG3yInt5loeo6wa0dEVeRU6OqsjtAWAoSZsz3PAScmFbfHhWeJos7DZB
4CgGPmiLKpGDuMFdB+4zKIHVLFFSwckXH9+/Nv+aA64EwoBzY4Nw5bu2anN+1ImWSuCw3JSaOYxC
Y6kH6SzOOhEu2qpPCfHL+ON2/VQBn0O0uHr7QydmPPoKIo12/Yf5VaFeUcOlwnQmGnz++RUqPwrd
M1Wy+HyEthUUcIHeVyClT4OXl1w9sN4McaPflpd2J9B8v3byYKJCtQ1ptLxUJiidMqVPtL4mBtL8
CnEppf7n86jZI96dZh+VCMSADibEfDFXdmADeYvXiMyv3NrKb1lQoRKuIhD/Olz/OuB2q7UI6PFa
XMTDkYx4RhX3ruMY/pC3OKvVPtUa1MVLnpoRmDflXi5vXQ7pvzwYsAL35EcFalhU80LR1T2fPMH3
+roAC6uVV4hZwyezFCLQN/76ycHznpPTZiQxyltSqBUhpBjMiRO+3ib3KTgQ5LlVEnzzrhXAJcF0
axvFOONZx/9WejNRRJ7ZDKmgnMcuLvIgH37TajaR7Hjhnh7PK6oEndjVKq2qhxga4sWx+AdAP2Xa
qzRe4hXP2+gHAhux4XLfEfssFci3bOMLCNe6/n697D/SjIRbxKJtHqhdlW0USAfsdVk9QeOLfNqu
xD/e1YFsUUGTbzCPpQkh0dV1DfQqBFA55rg0mPklZufsEFz8h4NiMj1klZFeh79JG4dQNP0RixFZ
J/j/k7HLlhV3NCkCsiztj9r141kyJ7wRZnEg8t7j288hp0uEUGrl0LChw7VIOJecOHUKEU4yiOrr
AWZgJel4LuaTvjA2za6HHU/olp5TK4pWMTjc4mdkyG1Gv7PY6J8oN6+BM3XRUFN4bHR7fGnqZHvM
zg60k2+nTQ+1pozi9rEIPBtL4D3vfWJvMOC7N5HscDGiVGWlQtSJR1sED6FtPX80rvggDCoD7nIf
jYiEFk7Tga4c84WWxO8L2tmo4OjGF+AB/HvnHeKjjlKMuTPfjm5cS5whg6DZCm4Le6Zw40WEXa20
P28siyPqIJ/zUEYGSB5XEMan0JUInVeylpluKfON5YOM+0U2V1KUrHmXZTK8QgEQOk2J0tK3JNEW
1UjoDU9+tkaV3Nzdy5p0U+yeqr98QMSgfq1QIq+VvsjUZ7MBI17BAfpkAWT8qmZsXFizbWg6sq15
RJTzXkbTsrZFyykpiQ7wNdvv+et5XuV0Qr7RWmvFZqKL8wp065EJsGBR2hnrJ4UeLHFXyNhPwaMH
AieJU4cYZRrfNISrlf/o8i1ckZCz35cruGW2WcNxvFcLk17OIBTiVG2R/bcfdOezRDYlskwxAtLH
e5T1Ch1FNNnPCB9S8X6ygJtzagioE8BpHxcTE9gnXgWeM70/naC0Kl9WQpUUirokmQcWpTXsZWxs
nyBWfOVPL9ZcZg0r+p4UuAM9608grcf71ISY8YTn7TiZ2e9j9Kj2pxcU4kWNa5NwgxlNjZg0pmKE
kj1hh3Ebym6MyNmYbE9drCylI249Y6zdTAwUdhbI9AsHw9KmF7Zh28U46xi1EFcpvQAr6sZ33JR6
vBSVTKNB6g9rG36WR8gIQlYbZUeYU0f+XHiD8h4Bl2DGEMiI8BvRksc9fG3QzXPPFLFzZlgbv/pq
Bh5Lmt9WWSKxWiHsWP/f83B5003WJOzz67I3s3phixLDrHvKHaxjBJ0RiRcPQgwzuXJtETbC4p6S
RSoQo0TYSpriXhO4FgCMBrS+Ff4mpdwsJoBC3p6AG8kKsQyu5w6g000+Um/D8nAU39DWZB/UaRjy
k1Wi1jhMYdl1lJLJxaKe8jBVCFLvwIWTh2dwlgYUuGt507rYYc8Ivm6dfai+9i9VMp8KL3tGbITf
pUL3NViKV9LKFZLLQbEbKuKxk3e0wPCOqKSFx3hlvCiLKOxId4Vqn+sruAxH9Le80smiAp5ipyzC
ghl0FPl1bTD60WxG4HATkih8Z5tYpCjza/Uk660IGONjoVsTOLjODtGcVpkN2yxLna0o8/c5TJiD
0Px8bLnN07RxT8MiM6C/2Lga4KPl5KS66HxZlVOM1Axae0bGZb4OKpeS1JqVe2xaLkUUcXlXD711
9tW7A8c/9O5tFnu/G7/n68hf2r6P+NTlMeAyzT899bqdAHa54OdCMZf10/34VSsi2gJTjzq6E2fj
eD6TVhy3yDdgLTBHDB/vJ/t97rPFH+E1db9+ByrzvEhw/Z+wXxkpN+ICtq4wXkIKXVIbm9ob51Nu
5Yngs0G3MsLxMHOCm4L4oDSukTBMpDvM21Ev5l+0jSUdM2jyKBlUPblqXEBw1VNxDpzBVsRlnY3W
wMNDvevsylUt8J1935TP0pz5uwV6L4XUsVovGgWm3Wck5a6Ml61P3Ve5AWhiiLEFMziGfqER2uk4
d70Q6JVtaoPXUXDfenh30ePqLJZBlALulGhkhtO9XpHw56/M+/y0NggS8h6NFL3PN9WyI1kvyvaE
h+Kmn33nu2785gBpCM45lrhUdBmi2L+ULljoUmKGuwmrQ5/MGKl4K8x+R1EueMqIcQVFTqG95fYR
bH4PQUJGd9cqs2uCgnoNLT3CLMidsLlwVQWEJ02hSbtHEJAff8r2kF1uQpbrs2QOevql/1/LGot3
DIiJxb3t3Ek/uyPOyOgPk/qDKA2lbrCb0LcsFkpt2yRX/HTuKJLReeQncPJXzfX798CVMRKIy+lC
7iLGwGAj/KL1xR8ooDOVkmG0QqQDjm2NIGhP4GMowJahUQYF3QpJ7yCYnYQQPf85ppZQ7N0STpc0
7h2gCwL2aN6PaMarju/68ogiDP6xrNLbqZM3VECgfBvL6HuSw4VXnzj+KA11doPrvp49CFILFm5z
C+FvyQbT33r3U9jl/ThCbUGI6S2WpG1LiZPaXk331zKNuHQLzYkFDgbwAZ9kBm5+gjnWXpReXBfl
Jyhp7OuI4CDk1sf8306MvUxlxH3Ugz+P4PT1kR1mfKAbQ7PFZRsGsWYMHl8QvTlZTX6XLUl2BMRL
81qf1afdmsuMLgjuHCu7zVEy2wFyJfrDQEa2NLecnnl4ZvCnAaFA7CdaRSE0T0RpGTXF54xuqheD
czHoj8KJ0nhlaffH7VJWGKXNC+t5LYmKOQ5psvNqyYMWQjfjqUgz5LLYSG16y/zp3p1wmSP8DGOj
jzdK0av/B2WL+2fsenCRfokQOjLqt64vrE2FrX/r2orC4hl9hblaurMYWpYpK7Sfs6tuH+XKL/IK
wEYP2ZPxaPlkIQrW7xOLz2+orrNPcfXBXYI4MnhDB0RiiKeH1KjrwPVRm9/yKJXgXyb5OOuIG3TH
2KqWk1JXctHGGhw66L6giCwK4KNVAdaOwTwpKOAoacR/MQ0T9LIq1V4dqvEKkJwSTIcpltHlzNTJ
zglJ9J0nKnIfx1rHExvVU4aNM7HsBVhPM5/GQ72c2L9FuaHT1Xws9/sOOnledlkg1FhOVMfe0x9k
AxQI8Z/RGnnxEWa+rHWzTzZOPFICC45V97D+OPRRYdujd24XnyS383mBFXBm56S5lOtVMMnOGpqW
TSiq/oOnGQExsIZiQUzfpF90h0IIeIQO3LaEJERaxpn3fW6Anmut3O51RddRCl5hsNcJzSRmU+Y8
4ynwDgSZuVVS3fSTIYay/zSz+OzJdyDra8yOxmmgS/UdES7zcYjS2yFnMPD6h8ytpD30RsOczLVi
Vn0EtfVV65t73HwIZtXwzggiyd5JplwV3ToFNNOFs5ZpzUzwwnh9AXUvKRJDvFYso3pdaHl6SEmz
Tw4DFIZkvkVMwQTA/6aMNDPYAMKbake8atflr5xvG2XpA8FRutsPaMoACBs2JBsA5AUWn1W8jcnM
v65O0RE3nYQxG/ACcmEK8NSz+Lru65koRQGCleCat9yh+UOCX4XEzVX8Oag3r/qMlBD+VGXaI7Gp
Otd1hOx0ErHms1LLbQQBsCBdaf1/apFLLCp0m8CelRcbG8KAHkAb/TlL28OTFq8y3oxO6IcVm3j8
VXtvOjy2JPETG2fivpssUN80iq/2CEDWsSSGOBCYLHr/GYyUD0xdbS3dnfeoW8vjr5gxWzGO2ch+
uV8mKSbNjFeGIqq0T33JYF9Rq+gzkwVfjLdU73DUNgUX0jpjg2/B5PSXbO1bw6X3V3KSFQYyDO5N
WuEzrnmObHfqbwXKctKNBFfIRV8xLy/FTlZl9qkD7oR1VvfiiBbelO8cCeRwxk6GPQAtkKPqXAgU
pghk22hPYplykJhVw0vFV3lFlf8SKLithLMf56YcVOT8EGDzHfVYL9veIgGVhenuhkvu3yCl6AkN
s6ZN/SF0eKa+lMJkXRbo1WUXSuCTQNyL5e7ToxoALilQmVMeSqSIOBcIUnc7BCt0YrWhQnzeXeft
ZtAkoso4779ky3Vx62oEd38P0XJl7qWR18DARbbcQw/CvDjDt2c2+A3WlLj7M14A5wtpHy9zxhRJ
YoCXmiP4sZuOnV7ewGvaQ+8fwsvaVv6FzZsG/FHsGk6hioHWzE1qoDJ0V8FsdFbvP8jolmOQgLUN
/unQGigivfGT9OBu2eqtcW4OoXWQEo4YaDwgpClu+HPG8uSNraUD7savLGp/x66gNnhd9U7dqAte
v+FsBI6iiJOnzHAt9HFJBhvIGArJPrVv0/54Vh5L2G+NaVhRjg/jSjrkHMYMgGtjLVrV+0LVPISX
f13nSihGb5s1vEjKBwLGzXyc+NkphSPNmBBUgvloaSRYh/uBiF3mX7fPZVnow69r7WBciLj//TqU
ETvd2izxYUZ80d9smmj57J6oGh8+CIjiwlbWRdsODrinri5ltrygDboFRuK3HmMl5zIOxM1NBSWf
oWLIqmxK9drsHuCpgv27XDcbUx5CyVaqo7IDXiazJS5v3Gdi1fFeSSmFmROhYs5SpLubqi5PoIyh
HvyzDe/RD+BIrFtWsy+eJndU+RStlV/tubEzvz+0MmcCajzwVUCvnA4NZF3k9aVltuyr9wcH9nby
BJ44VF5gjTJUWzAmuA3Gt/ePJMTj2HYcLgDZgXbIObq8hwrBRWTg2COxIYSbm8GkhAkTslrr4eit
2BvUk6KC6BHkMRsnl1nz13Kwin4fLLnIZFGMC3nddgOGVR46o4kd6EEUsohf0eFsl/irZgCFqA65
F3VljdqhK2uELC+U1Xq6cwEcycOri9E021AQoMJpXPIRpvLzLuVd7jNJBQ8PhkHIfjzcwjFVqXYY
q08fxXL8UMwv8dK1EIwCob+cOvRFuZWYzIpMyC8rq0/uQsFXjkJtlqifS74cmu0jnQbINGcwXOij
dQHDbiHHlh33OZnRHoYyNvsFYz/gH/zNS2sTD20D12Td8ym/TBz7fLGpKxptoSlXj1/WuwbEhO8j
sD88s8UqTbjpoqOmvrwqXFA1VQ4vs7KRTRe5uFwD4ZXJLlD0CPwO9au8x2tRK9Ny9TctFw4u5/5W
r12sl4oVPFMnqBPk01xUIvutt8UkxBJmLHVe2nxXSlcAIBjU/GuNN3MSnW37IsSGy8PHBILmql46
G9sVIn/LmksFDir0dG67bUcM6H0JMuaIx7zEigP6CKtu2FLPoQhO3dY/kSK8rpCO/4NRkdnrjR5y
dmAY9F5cLmYOHlqkhCI9uPXSon6h8fMdaEhTL+A0JRaCxRPOCA81iFhS+r/RP85xmZUA8RIyyLU7
DIBaH39djRhS/2mvc2aRSy41HZq5uRruuBaxn/TMWU364hdZTHgb8W2BPXU8Xh9jlbjT2AAn0Eh6
ZSzawkGuIdr5MXkKSmazA8Zm3da+TFFlRxFNO4G5ii0XG/yDvls18kR3dFQbWDTjQoI1gkYhsKcv
yhe7UHiB1n3ueyzjdgVmZAcN9iVNLIFCi/OXK/KypOURF+q3/u6QCvPjXa0UWmjSrTZ1Vw3pFMWu
OUMClS/koHtb9PfaIZ7v5A1Kt/dZ0vEMiB3ngiVlJ2qTwhRa1eZarft0yUgVYjGqTLDJlYrbTGKw
wh/AydHZiseiqxQr+f3wTGWTqWuAEx7uLVsNXguj+WW/lq10xr4/z7qbWDpBjKSggyJkuaA/QymS
NN2KZGfXzVDhwQYfBacMt0q/SNzYfwslGaZwBE7lBSaH2SIGJSmqJ4ooR2r92TO5yt+PghMsWWca
4k9COmqnEfPxlw+C+g2JYnUphj2lacnoUWyzXJBrb6C5TDnl00sO6/3dJ6RxQwOT9iC5lhCDiIzc
WYnQna9GXfYL+sfvOpSRoJQMKKJlnAM1jnY4qWy4rRfgut/CqgJBZYuBcCERObmIZip47FIh/dj3
l6ZEe/9/FO49UW0op9Bm9lm6Q+LT3vDX+D5kRoZ6E8+kTRP+RaGo5vvU2J5uqInyA7hrYqmJj5XV
VNOhHHvN2HaiquHKx2HQ2c8XERCwHhBZWu+11cUulprj9k47tBrNDhjmFA45K/NDSvPV4Cwp+48o
wUtdKO/QcUhL+fU+nc9IBJnjt/4Wxi07Uki2cbVN5+zTEYagHZ+42+pRcgkyTn966z3W/tMyIXMz
5bGkRXFKCFF2FMz07Al8kgTJ6G0PDMAHScIjTZuuGKjBZSmJGFVG5mujvQsUVWh2OIh5SQt9ErmZ
aXH3/ZBCkFXEMRXZXaiR4Fp1n01H1G2DDNRM3izreygfxC7M9I1ymelcAbX3FeSROt9d8MuI0esv
Q+48TlRJaaV2IAK5Kwm9j2wsFZSjvk4NmnknjGszAjbdI94gRdA1sa8nEgPkVacU3uqEsBJfOyHz
SEMY1v6b9pe2VxhJZnMGwv0yCTHb8D7JmlHwwD4qVPGt0ssVN4isS8fbXc7NceJUSYrzxl5iwqZk
KohaG2xX8Ah51zUvN4IE2RkRQbEJLy//XVZKX4jwU58gV54J/wflIVAvjC0EprDf9eKxuHNkIi1h
6QWx/5vNtCi7sdmhnP7+EJU9tkicMfqpDRTlIca/mQ4FP+8K+g9DoqxbBj6xRLKC3UttkNsvAyYw
Vn+j7x9WxHp7kyiXhStBilf9MIe0kpJuLEsrFs3CKOtbKI6CEfWGWGzMG3jnUA+0eOP1x4wzfIyh
r0AguMq/vnUVtvTuWXtyASzdE3te1b3ysCmGkqO3TLccnHcm2JqjTvosd0+3B0tbKSx3dLNcT5BZ
P0KcuDuG6QgR4GpDwb2Yg8oDsgRs65WjZrtJoJyzlFaxE6gTCUMhk4x5mv4KwtcMdLAelH7IyyCd
vXKOG8ObrV0coSK+T/QRUOBUt3decWxzzwfmcUJxCu7cJbH85sd9rGOiHLh4bohMBQ2f8/4/VIRh
Ca9KY940Hs5Xni44YU7EPcDOCshri84/eflSTxU4aSEe3FAp9VwqTF3VSuyiHl1B8LiXVsP9jI9H
wwBDlfdeRtOhlEH45kMNgJNggnDEFb/zImbPJ270QNEt0gsI6Vapha2bdcqRWPWB0WIynpQiwq+Z
jl41WYLfsYJnCsRm50vR/COCBa8A0LAz8fPVDi51WEQhk9OsSaYKTxy+7SEU912Cyj9IXhgIgK57
1TWM5sAdPFpp3rFd8+TA6Na/Uas/KEaCKEtyDT5+RnFC21A4HnBqPTYlhhUbfs/u2nPQ14bNCk59
O5ZBG1jvutjmQ5rzwLC5nLENGMKoUGMXxMLT3lDGsb7zFy1nmWt9ZmKyDGsSBwHdAy0dzzTF+MIa
Jkwsj1D2G65f+SqfXOj08KKKYV5e9wEK7gSPGhSm6mon/mSqw2y63I4/Ggw1cwoccH9zP9960H7F
33voz91pj9RoQVIKbsDNl4z1y5unIF3EFJ2peSySdvvC4XSviegsKQyq2vuy9cpuyUznuykp2yXL
5u32U77WLoDRp0iYAJHMXYK+SzjYUESuhrqDCqcY3XY7rmG/5ye8LLvhZZR7FvLBg0I0nlEfksML
k9F80wAAaMDjSW9wOTcNTLR1UMwkqk5t/bmfXMlBPakbhBokVP9aLMZW2tZ+dSWh6HCWZbX0KR3A
iwOiQYhKuCtChQTE71Lsds+cAzU6r45MGR9fdxkBDNXEkMoS4tY4AuOCnR54n3Qe4/QNDGqVCrE+
gDNmE2zoCmj9p+HXs3ynprveKtJ3wU2IgHeZIadYQ+K43G2JQ3aE8nvWW72pIP6Hu0Jd3H1A6Ijz
Rkxnreyk6KBZFtPthCz7OZO7d8ig623hUkTMdFRVCwZ85xNw5XYTu4ZImmi5SNkD029FUw56h6SO
/t8lII6NwxKXvaxD2UVRIcMiRTv913EledQ7SD4aAW+5O7En/je0sXko84qCW0KPVVuvPLRgLXI1
ybEoHldentYsFQgd/7Qv9olmjg8u6dgyk4nppVV9PLbqjy4DFLlvQg60v5mYcW9CLl+DvfB7icgd
gnxoTuLveSqKvRALPyWIcxZ6P2lHA5lGHOBnt0zABYUmWswSNYbRP2TYRc1DmOZYfBnWLYDPN+BU
XIcYoKgRae2J3YUNq3B9yPEI5A4OQEIbMrtx+n/BSiAx1JUUI2V8c1quPIhqz/TbHpyYgyFlDVVE
FoeLxVDsHUF7cGvuuXzKyRbGqGZA2FaQ/JDzQ5InyzzXKy6E3t9hfQL0fRB+RXlZHEXHGM5hOx0i
RT7TdHBOGR6A1tzV+3TybuiNj6NkirEaH6i06xNGqB9BG+GulXZoo1/B8+uw39JsV3IiP4If5tAA
fH96WnwRXGMBBoZKw5qV7eJfzMpzUbe/j7Q9R3jBHu5vxT147ifgFjTej/SOdPr2A6pVF+KzEvU2
bTeGVT9vELci9iYlfTk4TzuY3DGpZgFvoSVALSd6x6wyrlapnafRLIpuBuUTPawkXy3B5iFk4B6Q
E6Jxe1ARgveSxE3TPMyUdFJ+Gnf/HUQ5DeHY353jeGHclH4qpIuk2wsXHZSStv5h/4JYZ5GF76tn
JWreLq0D/QokVvQ9Lyn3ewzCOaSVWx1OpTe5vNP4nUUYzplfS6dCat6TGhIswLZuPkdxV0vgJThs
3lKl07X0vRtPEbbG2DDcdYGo5En6y9k84+hCQBZGhW5zU9RsJS7gBeqm1szMC5rMmRin6QiDmrtR
xuLUmJrWckBmEzR3c2f2Y47MWk2sbsCQn6jfJlDRS8m+a/L37aLKrk9SezWZ1mxrf2F6kDlEKodC
jALgxCYOzTLwn/H00rZl8PqUbC3MCc3MlNzhNjSNGYrw8/Oa3p/eSjDUsxFWHDHMIrMY5u4gYiqO
BEe9QU3fPbGjxmldH07BFsqzNBmFKyVBL7XhNNgIdP48lK0PxS/+35hZ5obnFpN1ZWO/3iV5Eb4Z
YWWvpySjclWcCmxiv/CLzC/mRTBciOqoAk4alRq+iJd7HCbPf1U4Z9882A1EXH1qFjrTO2T3et2l
5QFj0lLVygbtnavGObS2HiMf54Dx5RbU0cQ9J/1BAx+P6qpbOFdjj01WFmO26nzrHNncsSrPFrcU
yj9vf1vJT1Sgt0CYpSPw9qCRy68d3rU9vhuIpKVyQE+yD7jxDJVQYDaaMZb+8k47wIzxzDcjfArf
n5XjgPVUD5+QTWP26Tvb5f50JqLGDT2JkxXUOje4QNHQx88/a2+K2N8QWygnna7oPalsXEuI5W5Q
AVN3gUQIN46XGidjRaQ3VLBuCXG4ZJRdrIodCOclBeDFN06ZZULCiaSuYt6Sb0f69+UhCZ105MuJ
PkA9v/lD2lU0ECBfgo0N11OpBVCM8jdF10rK2O6j3xytRKU8vbm7S8BcajBnSnmiHyBA+8JYr/nH
fiT2SNbJo6uj54G6qU+emTbLhQaqg2199RHLYorX2thB1nVkiPx2NPMcs3XKMSwcqkFDyuv1luz2
zF3xLD0dwMDYOBZ7hiRd9O9wryGaqpE9nP2sfQqqaSDAHoqFuT9FPucdnzJFQKwPCKvtK/08Ewie
T6/M+khsowYl5bt4/7or+xJ6CTH+2I+uHz5ry2JnkVDPFt6w+DSWPfNtzCMkoSciZpBDSSpJNCOL
cpOmR7wXqN7Y0EwgsgGkxOae1KROo2MRtEaJgikwI+GMLoiuqMpFScJ3fg8T4MfIB/dTU+cV5eNK
n525lim2yOKefeNTP6JEoHssKsSCVfAR6556z6HamWlTqTo+n18HTwm0UY5+xovlTkJ7JNEeFlkS
ZiAUUC0YjlYfqXLsaVxvAj5lBPqWwWxiyoxs2P/EYzVYsZGHCLoxUfRxdOaNa7lvfTULNA/JoXna
PQ32FE0aox4LMwD8OvoieTrEH3QF7KTGgpOp4rt6U6srX3wN3dBr2KAnz2OrOOfRlPvaIIFgP+u+
jw+DpUq1z9khgKJeNegiDzStTLFS2dJBk3PydYe1bMGuMT3oOrmJdHEq0WzChUtFBvmHdPQIc4x7
UWDNUesNPytlHV4JEdngbY/5/BPYUKeUes8KamdEsZfsTG6IqGZL478xeI2nEhMlSVFzciZF3j2t
E0uah5JqY5VJ53C2pCVKHjj7hfbZwxdDoGP2mSAB16KJh22mIjYD+jSr5ae7aicL9uOLX1L+zipn
sXxfmRgRtfuQSvXV4EKXX5h9T5k881UdsRgTXJUOziyH+jgs644K1JLH1hORqQbtpZS2NqB7XDXZ
zjlKuTwbDRnPd610Dg5wWJzTUSKBfUFceY/eyuByLiTwZSvzTcRnXfaz0USFYutTsxhhgddwWqur
3NYFtPUMTpFE0K6XOcvaQqnfkEc9jX7GHl6+gjE2T24ykyJb25txQq+ZKwm/0RdFI7TBIW7U026F
ndO1jjc1+VB0KRH9E8ma2zrDLRFJAlId1n1qhH3x0DQ+OG2L/6/+K+7zblEObc8JOtUx3o5b+dfN
vaX9L8euY116x+2/EA+jGOp5dhGfa0xlfoUd0h90JxrZAf5liP/H2lK6jvlNC7NGJUwbbkJlqJdt
6py2zYh5jBjXFAdc2DnaisAdSMZDbdd98qYCQ6mSb2bWiK8mzICRU3q2j3lf5q57CHTbnvI6Ryi7
ItHU4BN5/YQgVBMawsCTmSNS73t6mge3tWIuryg3l4eCf9y7WDPylwqUIEvMon6ofO+OBZTIzc1g
uqRjifVoYwfZ/zBesMf/NKo4FQdf6gQW4ayZWDGIjPHkGHIkm4s1y2A26/1RHwvKfUUb+SW7NgLp
fDZDXN5nbLQEiwjA2z2UxWm0a0vXqP5MSsD6Pc5ouKEeuTiWlFtbZAxTL4ZwkxdukokOYwj2eM47
LBx6hQ1Lsjevf+fvzsZbPgpcZtxiEwkiwgDaLqVRFR8j7PYL7sBEQz4ePnEEbrLtp4xrKzJlmZeo
qp0QlzwUUmQy4TJYtHxikJS7q/9KM/lbMDPpiBLnLGZN389QZMGTlJE2jx9rZUJsWKjV0rtjSum4
qEG8t2bCStAr1YOZMAua/bDTfVjAhB2tPAnUJ3uiDKisH2I22aoPns3LQUgF3krTKGK16DCxeG3q
MbtuGnD+MlkEVMl4TExX7u2GepLYIg6tnJpt+P5yVG3S7Y+1E2SXxn272u9IEbxO7Ph7k6jkOBIe
/fp5Le2/NhRIE0pPzONb/jfYxeacJ5sr3VRH5dDajjN4/XkKZ5EQPiv6bC4QFg/b2qySxJImLIpG
HUyKXK3pxr/8ZTvffnjP16mIyXwx8ujinLa8fzBfb0xpT46SmFlaA8jKMpPlmNacQoR+9m/GiUCW
wxZPjMxE/4sjWxYD/4qlI3qNRJ26IWlBgF26GpXR8Qg00VFr1cgLMOhXaZKIpGozZmfNoAWLHN1T
eX9F9BOwmH1H2+stpLHvFpPTO3aT9FJay9caUOL8ob3+t3r8nFIr1Bz0U+TYjy5h9EzBjmeYBsK2
ekAxXn2QLRdRDhSZc8YJGPu/GeZkCB01QMzApZoha4XAuECTz5bnYDsB8vk1KGLWKxWLcAWsJWy8
I0P0TX2sXEmD4uDz6i9jfd5pVPOA+JmIcrsoMfhU3e6cB5J/QYnVyPSBdmVVaBaO3PJErH/caXiy
biW1AHymM8Wjg4jnQ38XZeeQH8rTtFKXWL6EBvlOMQWRI4pqgvpj/7ZjD6fg89jB9Fqpzb0OxALU
aQAcIUZb4Y4lr8vo83EEu7ZWxg2Jr43SxoOhbYyzpwRu5R3I28HA8wcPEwfQy8uA2EshtGsESh5o
3dZcV7BbQuxm+8YQYEHektzpTdFZ6HyoGIKKRDBF9+kPf4BFSpcZoHyAwlbBLfu51D9BA/xLgd3X
MdAtB8ycqqibqdk9iHloCaSd3ealQaGw2JPzwRRRUs38uNx488oovOS6o8cCFOHxUJKI2X+VH5RS
Z2Yy0SQbTIFQJ++T/mJ2MgG81zpdPQIfOcwDO4MriPmiTLo5InXRfUG+irKsHGz9/Sd/zHqSTKYj
uJCRVTBVKyGYFY9TN+VOMKZzm+uAWHVVro3uR9CJbIn/ngD/olsxZDV5YDuVo+Yy8+GxZopPa9Yi
c8tD1HDuoSJ16qESbn76Zc6dKTQPtAVvcJCIxx3+qsJNuEqRapEiFvF1ReVHll5SA0d4WHakwsyH
xJxmJo3UvEHqPHiaFWdxNjGnih9Iuk4eRVZSt0kcRNHFMgmAbANIIVzq5axbCqqjMw9zG/ao7jZI
orUgg1co8trf8T/gDPHlP1Lgidnz4qh7d460gvmSmdZyQ8/YGGWsOwp9AIfgHG1V+NdZpm/VALcJ
G8qNRs1geJ+/MQaeXJAqHKaUj6u7jI2aGfyi50TRGW0ysYrny2K/yKZlPZseZsOUClE0DayoCwWQ
O+5pDHQGZJUIaVDsvC69NZi6PgVPW7wNGICCSneQoSIxgKAZ3DMhQsjKxPLS7ecf/bjjh86vsbS8
2SiaJJ9KWn/S6BI5II3zA6aYHKFy5s/KCTG891a+Wt01mSIWDKW/YQsZnd63uVNN0VIJ6Orl6SGD
fcubYeKWPpRbOhNx8Ik4/X0Bkh0D+xRem3raDy0bRdCWic3dqm2lpIenEZE0ZJC3ECA+yhOTbR6m
hm2Nt/IR992Jzio85fu26tFPATMp7DTWTxJmD6n3D5A2obxd+rVrGcBQmjIVej4QdGAM64ZAGEDW
9RGxIE2whgyUIx3uxz5nsNjWcqxOHj/D95aAkbvdRwWdrIYgwsEUqMQ0jm9QH71BjfVC5UVeLbHs
YLlfvYv1KFo1Io+PtG+VUaLrz5hUceh+drbbYZllCGfJoEciD96z8n3z9puaQnEGMI5a7CnfaU+v
1SBlJROneWB5M1Kk88TxkMBUd7lvR/E7t/1yvTjiuqcOWqDyPONDpubs3Z2PewtiSfK7EhrkC283
V7NYi5QtW9XS2GvXBO/kv3AMeorZK9GSGsmibB4KQcuhnG7vZgmsF7TGPRia/gAWEDmtKoFs8vDp
eTn57HEsBz5UxkqlltTfiphWKpPVjHKIkad4V1UwFS9g7dVOaLnxJsB6xNXus3oWob1GR9n6utqP
X2dQ4a3+45AwDgQdyTTSj2xf9MZ6Y6hh5dmeuMxoV0HrqB4c7cyKj2Lajo7OHrmyUCStaEA80a5G
+VzfmM0/soXprTPfFy1B3lEhdhhGic6sUkJTe5bKBGZh5SZD4COOXWi82xsZCKJSocoES4a9CJOC
cp+J2+GO/pxH6k7xGxBh68Xo/vUKHBLvaMol5kh6L+KR6AJeklUYuIzFPp7rqwjxaUBFGm4l2aKX
Ud7g3d2MvxdxQHiBlIKy/NEhMI5drlvMz1z091CdMhmaIWzGsTLwX1e+iGj+Tdf2kiC1bv3rBMgY
rDheIvwnAFGCWSnmiRWuhD4vsPQ0nWq5m6CMlClCf/PqQSAG4qtJdQDClZSL2ztqcbIrx8vPSnUl
E4dk4Ipp5KFoQfyoUuGUVMhqRNQtrUSNsRUvBFFUdTYEYiS9d14Ljevdye1iXt1USiHkoibSE0qY
zOfYBNPp0wfsn3Z36fFX3867nVkV2DkHBzIy/DjSvNfUKyndvHgBKnh/UCg+bKCrlsrJaWO2S+Kc
AsX65cP/TjpVGiF7X4epAA2b8A94EPJo3BjqMMLv+r2ZR3p5v0xqnwgvl6DKoWG57BV/FuJOAPTe
EtXDNeeVBacbQmXjVCh6FgAfkd87+7btPiYQyafDwka8c9CraqUjVzH281nuO7hMfwtXN4rquryw
ZE3aCM88UxxVPbQ/9YaPxwGUgY7s+o2m55hamG53swmn7etcFc2U8x5RJC22IiRDIIsl1qOHRuHl
llbyMUMWKwh8P657MPm+Nc3RGzPEQReTm96wEdH+Ggk8auuRBgTW2+2etZbaiCxKoo7XgsYFOCWT
XS+76vdVgpcRwMOTIrw8T+yHuULfi2uxHYTG2L1kB9yfTXESRTKflIs5PV6PNbY21C71+adaMIVH
Z/c4ErM+oMDoch2sR2EDasglJ9DGsoPt8A9qjbBHnQqrzWm0ZwqRIVnuFF34mAfaaMrWP2i4o4Ig
7DIT0zH3zwXAwtMKq0b9VdnEBaZAA2LAT3TJfO8qU9VDX2SUtAZ66efHsh3z8nkKoRQQiApE04Fu
HC1o5NAo3KhoGOjpdjfNK5XMV1U84mRBAd9BMCsNo4NvzcODL35Xjx7lPuIALJaIpZ7MHqEG7GAO
AXDW45tAEfuLMbh3RfU1jxD+tUI6kF+qJjb1Xm1GItfCJLRqE78wg5fcARinlsQUyJMBvvluSObS
U7UOuSKY4UVP2G00SxaQ63HRGTbMN1N2f5NiWG7FViZPJADCIQYx1+T4K4aT3KGU+kWnMiSYbeKp
yD6tgQRWIzI0B/OS8bMTCxka8IfNBpSJTEPpDAZyLRiv8Gy2SvsxM+FRQ4+yWZTZGNwSGP+G49r6
xnnkq85MnTVPut63Jtns/nm2e4g7McXVZnCOG1DcKzFjPpP1Q5CRbedxIdr4gvh+1GrE4hDgxffm
r5rtJMrYU9ZmM0UILqm8k30bPgs+lNYydhfG/iS673+NqEieSk/wSs0A2C+R45ivxQsve88h6IHN
sHl8eti1L4A8YjDmUkLaqtTXZGj4aEDxKC0IiUBXpFAY4JSO99NdD8b7uHLnb3HRaJcO8rPWKYSx
ZqZnij/a/ka96EwRH01q6U19cT3zMKeDdV/scDocuYE8uHaF2M8OGmzle5UItcBGSLIZY2c7GUMi
zF/jKMuA/a8kTAzdYJtDcqEADhWMNrep0BOAr2z8KL8zWKIyNcQBHEVp0z+/Ok3STS226opzSi1V
5UNH5xtxXnaVMXbG2WQw1PdBf0BetOVEWfZawyFy0PW0EsfjgRDOCWivbe76pDcvZwpZD+JWDHn5
pmMLG2qanN4V8ftkfRYLPk6qKabWdG/88TDOruqJGesfmcM3efunvS3VKNdBByaosWo5jfCcUMrM
wx1Gn7lsoK3Xd998gX+8s5zdeA4DW8Ed6P61yM1H6L/gLjCM2jZHoDih6gdrEGoXYKePJG4It4nt
uEGNoYzpTJAIJduiOX8NEyMjBHgoUalIOZ59vHcfiKEDl6GDOMvFwP7PUH8xrQInQuQigwzDYS/7
4YTc/jWXPTpzZONYV3+vn3/7jZxJEn+7npxYgBLusEceMu6J6bwlHvCRasFG8e/N16UweYwJLkME
btszlz6ubJCr+JTcmpOnRsAuMPIkw0M+RjhlRlNG4l/+ifKebworAFgnNZJB3oa+WTpRVnT7Vdbb
wDWyiJ3hDG7FHAqAsCSUO0mu11krP/27psaT4oHESqZYjJ17lY3M3mXh0hPLisHVqvxhVTVuaqsU
BEOe2IAzWBn9qiJ0FVuExBcERxMURGjSGHguEoHKFmac0ba/NlP9SknCbcnm6l/TDdo/IzkHY2L4
Y0wLe1c6qdnUC902/ZimxKBcVXJjkvxw937MBBMaECZ34ZzJUkDeJx9HLzrfjzk+yeMDSr8y55s2
DfQYBc7ku1B2cX6GGJJMtZQpC5wH1N6IJM7gyztA1hDz1zvKbvmnp3P53jCO4zSTkyAQop5vgQMo
R+Kwdi05j9jq++cBMXnx7UFbNNYIilOyJBfR1TSnBM8R6yEN0NS60MnQbZ7hT4PJjCkJ4CYK3aII
vfpsf3/TJ5Ulice5hGSxi5PDchqu1RpWRcF+dZUoBmpq4FpJituYFz4uhLiTijuHo64xOzmbmpdT
tgH3pB/q+speDilzPCAU7cbst9aVsSLbEyoYsfHDH+X9g6xpUSyss0+LkXVL34SmwGZayLoW3uvc
nig/rZ+0MKrKyXBp3nST55mNtDp9Jtc5feR7JUSq0h2aLtcwRUAXxZjQEeaWJx5GAd8aHv2R7Yn9
cA74KRgVFppM+ydxLT4dQQ879Bc8RI6Rg/Iih8Sc0kANOVcwJnYoe9VSAWovkYoPNO5KLPzMLNX7
Z0Y4jAz1Ah0x+I7LTxRISbQTnUYvk9y76mTRjbKi8MhfkTHsg46PISEzBfypOqDztkgyq90E+4PU
UXZuZ6WN9iDmzng+tp8sefQPbfcPUTqdCVmWkeiPTwC6aD1Y1zUwmAOvFcAefqOFYbV9OIlNnzjN
5joC63r1d+lcC2KyO0mO6qUXP+AvotNtE8fO1c/QLgQ9slZ/h4r4783ASYFxRcg4IzH4PrhYNlU5
ujHsopRdtZzDIacfkh+tFlnaL3g6HDdKjUBQqqqDq7RpkkhEyRyRA8GmhOccPd3cg06QzzQRIuk7
9eHmvAp0YJ9zv965kBgcBvPzHPjykrMTSwQ/FiJlZ3kd09u3fUGeWZJnMvNMNK6m3hATzW36loN8
ohKLSap7nMLrQOmqIxdkF7J2Mtfh38zW9evFl6tlURt6UwbyexPMitB+WfQCTv6zjin77WUnRcF0
coUb1KvWsgN1VoBbZAhuY5MB3Vf2R4OWxJP0zdDAauw4TWzVK/gGCTayKOg9sMZmBXDH5w1nB1Nb
E3uess2/rLZozd3Y/UQG1+3uM5DbcMD3geu3M4e1B62rQKViOFeD5x8lUxkcRYzRBAHtjkQExhZz
fzk5yWLbZtnSsQi0v3xCPadf456LrhHqGA7r3+rwpW8N+5aBcvJbWrmcSPkH5DzTEhcBq2uvH4b7
eWVG01/i3Euz+jJ+0xaQuhvW3WqZFnj6NdHVxDgW60wJf+kBs3bzyqkGf7L6AzsNLeO2EcwQp5iY
i26z7hbWTmeowgPGioEQnbHg2Fpm5mKOCuEx5mAyWIBDNZWalf1fNy5TjqCYnOunY6dnMTcQZiD1
jHFxNGa2688hlB+AiMvugeTdkn2S3fbcd/e0Qt0CuhIKOkykHdoIXWXyH1Wqfg1N88X9ypJqoHIn
WW+SYObmV4GZNCQtTslAthhzU+MNFq70PHj8AysH0eMbV7z4QGHmF67DyjTGVQ4TS0d+wLFThfYk
3uzB6adnAYU0eOPuVaN6Bu4tXWausUY/MvZ2suklht5i72JOZsNCrZT9byKp/8XUz+/wzDbQ7+z/
/dwZyOrumFBZx+b7QXhj51mYXSDB0LGnVtHhG+RmJYrtnWE4yOLgMN8EMFGozO7sGIEsWM+IMENK
MUVixelS/zAFBWVSMqI1yiVmJdMmIe8D9TNVvsQw0S2SxmQtsiGRks7JDTKIgNgh++UMYqwLekXV
MsUjSaesms6YTtqTIkhK6oJEb3+HQYw4PvR1zh/rnhKAkHXA+IUvKlTyqiD13hDWVZnLr1TnU2/q
wD3ZKVnK0qNFG0456+gFivHAjvQ+Wr7Yc964FE+rMr/jVdMkjejnASnj69cadEr42hNLKVWieVhh
UhDUlr2+ukJLod+i2o5fWpgRhM7PVTZ3TDzgVgvCzEnMkrbxEXF9ho7ZpshUK7sYpynQtaa40+l3
3wAsea6BXYMSprb//O95sw6xz3hiBOjC9FLDvz+lwnO36fJdmTqRe82kK0sYcvd4/bpF+gArFtCH
l9yOmn/5rxH803CSFceER/sJ6WqYkzYt7yFmf24wzcx4BuBfwmvQZ1QpQhSRUH5pcwSxW1ftWpYw
5GC/MZNXDUFtcPkKrIzR4e/uAO1W3rXW0VU0vQYKT9SKdeoHG047HO/I4sqXFGEhmXNlfZvFOMBL
BzO02/R7NmS8dMOtNXeOGB1PTHw/f8NiPALF2qt+vH88tXqYBR9bOhgP0LQT6ZzOJtrbYgLPmxWb
XvJDsySqj+fpiZFIYGpkQzMaAUI7DxjU7jpHUK4iQ4y3xVnDToXlqxmduSwRX/s2FRm62xTm3O47
qd5nYvl561ZHDGC1ruoklEof5lfTpQJys4GHTxOl/YkIZfxDrEMN1QBxmI0WS96Pnva/ZxFo5vLS
hhupsk8YoeRbVR9Adx++iAJHF13g71U3BExcagDoZ7cAuSpKxyyoNcVZKJoscy5d2O9RndUVG+Kr
BcAzk7NntSahnRMxoPgO9CuGLt7ZR51tWslDoDjk0ql4E6gJ3OQvQQtBCFYPJCsxk7KwRpKCkU9q
zANsYR5IAgTgHFEHBfnVatfpDh/+o4bLh6vI/nBPh7W8vSql2NGfVJAHL64nzEJ2au9ofrd5OTnD
voFXhEzlDqmwvVGMG68H5mhbcFxMQ2XuoGpb6xLI2esVW/retxb6Jdh7D/c/OTiTQz/GZijxWgCG
9nORrF0rxvJQeCEaqP1wyl0K/XJSwKFTO89aP27+j9W+f2qsY+xzonlsTY9eLi5RDOx1nBGLIb4t
1VvzCIJ70IBb13iwRL5gDMCKARkXK1SXnCIHhmwyKINWV18drXMEjihlitXbAOd6bmRIH3YkbvxQ
KYRG/a8nnVBfli/GOA/FoL5TSusLdEaN+wexaNywgzTUI/KGifd3Lpho2guGWJg+mY6/FPGaLK9h
FvevICcMxIewacwKl+wBEcD6ZvvO6r45evmFS5rQLBa+5lBO76Zsz2DDmjUsZ2uEA9/esxCalaEZ
mxdmIz4i2WRMxB/Wt9fvcGQmv+XJNUNznmsOKFsp+of8puROXeBJ36koGyDJqmEerUKj53cHP37U
q2irsBLYU4YvrMtEyTO0T7G/P7+egq1MfPaBHUKCTSCTGFiiiKxuz+O8NsUpTU7hHutAoqHx9M7g
6IeNClHxCnYKVm8jY6LGmaHqBeTVRmhaBZbJn4156M6GPE6iErpuSoeBpdKm2R9rrN/VD0/Qv/Ha
dPqcGFmqECfzs26GSiKmCTZMr/8nFflrwHbFvJRQzUV2koCVriamKoq5OQnLRqSmZ7ZH16dmowl6
QqWe3JsX20G5mmo6x+aA8mhwOmqh4iC3whcEo/py75oyuSgA3IICEqNHI42EJG3xBds5zo8jTeVl
8EqeIZ7zcp9cYf3ECKF7sLBLjiCrSr6NSmP5vFINfxfaaiehdMsoBmqqfCsJMtmLe6CYtTxiT/nI
W+ARMCI+0CRykZJc199C0FPDZCSfH49xWB0iURtFxEBaLjRMAo5tA8CnJdcmhZJ3UPVfFmy8C7/J
jx9iE/SDp3S2oARZdD4dvi6tqjxLosbHx5WfhvZ+MF9QMxPhpWgx+Th2vPYsWyW6+zmTYklTrswK
fXWjgdaq+NN8KWHSvTZYp5dTL9YlwapRrbwKXCx1Ii4UEMqNx98dBRTZ+xLypsPMiwwp+1VZu5/S
HUMSrpClK0txD+4+j+6V3hOCG0UnyzC6I3/xISqeBdXEyqPxsCyTwgOh5HEnYem2PL8upxt83uF/
jDQHdtLzmF9Pk6i2DDQC7sBkc8nuOsT1z0i8+wpl/3I8Gy8eKyUG3HJqrxhoL0p3vbnG/Pwdi7mG
utozleUIhjagrQf+zZXtKlfMYbrjmh84p9V9lzv5nEkw/cZCoJ2cbrxYXKUQtjC3PIsW7VPwsrQ5
/jpX3Muvxsu9CZfUdWJqdsbKwJu8rOi2nt2mSYsVrZsJZqboyfQI4JtKlsq12fG+A/4GNXBRl9VK
YiDRJ5zvMx93e6DoQfz04E4WsVAfxz7J5S13hf5g72BZwLeZrVTLBGonLlxN4BfwTF2aidUF+UJM
/ZbK6OoKE6ndByDiPQEM0eDv0R2hDKL1K5JwkzjosxApEp4O3nIFzmwJqKNBhQr93tWywSrHKaK6
33V6u7U7pWIliGEsFDHj1tuK114q8CJOK/EizzcCIB0ELzGMYfg2vnWdzaE3lMct+xyPoa6OH1Tm
Pl2HzR7Zi5qeNY3Pi07hw9zCxCnlwJ5iJhDq7WkdDz/W+KaMR3yPgUFTTaftort0wy0GIJTJ/dlN
E9o4OjSqiLy/8UxYoKUkD1LYEyXVu0HJqhfXNWNQrh9WEwaIUeQM/PeEvt75nPpBd9XUYDvQTg/K
P8hkSNlf/PKYrQ8KMd5QCnVqHkvG56sOqt5cbA3ktgC0ypFkjiDsSjQx8c129yvBN+S+epXRAu1G
mwQh4wois1lmE+fi/qtI4XA1SZkoISvxhOr5RP28JAvbFQR2otpjKPtPqHxKfeXuK+tSBg0ucrkz
VM6/+QZf5dzEoNr5QhDcEibwGM+86sXVm1DI2NHCLc/58krWuFR3WuGwZf3OQpbIkPmbGXCqUmqu
fPkwyfAyVk9KPu7k6Urk2Lcv+uHhj2w21TtKNiVEyzZ4ve3jMwnwJHtu8zOmfOoaXS7auym+9Ai4
+UsqlEAd92wgwBlA3cVCKyb7lGHM7+um06pxwd4Qi0HaN4Lsri7VVuzu8K6KSYZFKEgt/c26+oT6
2O+ioltXjXcvj+6c+0F/jaR12BbaEzDQOj9uBEmRK24Qry/I5ZtZNgJ2XMoyWH59HZQht8sFR1oa
fQzhCL54PBf0u6/bKqqCueqpAqDtBU95+jltMoTnRQ8+m+4lFisF77DXph3t1KB7CdYau0HCM2sr
LuXUFAGgdgrZwkMKExGf8OXD/COb2VqGo3Y+JRZsUndrinvIxBU9UycG9qaelu/hBhBujyvuj+V+
NF3QsPEegnntA//x2T9VmlabAGxRf3mFlEnvip/UQmJaRUWTkW+EMezSgLPeAFPYycejmaxG1E12
2UPVMNnzZ3hLECt0wXKvw9PAKCmNEkH5Y33yjQIejSDo/9guunYeW2O3TwJg0oHvlOZL9XL998+n
oy/LWkfCEfM53Nqeq+CtJImft5bkcapmD/LdGJI6D0XL0fk1ZA3FtLfrp+NbbpZGsBwe061S8Zdi
oXPa8TgICxS+KoPBBt4k/qmXK+Buriq20Ve1p04Sm8XuH/ntsLyHJiXY1VrvfqCBgRy8SlWOmctA
r3vaS/dsGPsw22+GsV1g8xPg/DIkVK4xnU/TSa+vG/Zs4VEzBeF2Ve24wnJIpwBsNMeh40HHsQgO
d6VhqljtcwwqXmD9FuQmmXzEzHmtlLgieZyxn+SUxLQrwhIyJtxfWKdijSeC+tctHKWnwNBwh1qa
1/vrI2TjOr5k7xJzyF36ZjInOr+XJRyQ80CwzyC6lRLen7EyxiDAon/9R+lpkoYLOF8qIVKALyLE
zDU37GMAzfkQ86RxxFnDtePQeevZlXCyOtC/kgK3t7kirgodXVTAlBVJHXGf7h4nSu0sU28zF7aB
pkF8eL++B6hf6oB2b5ysZ2SLSMWzPnf6TVgmzXY0U6ASvwCJ5WlQOer8/UTEYpust4qVWOuIDRmL
dKrX72uKJkURFiHYkRM7KBG0GTJRpOBqOn9inytbw3umFfLobTpj+03LixeBRtcnmkQbRGqaF2Wn
9Nhoe/GpiL93cjfxLO4/JwlT79rKmI18B9jfaxtbY+t9BdSaQ9HwkuXoautbITD6nFuE4sHxZOSM
bvWupQGwMKBfJsmB+P5pIodzrbvIAoypUYtUo1l/OVMxoMBh5/4sIoEnLC0DyBmwv4wEFa1a2W46
GhgMe9kmjiSSSvpIOHLMz6JFYwJ3ox21LTsk/ULbiscmjpOD2YNrFzC+JjPoquftsTAmP4vIXW38
RkXAntDV14tdFTC1sV7DVlnXnyZSK5h/PTkTU7e7RNpi1YPGK2JB1nE4m1uzG+bKx91oudCpboIs
mcs+9okBGMfHwXjRm4OVL4do9uYUAb4zwZiQe+d/CMyz3JhzMJI0/rrjkcNw0hFzziKceIYnAe+Q
oDPiiw6CEZRndlIO8+CWpWmJynMK9SPhwvvhCpc/0nCNP5HQaQsKpxt9o9nHE0p3n5D6c1MAVPrF
kMVOvFP39IyQd9UJTSII4j0+FAoS1AowOfKhzVYhIOXkGfJ97e9mNtx4lFJjeTP2dK3AjsVl4/LL
+KicSrlVhH9xVaWF5E+Qy1PJOmHx74XjODLEMFOmhWY+DqNnZSQWw0bv2EgbYLvAtC695DoLpzXO
2RfuoW8ZwDF6ld4PWmcnOTwzlalzdklpMtagxf4558tyyXU7gLoOj7pgdNuguPQ5arnp5X50iH+l
7FzFZbyDagZzMvivmFY/LPhxcfrVu12FWE/TaZvhJQJTwHFulSfH+qGNKh0PLYRJk9wTk5Fb886N
auMwvs4bwkNsExx1TALpuf1CQm2Sn/zFKVc/VkA7tZQw2dbyB3CNe++JdtjB2BEsnAp15k+PYJNu
IGcnORMipJEYg5yuvDAGCX7ygVV5aNCBWP9QI/R1wwCOVeLNKqy6GBTpSAy21o+Rm9eonnsNUP26
ZznYwNjsqobSZY1cvpkazlk2wG6f/rCS+x9wng4X2iCcKhO4lOb6RJ2m3jIOdgZl3nvK486yUgst
Zhqa/VyLCBEaxtpXcsjQzGgGeKhrqMspSHRVgOW0BeKQ6QXl+6k+cDbhT4oXGxeX8gsyk/MdsH1j
oIpMt+HCc++AA8N+2QEySHipPd3EB5xr84eF3r/sh3HEGSvENwP57BIKeil7AdhKIsVBPXJFpgrq
dHyU/vXefpeDBe7vdy0krobNBA1dgFapwGTP+FOwCTe0xCqQCQqWAo2A9L4pC5Vi3vuXAYd5J48W
ks1xPg/mZIDtHhL2cN7Ws6xhSq9ssYC8akPULKhPLjDVEouT+0dFCFY+t38nT2P7GGKI7A2DL3zL
OtOuIlziRAhuSS7WCBjQSy/DxAFONMv6BjluBTZ7o5pCqFvR/A+PZF9an7O9ZwZxRuQ8j7jHvmt4
xoDvfz5zbR9OUK/y93B8fg/fneSY2UncIrM/nh4V3SUoBaTLIGAAgMMktAWpeskpNF+sPvQ262uL
qf0zAh0V6mKJGdRfFbDkBy/ywbFC3TcpTNqXsCxuxSXAEVcUxhj17gjtpPr42+pMWWoXXawNxhLH
9cAxHQjfn24ME21hSKbhkdnr9I0dt66r/7SG+Tks1FxQjS9kpxIXfnugpbdlnogl8d5vqenXGgMu
fLCo/zMV8N7buFO7m/6fwTqAsyDCga1wAKFiaLbVAgxbbqavFDW0XNL6Y4/eSrbApgCRF0xRlJkH
kIby19a01UDt3k7X9lcJNSjCQafp9l9sGHqSIx35m2WXgjIi9EbMnxlUctZWapX1FafFgaRJE6w2
gHu8pdGDXkfM20d3CWq7+ieaBpeixncqPyjiV9rJ/+a3UgMDE6t2L0DaCXy678P4I4WdJwrXUYIU
E7H7KORl31TpRcWJZIWP5BSILrJMOlXgLM5VcHWdSN6Z9S6l84hIJBWkX2ZyqzS5ICRlOmJazXCR
Ry+BWaxnix3/yIQrzWRQ1Cxq9fxtXnVE0HUzDN2oDslmGdRVYoJlLeg98UCaKhmqYaGCOk8jDKkh
s72r49vrkX1Vb0Xp4ef/5dVGTPle0yksLEdiRWHpZk1myh57+gWtMAu06aJwUQF2VDXGNGBuB4lA
JjxI5uWYSdIgjZuekJiOViliAWaj+X8GAna/FFxY4VgABlTqcpYQ7fbtAVBsMJEruJpsF/o8ina2
7Nf/xa/0LNhvgnDsdywaYHtSDHgTdeCmIxAIJak3NaYU1nNdtqoy460jfhY8gJBx/QZJXqHPYcEF
O/g1JOOGphavBm6pZh5+VrbezwarBnnX0pz++McKiHyka0+q7Qt3lfUUikxNuNI2iwUmH4Bn1tnM
FzwpTYt/R7cxceHaBLOZYjP8uOvBtXaU0imEtstzq67MySIawitxteMt50yKqHNtgSyQGdiENRa1
Dx3cArjpkJpEFCq3MXC7t5L9ZvvyeuMjttsxsI9LErfBbaakVXns+SzHvTiTwRS1Q9I4NlV4jB+O
vJx14A+97Z3t+XR5XgQv32EjeSgzgspWV1MRILOIUkK65kGKpxTbRuOxA6g+g3JJn6XkNaacuksi
C/lv2V937HvjE87+UX3hRTdVc8eMGkpxaVvou4cj+3nxdCg1VsfoN94dKorScS+I1CV7YY6fF9JC
s/OYRUwAvt3Byqtl0j+odHuHf2cKLx/R403aAvY5aB+55OKl33nm6/+i3AuEMQZb00EZpBcHyPUn
adLEdaiue7m0u10YNQEqdARqWapXK9YE30PRXZ0jh16HjOnvXe1dW+dW31ReFbiibJsXI1fAtner
xEPh2fTrOQjc7/s63jNkrYsbiyFV/8BuQrMaeKV1pLNXzO+Vk2tAlv6wIf5TMYCSvRjQT45O8cZS
PkkWwpy8rBtZBMYnLh3yBZWd9+dI+bHhnzDj7V41BZuTxgVmNktZanFzD6gSkrYqoui+peScDwwd
+CvEcMnNaUalFLRV1uODZy1uh4fJVL6djyBC3J3/4ts/Z2PceKfIMwnGQ5OEM2bU7EVd/S2JCVo0
yjRnaddXwzrpCzHn8Yx0jcanzKBP0bMAH+6Hu969vZQf5ZVXocl3jsN1N0ttxDHjAmOjLw7WV3P6
fmN4iMQoSKI6/WMlLWgMpfilQzTDoXXxwhZfvBaOvpxhT3HMuLUk57XJblLE5ezcpIvTYX0WFsej
ECT74ZBbh+9qILeg2WitQml4CjynJBUAO7bjByQGC3sI/FZgUGV0/rSiy/9msWEGOUrrzmwUXf50
xiUKWRYjvujx0ZPHcjLqC0UDqvLYnxA9hTZhwLLYRFlMmrbYw9/M6lgrtAuZCK1V4sga3lzBsZW2
WrMx6V2FHuBXWJ9AX68dzU8ObKbRcS505kaNI6X6wc1g9Pne4LILa1iDO2DDhyG+xGnticTBsD3n
tz5lX2kKxnZ7v9qMY4z76wJrN5uAUnwGY4R3skH3Mab3YtoG28XHZS2hKnznkdyDS72uHOmM/Ul+
nt0wYx+FlBF3NNDamjZQGY0Q64a3DPVpNhaI4+Mq0kSopcm0+D9tnPWIVh6vMZyzk22trz4eDiDp
aTZmJtuNBuC54jXkKu0jeyf7y8hZKRyC94WbcBIGfjdReYBdBq2DA6dKSGZo+b3Y2c+KRBX4JV7e
OXlWzfLXMs6wElMAizMt8uaSeHQfuY1Q5oac7NpMlj2bdiuV9Lhl7Go5ohyA2/oKC1FHTnyy6A6q
6mlgBa0VVqxFwZiQ8eb/lIpBycXRYrvdBJsNUcLqAkj02GPMlXYpAVWTsc6eWcZsapZJ1I+RAnHk
PV27kmMi17S7vzgCS3gHag4CoXN8TqilKkBxymIGGr6TGeZfChONpcCpZZUbgtwiwxlqthI4LRPa
PghkUO+G9QKnc0V+HF3TAvD/ZSY06N2LUXKC2NWaTqp0W93YghFyqwrwfHGgq3mZbvJKKaJBTy38
VGQhtb1Thdnh6TRE9lRZ+CSpajjATw6C0HeoVH2BJg3RHepTvgoKNNzM92PSSBk0jkq2pODNsr8n
Ci1ovdV463y/EUBx4MdTWnlV5YAxpufJCi/ru5P2i6BywtsjJoJJ/UDLJSGHpDqpgKRtsGgrmcoN
AlrM49Hw7+oPsfJaxbpALHcgHhGw8ryvfTa18Jk0qWt6eAaL3ePWkj3/lLOMCSM8RJLOoL3RE6rz
tuyuvmrxET9K7SPyHRw/I1fRnJ/UdZfYIHElFiVoJGDlqh/sguYvXKMyOGQrxiHFUZPmMZXeubQt
nVe9tpw6EYTrEPkm5Py3eZDfGZwYreOjXjr77X0EOjhrVbyAbdlrG1A6IQnqZUGb9toIFnIAxabV
qXWpFEc6tMJJuuW8HWa2cvKi8Au/ObtvfpFYWOwIVw0scVmbgwMIYG/aMShAkII1IzSYG71/giqW
eSh0RZUlzQk83P1tooVB5OYEjyy6d92g849kB0/NLJLkwunbxGxMxgTfu15MW2Z9A2FepnmKQXNm
/4raZzzMoSofPwrTDSJFUwowrGDTqUN++FVv5S7PCsVwerLPFwh51z1MvuojxTDJ7UE2i7cGaZ4r
n4HtVQccjYT+lF9a5Gbrudu1Qsyfci+P0aHQnV07UHWY87miRZkC3rPXmR+cIwkhuDaracJz8K8a
yebL9vuYQpUDMv+L3jG7SycyPyQ1vk+2hceeIrqxCPvxQ9hQ1ZPG3bwPRq8soVf/rEKGF5WmRXiA
rmH2bdN8qd1XSLoX0LpWZkLLIVrHUt+oVq8bDFFSopUaX28X523nMnHZjDADnlKsQE38/yvqrN0o
tDIU7NEzuK4bTg3RyzJPVuOyTnNnzYz3XU8pls434j9KICChim/58aEY94+EY+fRiFZCReOfYMWt
2d/dHrzV4+fQ7kFhzVZi3A8IcsszrCeruRb6Renc6b/cxlWpAvHQx/LAtYc2ajYeMNlhGEtwxJZ6
LmIupfeeZh2Zd8TPG3Qx6NXnKovxW3txnsW3wnfPwbb7qBzsrWzTyyVrKbEjTbySrUkCY6cC9IbB
/rcgEMN/qWIpOQypDZ6T/HjNc/5ncejoePMNj5EUci0wIVtS69I57gBi7llfLBP9Id7OIVfhk/NV
sRiY3nJSTKyad9SPofczyhwhX1xzLgnU3Chtd1q5tfw+Jo5nKCyYbt7ZpEB/P90RGSFZAAcJzpPa
LyC8Kbsck+Ualm7lpY2ZOZyzLAQBqir4SuCa1zHHxkOvDIETLdqxN0gsDtSHvYbBAxuluNkH07g5
2jqVpYkF67GjDkSqJLEvux/OoXVv2zbqNy5o9EAZzU1fU4eqrpc6QqwxcuB0Mvxism0kpsgD9oLN
wZflkAu0Ly1QSO+1Z3vFkezecTmUUsyJv9QmpEssTVCVnjMIBUZoh7eYjKuWFBEv10DvJwj1XOx1
1ZIj6rHUahwVzzZGkKNA2kpou7hV0yaFVlp5kFZ7wLfZZzg1QZtIHkDAl4TZ/lBsht/8lkNuRCmX
lLMg5PU86Vx9IjoZjbyF5MbA7Cl0yrysxAIdDNCrZCmVyAvv7GFvoZKLyfUKm0ngfzeNFEeu1aDZ
aS0PJBNY1ZujdVp+aK/PnSkpuc0TiPUQ1jIJDEtdAM/yx19/l8vjJf122x2QOJC7aRCxhjmjtiFZ
XIk3H8I/QlDu/W4r5TkoGTwCxe8tGQZ8fnMRJN4SRCyOSJy9Lw2BKa4GUmpGSm6kNXc6331p9jPz
2iHJ2IsVpNxzYqNRB/AJ5kCNrkJu6T1mWywcE66qWoQeSGkkuOR9DB3t+5vK+Wr5C2Cohel+S3IV
IknL5yYh8o6oy3Iv6wsruZ5UUSJIkTraX7KNFw6ngxHoUhXfDp/DpweANE/HrwPBjzXoLRG+LjwN
lYiIrFjDujjPULtU3JIduVXfFXs+teI8UrknXo8DudQ5SSvffPl24/TT1/IHr3txaVDdZ17URJXO
tfXGMfGBjTm2KkXCoQEC9PdyS8zmuNAITmjMEy2vOAtj/vLyPMVyKdH+5wmPAVdS1MuEKaE/PmTx
dZX7DfqB8XLw84oZdX/1PROrni/scr7DpfiPC3jhYVwrlvtn2QjTPaDbfxvslpTLziw+Po1OONs5
qpIOmEEnYQQVvsLj/vcBfvlIf1pYPdBzqy9uksZ/3t2hxCU7NbI9JFYRSSn5ALWQffAG5zPIF8vE
g/Me76j2t4Fd+KHVxZwRsxyzbsjkQFKsuz5jyNU9r6Fxg/CjquDg9C1Xnbe8MkTGX9laKY/0MJ1Z
DsyvibGo0j7PI+RI4tkqWxnnBrVjR5Yem08bNkrJzUAP7D5M1t9d6Nx4cSy6nBGFaEB3LxNW9GY1
CN85TZrNQ3AAjaL7Soxjt8O3JxAVCEnUqwj3E+JFqctM3Ma5K68YQAtrwHBS8OupqQK7JOdSMDMY
UJ88iqPQk18OLWayo+m16OA7Ut+GeDuRRIREuc8lGY7zSmWats53ud9D3nIDcpr3rQr4Q75QBoVD
lYuncSCPbwkUarFL7A3Ths0DczYmh3U3+aHUddKFXcYs1CZ9wShhhRJ4GBDj28pppXwLH4q9pyd1
J3A6p/QWIOsh/3bYH5fhwbNjeW0uLNIK24F6+yAD5MRMJ0qm+QJmQhVDVFhx0U8ijxYjuFxpC/dg
Xb4av6BKA6l3AzmaGr2rnJ+oGcwsaexxwW9IRVWxj4R2dOoA4xSwLyNZ1ccazLyERVKK27cwjVmF
zHqUlTlZWGfbTobIZWLTdgcpIkYeHRCQ7ZEYrbMu6RvUZ8qXbN+mCJBi75N5LuIYzVN8MhQhfSx1
aaK/GS5Q+jEFAdfL8nqhmgm2uBYu3+i/utZcsKd8ZHs6Au/EWY56B7hKUPKATrxR6+jAyhwcOUK4
h7s9tiyuwpopRggHSLLVbg5cEY0+djkYRgX8CqRCBVroYXNXilDz3nWRM03yoCuK4Obbyhr7Ki0P
QsuCX47uS+8QisFTeZua4Dgsd3d/K5NG/mJ2zWWx59Wc/QWPHqhm4YTcfW3ToTd85UXrAZXEr7yl
eS2TzEXC1dD8x8l5c53PV8n99NZAuSLZW332zItegl/oSg0b47mTyNb49XJfRwVm/UWLrzEVweJe
XAeLjK4qR9MKsB4mCVPwsy01eHBuHqwrNw2NHJk1HKtezig+b4C71JDQ1cOBSpW16ioes68+YONG
6HF32F5PMpWadsuzT8kwIpD/ze9sHyjYi2RfAVfpK3o/QIh+YpOrp1CM6zVKjs/5X7MW/UJL0DWs
6IUUAYOxw6kqdvD1izwwqR59XDrSi1aKxEBr+R7LCTXqWKPSiv4JwpI4seXhMbp3rNkXNIZfc8E2
8Tt5WenDAQNvf9EEdLtN0j+EUiiEN7VYJXVSVhxSl/4daiaKeaNbYsdJt5yiOtWu+LdF6aWQi/i1
e5HJrZxyAOkW26mTm4OhtfylO5Id0hwLDPKORQSrZ50O38mgt/Ny80C4lCgIeTCOA93Eo01oe70J
C83HLH4KfXMq91aFFISGSP/cPtZ6Ga5JJWqG3a0CIOje6dTZNAciDFwT8IFz7il4dnn6zL4hNlt3
TKQnw6Xce794v3AcTP4VGQUCXczvbB2pkLTsCS8L/oim+vHvkUyujh9nB4Y/jEjmi/H41mrGVb9T
U9AQOFo7xtHCtmf1DfH3QBwoKC2DBPZZ8uh0J0B/x9Elnf+eSLcr1XCIgiar7UNY2yBe2hkPheTI
JTEsVfJ690XxKtcUr+jjBhLDQLJ6QvKXzO0OFmbxfeGTBMpquFgCo8TiLDmhEolWHQ3gaJosqN1w
sbwSMLtgDK6AC5MpS/f1k31E3jllg4EsrOzJv2HZoBqknoJmQyn7Q0Sck13/lwXTJ7YM5iokdiK3
27M28kkZIsWFzvbGqMfRTg0w+pqIJkMVJSoIKEXcKWQekDOd0/HxIXHyqasow2ndLpNMvyoVdETX
ylywqwAPxZ6l/y/pRc72e/cfvnjiX8fzDY53aRvMjykqcbrUbmkNctV9HIR+/HG6mqRjMddH8OUr
VBgI7yF4/WZUe6JjoyZ+51OspGdi3ar49v8BU4pt2L746NfCTag4Y4zZ04aaKgRP7OyMPGZAhAvv
5JEUkaQZnfIOy9gGAmzPVK4JYaOJsBi5eeaG0r5wm0g+So9mL/sAfxu66zI500ZJnhBkzuyyqcX5
k8+DL0BzEg+BT+ktjBXeLfcxvjuZ2yzXPEOwM97tlf5nvQJyLirSbhULa4k9BmbbJ7JtqzSOLfgI
tdMhkaRvRan9fTvC5bIYvgXwACmmIIgoE8J1yngu4HCprN0n12FYXVhiL2DXoGW2jRwEQw9pOML+
AJ5UIQGfLjDVQnKS6vxjE2/5PYgwAFZh6SK9wUaMbA3e+KsubnEfhSnukeyaE71FK4B79cOPFbmC
DQL+QMoTLVkdwKXh9RNdedLb1wDVlQ+arw9sa8LO/SbVSMdPtLMlWnErgRB79aBBQZzaRuajFP33
natmvLuFE+pu+ZZc7y61WnI9Rr3RSHTYV+lwBMLukJKM8GnG93HrgD6aGVO3Yqt2MPniO/t4D0Ur
joc17nqwgpVfNUOrRwrZDeCHWN0ZEQXLfCZKGT9kxnG/4iJ94dEJ88XwtvY9w+oJLXaTuiPttaKT
ikxOLxsxnES2sFjgv8OJhqaIfnPNrRlhjRBghA7SBUd2G8KXYOaWwNXcxdRuJd/+eOaT7D4u+CLG
X4LaVzAqPflW5FRnwliC/R3YAgctRcQjRq06t038qGqN+1wzY3kQo1ex8zEaav7e7Tn18tCl0rzv
C+jOOZQ29KQ53j+ObpJJd67zSjLziV++sJa7wGyzCw1KwwruTfi3LrtBEpKfqvD5YAsjV0Kx2tA0
jbR9ZyK8DGXRfHYHPEazHILSHZb/g+k0LsnAcoUpr+UXsKhvCxyzmae1mIYvgKiT4m84J+3Fk4Ib
TdjzzdD+T8rdQvjsBkynr+SNz4VPWFhOjbW9h10SGDFLFkx1PtiqI8AlKAvhVFZJwab/C/bP/ZGp
gpaJRXFzWXT2nkFe7w7IO/mzSF/idMUbOGytjvgK2GfvGsLWBR40s/EDEiq/zOqtemEc3PutRhzg
NT4beOl+UsVnrSCEOsKD/frTs8aCd5UV26cemuXx+gnMfGF9DfvAXWyGNK/+8OysQ+y9RvRe8bqr
sPOkmLEfuYBb6Nk+Cp57cLpQX7ipSUW9CBr/B7TVpmogKsxXeH1jrECAxhlesD8QxV7gSVySYja9
foLqoGz+8L4900OBs2cS1uHn7EU4k5Sgtx+pdha6OmPySilmtd6lJIIlb6SZC1bc2OXLpk4Dzmh1
yQ51r2bZBQOGryvj/DPM+z9ZVyDAXPcLcQjjIJZv+6qsQIvx1/6Y/pk1CwOCwpBmE6+FvQLvd9H4
NW+hHuZZUE1mQQkV2EsBAYUkShwsUcr9NBcb2SG8ha7G/V23mTxm3ClE00bd0qAlTH+L7NGMFr7m
1Z2ZnfuydS87RIHUmrN2grj90Z3MTROuZtuFUA37pigL3ZsQMfcljT11HP9gRtzSuPXgROhqYJfx
k30OdO4O8PxPIKluAaCOdsV5BIzELYD86ejQOudxjo6ih1SVUxv2BbImDB4l78g0zNp2wMV/7DCJ
7Dfwp+GfS/mLVd3WzqkRFRvOjMOl5Bz3MvqR50SsFna6qXfdvYnZndUpCIsHfmwqywttxvoxsKRA
+jiGzFLTyPUi2JHAPbiVYWIBwuaG7hqUZnWAiLqseAQsjSIAsk824Z9CNA6eZ1vulukM+fF5KyHA
0SCOTV7qX5iUTJcwB6xi4zKEGObhEQBnES9hBcmqCTeb/SpoyGLZrG90ajyw7iZyAw+AjWQnZ8o7
adtnAE9WHCZHvBMXpJwPp7WZFYtL+yNQr2q/YXNXmhPtrRAuqx57fVxuxKhCwngFx+YHnk4ESc1f
QyYHCHW4ihUosFX9UmZgyhwc+xXb0ollxNpiGb2Q/AiBvoYwwRZExS30HkD49ujKhqiIZbzXLoDc
gX5zd2Bm4A+UTCzbNTP0E8log+yitkSAO8xSZ1v85KGPZRH6wk/TeQyVc7vzC37Z1njcZJKJgY6f
TlmVovvOIh0GrBWGepu3obF5Hd1kN6lIU0ykdOP3sRYlp8gUcWTEYiXUQQNuhlvwjMl51OjzhH1a
8ClBsrhnf8tDEIN45dt7ff2zv+BtoDNqyhZkBlAU9q4j0JD8QBmUD8ChOL/9MBn4xJF3zz6cC2SR
C0lAC91bcSwiD+qv7BLke9zx6El6MdUQlIv7/AqtJYE6GoOkkheTIMVBWnLdJWigdEr0HEpuPPp0
rR5FjZjlPpddBgnnNZ8S6onCeKFGKZMXwPpxN13hC/K4Wl0BkM4i/tkeEw8RnaBtvLjdeE6kgG2Q
ZpWQiCJn5jZI79T1C1gbc8XaQ7uJaXFxY7nkxX23XoAzjD2EmvS5s3kRfmFunjsc04YNjjfxnjmU
9lPnhNlNWUG/FvR5cJbQW0/rYem8E12btuqvbT0PtYWetAYW44a2BkocAjVaJ1x5s9AGOZFz/klA
WqWQ/keZWQjAXrKNfg283S52MN5Z4UOcP/TenijjKNE4zZfYFYb3d6IcDGFBkjzoq1u5/HWQdCpn
WQDEVwr6iHk3W/mTZIdWZuN55mIKzL5navfjVS6z5Iob0v3t+5d9tXUsP96ra1EgPzNXC5HXXBHR
LV2jMDpbB//Yk52/4Noopo63wesxjR5d3T8Y/18mL09v7fuJS78dyixY81+TEtSpnWhXpHUYaVx0
RsCqsDKapEBircUdB5ibBe0mE/z7Rr1eMulAwepAUpqortNp44GKI7urapQ/rBVBduXL+U/wI+44
YDii3h76ryyZ+a3cEmJOyE3CPgsQFirPbG+6xyBNnOflwTpEJjNwiWkmABFZr79RwdhQ6VQIjJZ8
M9at51EmL3v+ScbAoDv7wSXUHVaaY0f4280D3KPqH7rSkd5uAj4ltRqx4hw+Q7bnnaTdBifF8jov
OtxirdlRHN8lK+aEuujxEiW2G+mIC+yNKc+rhriSRDyPqREIQbi8uFBQ0qh2XxnzJpSYt9g4c8bx
8I1ZyginmeSI8hcjVBnS1wbaNCxikeEs/cFCRvUQ6q4+h1ywu2FoPLq+G0hnwJCZ+hfialOyFrot
tHtsy9pt2otOPkRjTSJKIknmsvba5DoEzK9jJRZv2My7XWMgTVHRzl6mYfR11BCWis4dNg/6THIw
9Xv1PB9LClxmUAQcL35Fq8IX6TQghIb+QZX1h95td6+GDRXhxl92aKpLtP7o5/uLbIzGGYAyPYAs
X7hL8aQ1y7Kd+VNzn0Ma2k+5VlSg05CvqGfR07eMQIxRsfaaJtsSG8WRd+QOIXwfXouWP5F3pP7q
OPz5A/0e6WkGEhMltOkER7/O9olDyNXbyb025Qtl+CXmiXnCbaSOLu9xZpr/zpTTPKMSMRQUERod
a18aMl+984Xr1/UbLPyLLnpwEUFbd/bV+BJ4VEudJUPhJ2RxfBoxMqpu/H3KVLtUIURST0036N68
CL5oJWZKxDNR/QLr/0Vkp0A1WRkrgtn830JkGm2MPmPI9XEiNfV/mPiGxU/OKHkBXybyocWjaVT2
inoZloTQNvJP5gahuZJ6jPUA261ZhR+oblmuIFC4PsD/Zdjysz/q/UHbUf3RpfjKC0LdxkM3/sD5
TbxBM7oSTrQ3o4Dn6nxfe1shJ+VlARkd1RnHTe5q3Zu4ivDF+Ii08BsGL/8nLHZrxDmki95Amwx/
8jDuAs2hLa8E1h1j6L9qUfGMP8gTJ7KdCkoiD8028Go15Pu56tgBFDBlKfH8yW1KSvJwLjInEXhD
Fxdt3NJXYl1PLITR9eDfNUWoNj9xQ4Cn22KelZr6XB2vQOK9JvyLW2vdxF3jTz06j4n9tpcZaWg4
kChQqYBm/9rSXrAH56KqAqJj17pmE13MrwtNPOQj7Y5RH6id1XoCj06ANUJTZT3ebnf4Z97VHAcZ
tzomDg7wcb288OsZUlIryNr0SksaE6ZhC99eV6hlcMEM7fe8uUzf2c5VKeWCDMymLM8ZZJh7hqzp
T7bTyHOOfUQYgTxcT42ffYtKCKGuC5zZi9NiJl1y6O4uEUUzqATFlSbHDKpdkgAIjj5RPBOGHcJG
XS153XtS+Vb11wBYkeJGFTXVDVzZd0ogvKdciLdiizauvzD2IU9YCj07I/9hvTHMgvXI16Cjb0er
K68zJTb3D6adAB8CZ/eiRYSoFhcFs38tXBMDKCQuWxXtHBJAj2w3czwUA+zPKlLf1YQgqKriyf/x
VepcxOSSOL0Jpwo3SLTrtXf2rfJlHVPda5a2Ohk+ybi/F6JrwFcApwXiNjM/0UyRSX5E0DuQuE6B
4rHVQtrW3byeGYE656a4fFV503mmVkQ/XdT4b+tvP0j7lQiyISlGcNT5klJxGX7bB0JFRZxO5tWa
IxqOHlv404XImPdwxH81Mk9Kq8guOgglOwUm63kEpzSA4x/f0GGnzqIykSzXVBc2Dt1NDHVsGqtg
EUJ2fnShaKxTrM2NBHpJuxupK50XRUOroCBy3s+hjbPo8btv2oJNbVxRQlOrKh5Wyu4RDHWrQwgZ
R+Jlx2TPARpq4kx6j8TkSbU7ryPDNi9F9GJtLoJnBwoW54Rp+RZr7uC4NMAngQGr8RZUVTDIJ2Au
H1qES8Y0j4bjtmGPpipy3JREsOAlbU1alDtkeZaSIj13QyJ1pwfCVPauPPdsT7NKNOOCAaPjEglb
6S8WkGCJUwMQhoxNESLh5c7+WrRNiSeiHSMzOKEkeFLPkNguknMO2z67qFei8iEhH5iRUonKcL+e
A1T56neuIuc2TZL9Zn/LjE2O2l3JIVM74TEdV98p8c0fUHHub9NkSIXcadz3roYEPfANA1jjMok9
SbZ2OsYBfRS52UvA1JT9bHE4Ctla7W4klBgrzJkzluM1o8O07JHsuhYqOZtjXRyi1mwzxfYsvjSD
qwipomojrEJSAuihHVsfOIg3tlu6tVABnoP4Ee5jObPkKyjYz0neuOvXJjYrPyQ/SthfpqKqdIJq
S5DL8TnKXM/NlouzXqKNSToUwxryRBVBZuwc3banpvgqrbdRc2AbY2Ep/LGfiFnTBUnNUU22/O1v
K79r6KiYbwM6tGhjGVg9aov1G/QIcjnms/cMx0VrdqqbLizXryXpREM+3UaOyHeVwZvntynR/hgI
zYQngqcpPvu7iB1H1orzzDpPlnp0ULsY5KwnBYru18xUvjrvlTRUtACOA28gFw+J3/tOJHWglbaT
tgk4L7jzCi9JuuEsaAlAxeBpBPQniUHs6vSIzLaCtCc6E4vHKkrFUnYf6oQPCfYzIvrlGtGcxyMk
G+Dx0cwnwqC8MBMDi0p2PjpI04Nuj4Y4K4smwFsSBBZoQe4tE6Ii4Tfjq87I13QnaJmQtYXI7rGb
wwggNN+x7rLmXdK4W2BEh9sBWMmMZXf9IweBITjrgJyOw8s4Du1WAyRqraaJ4fU7SvVCzVq16sy0
tHjpms4nCbRcAOWSkJLvkCsfsKg8afCtZXur3tZ/BZOfIGuCv4H8fgWWbWBU/ARGsFbzMdcEUue0
xSSolsB/v0fZ1HFbq6OHeUGN/i8qkrQTe0NOY8FfqixUtCXm6CcJ4lsTRNEyTHzMxOAU07ss2hx0
CBi+R/CWuXxi5rxo1X4Pfq3+CG7BWiEfbH2Vky/i26NGt5x20Qpu9hGGRnjJLb7rnhjjSubLJki4
S+eEnsnf7hrBCIxL9jTUZzyt671IvUCzu7GFo5XjynNUA4FwKotft61+UC3FnX4buPQbPXQO6RuR
AJoePOpgQoDtiUyoiejbyvpKCxu4NDQFdtnTBwVrG5nE+ymiAp0Jv3WWDJwJ2YDaD89ELQdmBYp5
IJQSMUuVGHNhRZXt/TagPJutfvQfrazTnuZ3xMiio3Vq5KFEDk/G7kwUC7MU5CUFVIHh4lC+uleR
fZ0JMnWKAAEB/l1JPuBYdh449MoEu2DDDM9uOEg5ZmuonO1nUEZA24bseWLbd7vRySgKI8s85TQV
bUiEiaYJPOqPmir46yfP02yk6k6/2KGYDGRPfqS3/62XjEedLOXNgGBiK7IV7PAie9VES+vfx511
DgFP5mtoYkWUx3iwlltbAJBxK908DoEDLigZ1wpmTqybyrTUp4HQRnwmXIO4gobSVkvLobxkrOP2
TXEEGVJkzHvt+cXlVPmAC9hoqAQLY+0EbFU+9F/37r0zPIOk+YP1tZIgdZ4D7E3gcs1fjZZoECtC
0VeBd+7XIJVT40H0+RlMO1hSc1h9k8mDlPTfiYQWv5uWgdlLx/kXE1a7anmHndBlKMOKLkfPxB6Z
gY231PMdn/zPCVMKFwKzwgq8p+TZmjLUL7vZCsTNEpn8pkUnx8QeRfP5yIFy0JpBW4UdCDS7tf7z
9VELfRcLDe5/u6Lz/qPpmNBN2HzDp6tPVQd8kba/Z5k8u5WI0gF6cwtSbByaYiwadwpUUjA7ulnA
HTNXA6Jo0aMq3xAockZozzZlHMWjv5rWh8qqX8Z6bNakYfg3dJU4E88wdUUFAk2a0ZWIPnGwoNKu
1W4nnSpMYPWnn6pUmzhMddJ9fdvn+IUXC6STmyHWxpjSg9xRUxbwGqkUr25BMhWpUPeYl8re2jo7
fcH50uZsYlKE3PuXweEWWG99a7RpbV4IPc3X9dpv4C5U8+JitY5bYk5ewVjisHc1wCTkrB2Aatub
q70ppR0CnFXGcMV3WM6RAX4kpC1VP1YnFj7YuuxaLQDZlZfwMCJtDby8V+6jSiFlPv7KsGX8zQh3
SgcoFazUQrft0p8KEu4QdN0SzoQG7g5kxYWwWnLApafitiveRR2tBOMwNBwTWfnjVJlsYysFJER3
tJlXvDpFY4OVICIDu7aZovI5nq63QfFop44Dp5sQWVzS7TvJCnMtFl/9Ea6VMUp9vd/yPV3LlBMJ
REDQULb/8G/bU5ac7haFOq0QyTvDaZ8GIfrpD0t1E2bH+U6xsKMRCls9iSD0KX3y8ltQRHO10Mxq
K6W7KiSagfBQoaAmCz2gdKNyXiXKPuwttNvop5K6zMlHHvyM1yE/C21axXZyPbAflyHtHF+DaHaF
JGvcP7cxPqh0WnBTcV1Nsbn/v87g+9PEtZoIR/bcsvcGsLRHtcA++E6gDWXLQopqLcGBmAoAmVvj
/+zNl//6HI0IdcLAZi4vn4ksU4cpk72/KVFXtr+cVPN1E9PYgcBPkbUhmTOgejVMEhbLozsRQWZf
vYnPQFwuUVkLIY1Iu6/nS1VXbSckzNvOCGwHEBph6qFfLxyA0ChWQHBH0EepRTVqqmh4q+zPeQPK
rWyhNjQN/WJ+yzr0L9nyQC5TrnQNFph0C1NTkmcZwKukuk6QnP2ge4eURRhSDxXnPxEIQ5gGZqMy
l+X/eXcpw6wDEH+fTESARb0jevDdOBa+63gm1tK5ee0TEb7x/Vqebt1YCV0cfxUuCEVhgh0Zlms/
Ih/Ny2xfXrQ04P4Kp8Y3NBbZ3g+nzTnGT1mAimtniN+J7/OYVWw+oJhzN2oGkxoDI0qUXsOrHDNj
7Ni/Hk940nbgeF6e1bhsDq9U/bQiogl57EpWFyaDUthfUERYvPoci9lAIiywNvEIaTu4oCaSFC/o
VI5UxOyjTAqAI/b42jNmIIsPMkYH0EytLLkcBnq87VDr7PKENWqaU2a2Cgg4M+gxkRvDs7AUVLo3
x+CqcTWfgTRJJi+FO6OU3liuTKGXfFzPEj/RtnWTFhtr5jQdqn4TdkV4B1bED5A9u7r5PhsuC0M/
+8fzHjOFz6bXc+wjF3lWrR3QbdRirNkcMh0RdXKjpFYZK+3j/Wv8Veao9Y7EDl2aXjCLYF4LPgif
gxw7MW+PAbfq+/KVQhyKFOseVC49mS1QeA/IC9sepm79MCSZaqNTFm8oBKb3UW/FwWvBQwD3tXdW
dvxyA8eEHcyBtxpXnBqhHNhIJoLu4/tUp23RDAyIay9XzfBcf6C8OGdWdKApi2THlgFBd/meY+4R
3omwwAd2hENfV9U8iPHMj5kuHmzwG47zA/RkOc5Eqq6SBYtL6cfnYOt/YdOQYp/VUw8sODXmw6zQ
6EnvqivSaXsf19Q2KjSnkfFHItbiHHyteF74P9oqiypErNieKtVi9aNJEKvK1VbCQG/2w9khK8sq
/Ayg3Z0aGPWM6Ryc1WBs+aBnezMzgr32GypNdU/7d4e7T1DO6/gNvfQHl8frVPJ1UYJFs6FgmQBz
bDq7OCCU8nJIEVEjOHx2Q79sVk/8/xYzhYW3bjlaVm7CV8uBy2benp9wvPRSogmxkmiVcbIgtTmx
6d/G0RAFxp/uAjpVJxxVfHbdjo3oyiL1JSyWKoQTVMWMuecapVOeE1VdcEka1e97SsJlaoH4fSKF
D5aRB3RBg0Z7medIIi6jibYQ2m49BC6MndD3gPFXe15TTdf9TTykRa5MKl9nuaMBx9+1RuzOLQox
02hlqYOLrVDyoTkP9AopVGok3+qUb4fyuMzTvzF5Kb1ZFekNXrdvg6h/FiDtWqK5of8+6qx6sGim
zHqfKXercrdh7361RkWKZgtS+W5GgMGVHQDf0w+cC+2JCxyEcWvpNU5G2MZodIzJDJ7WhlJTgfeq
rBQ9caTsbycz8tSEvE76B5nL6QSgRfXilfxs+RVqOD3vX5HzJTeYbd9gy9L1BCakOcXeULmxEEaT
2IyXHaOZ9wIDklpQDOoep9IN2rSNT1gf6tOuKoa4ccFPI1S/CGAhXZ12jMo5l0O1+2+xTFZy9MSH
fOcTUJEaib8aP9QurQYTv+s2bF1qE0y1DQy142sWAtf/KygeM5vlO4S9pmsBFXZx9byOsNhgx9vf
ZhcS/aMPOW7jzqgtpF3oSCvXIt9xgsD9kwWAMjYMe+SKA6OuxUAQne2Q/Bvna7lcjLzehUDmt4Mj
t//+EE88t5nQCfWzD926iVjCsSMLFaRVsa37D8f09RsVU37KxNTDElde1VEw5F2ae0jcxBGbzl7e
FDL+qggqLJhL4TJeFw01urlqBbpcXzbyyuej4guNoeDBSGbezCT3V5HSGIKVIwz0M6VuIGOSnVYS
Wa3AFPrkFNeZZWXpDVK5WWvx3sVrlGaxLtpIa9WZ9b5JWDBPe4myoxwPEw49whetRnTPhohwgbQY
4qHU2u7DaGiq24DoKMIfc4Zb3kfosJZ7Ed0UTw8IVuf+zTohH0GGRHgOrpYcByH939jJO9m3w4JR
EeMO3ouAPFwsy7HXiaKybasjafz9KRsEfhmKZUaUv76lL18zatLmv7TC0xaps9dDOxey1+ZZABid
xxKm1u2bn58HXtM0F5U6PA0Io2pI0d4DNbGzcuhlV/R6LhtCJnrO0XhD6l1HNhvsBb1abFhd20Oj
zt8UYzxLfa7dm34XqEMwdsBmVsY1vjoLdbNlIpT+XebAEyIt2Kqo6739UXqYIUl46di27HBhnL66
6yJS/mLZJzg6pqJp2VPUxhZUY/nnDZdBXdS/ydhs9dq92AozRoS1zNXbDBhpjlU3QqEfffAv2uC1
H85et+V6VqO9Ixmb/lm0faeJsegdlz7TonPzqbNEKDtdeXsoP0ag6FOImz3gdCrwhkfiO+4slXBp
xlm0d4ZlIzO0p+2nl6iJbLtXcFUAiplwTkP96+Stf2ZLqg+nnz+bXNRI4eRrWxKiWi3R8sTi6irt
ifActp6YUcO51ERk0ACZ2EvlBZMuLANC6gIOjk1zyZOtAloktCBAdHd7RPkcZldYW61+E+fgR0sv
pCB4aX3TKtQl4QNrS6Rq/naCTfty11Uxe3WtRteAJGh5IsGly/XNRNQDLt4rLRugEEjHF+SSZPxK
0Ck/F4BVN2m9eiNlE+zcHdZqVTNw2ioMv0AzvgTP3FBcrP6m8C8ntqILysBqIJDEQ7HVkLd1BpEi
7SPYsMs4ip57lDhWXunCztoWanIZ7JcU2rfxO5cvi8lahoswpZNBViVp3spG+xAqGi6FNGwFGs4O
whUCGHQQTpCbd0mqsM/4LQJ7AFLLvGHXNpSmFnz4wGl/vf0C6XlUe2Q7Yt0lQig2KyVEn4y6CCYr
CGksh3BhVhS445SH70VGU5k6vi93Qfo9ylEkDDhUe+725tCPD5cj7aYQ40ykFZNsMpB3dFNIlRbu
n/7Pqx1IgCWvlcD2kusN2XKYZIzT+pdQQzjnw48yKv3TEGaUcODXIP9DvM1NYysdmJidx82xlV+4
lABXFt3WMXgJsGSXDGx76LVfkvoLxbvtXcjbeN7OoYXwbh+2yQ0kKGpGXX5WYPP3QdHuC2rXKpEK
6fXd5ysq7OrtziE1050mGxHPitUx1jIjuEvjdPq4VtEsb1Mx0/GXQbn7k9GuMg403CbHogeJw1lH
zdC6GE1WO3jBmqjD/d2Lt/C7HP/m+z3DRrx+JzKNISKmNvd8eOKOsq9T3SUBEeq19ZmGCkurwP5i
Rz3DubM8fKiTcXk3/mX0F30xFzast9iN+TOzzI9SDG1Ty2Wr84inhmXpQGo1NHVz+mqIgsNUAeKF
yh+FulcfXdGGhDDzVUQUtnhgDgHHb62Ao/SZbxZoLGRfWc61+IxsrsImPTQGB53meeiKAVxEp5dc
hDdLQVTZoqz0RogT7KVH5DjNuvXgI3tFQTtjr+zqOtpN8CUOMKzCa+HFs8vwFfxl+2AJY8yJucjl
/2DZBMl478S8RG0wQT4m6ZSo5hKdhSKtBsRwg3Ejp0W0D7qPM8D3QD/WfwOhUqKkXmbcmLJCH3Vi
j5kDMGtoMpmcy/Hx24jNW4pEGcrgP/LEGnGwqB2U4I3dxkcRTE5Y8HnrAThIC1jGFSAgxXeKeDzR
dpFoiyWzO/XyQF6G7gb+g6ylt8mNihIUa+z7x1SQGkLQCJ1b94syNJjO/2pYthNGBU9x7CEK8nYL
zPtD5u/aQniPRHRmnFoG6Xcsb8yIkLj4RWfZDY2uKFqgQfhXRU7Yr8yXEqWh6mfMYBjzL8282GMY
dG2IBdKsxzy5LuJQzKbMvAa56JE/B6AUdl2X99+0A5RsSvLXyu0emPelxeyyPS9vIKGtYIv0ZjGh
sRLOfxT8iZ8eA9NLwdo8oIiXEP64pVoloVg1kml/k+ML9EyWbAeAs11buXLOqQOeUbXHftXTbcaI
P3fTvDQgowp3bZD2LpQXW5d2F2ft7drll8x61WIuamuE7/GKrw4IAI/DKuzJmr0juYgigDS3RmJg
n4pZJtwwCwqjwnrKR86NbdV/b3Cob5FoJvB7FXhJb9clbGhfFEV1wuwUN0qchL34VrBfrykscBbK
5R1N9z3HAu5yzD/jrvz3lSXqFh3OAHiYQyXBRMFCp0RQe8d+h4hF+wzYSTK4/shkfwXAPn+QLQ0G
SPLajx/2SN559D4X5G5h8o59ba2qztAWESNHpnIhgzlYRwVG/aI3Xf2tmoitEe8HntQ06dqx5qKr
mp+rWT8V5gUCgNYyyKc1QVjmVL1QSBKXP8BqMwFhITM4Yg14hP+amSdNEB801CtZ7AkwV9BUXFSA
V8m2yyYudqZ/oAgg6A3pic1R22/6bKc7UEwhI48Eh+JxZDE8lfR1tNxIvhWU4OTmd3fxMEgknB5O
exWTQymD4mWjO/mdPUQqI6gjZCIqB6b9DIFnrW8xfGMUi9Z4LAL5UhH2yXwzavRdjm9C7BSX+2rT
PZWZALRrZcx05dUFnwPf7Y6sf3/tCkmYhgG2tx3FlNXY4FAfOSDCgUsG+zkrDebXzEl3H3VsO/0e
1WBcLhFJN8mbvhfw+BOkuy3BJLFK2JnsclvSiGrT5DMQhTHl/ZgA2K2Uacpt8PKo6MluwS8MaVWa
AppSp/GqQsg719EXAdhi1HYiAddABAcrE8f1ZISZv1fZXKoDcxLjp65WuSs2VjkB6oSD5+SfRiwu
GgLeuBa43WJgPEhV45FX30KeBQv20O0uwKeaiQtABpG1SsHJeOlyUZELvn66vHjoobB8pES64D6h
VVt9msTl6E9fXoK1AyuTjplFvSGYRxOXJygzGFaXE+FFw7put9U4Zq0MBgJQJfXUOgWeVdvPgpsH
bHu9y0C5nz4pJ7cvKqQsS46+/4yIg9b9Q+YfDwFSVm+V9N0LQfuPwGWLDBK0mFN3+GrESngrgCTx
oSvpvxawwDpw3Ge5QEPr/8w2LVrLX5iJvk9g6mf7Mkxz23+law+o1KyL6SPAyeGokIpJP68TiUTo
8+uZPRuJCxQ7oW4xlQ4MfBWxAVpms/Agk1N8GjID+mfs3aqnQEdyW2Ll3QoFpjSk6+p0ltdanq0I
0NCJzF4y33PY5QOQKcdu6MhYL4TMz0TGeBlt3rgs8iG4+zsAhN5F8dKb/b/zRO3kTO6RFTOamXFn
qeRf11OggysmZr7el0nSmGxSMYadzyWxUruXBGyphAh2KLD38lo4HkFhds/feJTfNPXF60+GXD60
+kEoW74bw4WkPG5vrQCROelcrjZEWnJXApfv9H/N1gMEfumoaRPxg2uSZsbsYGWDbsUcl5Q+HeRC
ens0/YR0v8/MeIWX18WmU6j0B/OBP8c/zd+T5UjBPH3EdvLcvq1AzL6H3Rm6GG+p9cUOakXlXywi
OuiMhvlpVlHfud7mQBoikgPyFqr87iX3sPBPo3TgmelqCYs9pTg1Hovwi+KOJF9uyzErZhSkH1Ue
1vT5td3gE/PkW4j6PTQVtkopSXVzjCyWmb88QOQvx1G2X4vL2yIsRG410KkYCQ4IrbdEwq+NDC9I
S1qt5UTE7+/LtihelUxPsw/oBcVLyp///A15SWR4F5uIoj1W5IOrC/gdk3SllaNfh9QKlBOhR0+r
8wfPoOsVOleYRMJIV4IoIRc90k2yGPPtwqE1IYCckrHWmsX6skR9qyuIfmLJOqO8x0zp0HlW3EM+
gPHAdUQwdUpO9TGu31ptet4pi3jf9sDcZ0edygNpuZrJ8OtoR8vX3AEICHjN8MZDsLMwTysfgVoO
ljPYTd6fIzZw/r6QoBg1qRvLXUXHkXTYBmPcEmTpyqbdU1Mb0ptxNhqNCxaw+AQrISy4RabDTBEe
9Bd/AkDyEQlbXkOvUHayGucocK0z26oiDkHyfmNxy291RXF/LaDXao50nYYgk9qOPEs2AGmFQmEF
JK90rOY8BjSSXYJSUfGo3C+TwjS1YPdr4P/QHWTR3kqeFyg7wHy/jMdTyxy33mhWRvK9W8hwak4i
bb45SlTXzuVeKUGgArwEqY2QfM2mqTH4M2QaaJL5MtR0E5hYnmSeHmY71FlVUFpEMFQd0HCjSeFn
mtU1//jkZYCBJUuM1ImfcTKthjEDFpnmkBoFUEAaUrxnkDIDyxxoCAXRw0PQo1SEHVfs/3yzR2dU
pv/yv6JsGi1+9RxWf+mcONbQcsYAkcOhLUp/yX/ASX87m2+dNRBXZAwDpHO4IaoVPVRCqeoW7xJh
5y0cDpTCN4eEUK1DB9kTergtz3M/xBHRQyzmOsBs5jzj/NA6z/TGNEr9XRjHlTKUmWJW2sxqZm2K
FnPgqERWOVCmXIw2ALMO7cj3Z6pF1hGK5gBrp0xs2UIzZViPdsKnBZDrT5ltWkda8xuA4n36SC7J
G6qHklneblJa4ou2Cem4vKIu73I3rem4pcPQeDhK++iBB2fL5g3os/0394T0Mjw1cAfL9wIBM9G2
7Sd5vHQVHC5htXAkmuNxbWl1oChQ26B+UTJkns5kPh4YuhmYAXDhldNZRnv1izyi0cnGRIY5CHMM
k9Am7jgA2Hn6Nvl6RjFi7+Il8p2JwDudjCZxmomIVCVgyxCk27ln/SHHS9H5D1Otl5NxSoAPpNAY
N+LwGAS7diQ3GEb26ZmTYjcE9NXWqgv74LYnYjw4e13aS5haRedGoVc0sujXkwOgDdXMIT2UxoSW
IPE1s+VKLDtibOh1JcNNpdyC7bqJQyzOSJxuTj0lmomBp1a7ocqdPsCpk+wqmyNzXKmtCJDaXhtW
rWcaERFmwMUZaqMeEMySGzHKem27ocp8GPygDcox2eZ6dswvt+7jARquJ/rGy6qXcGkiy53zHpN/
JIbgRzfs4H2tUQuzhZPbsfXRbt8bbP6KAVM1ScmsLCIltCbLPhC/To9sjY7Gh0ZTzu7u2CBIMRCQ
53UgJJu3pWVmUuv5mMjuuBadE60qmOSiEp9lpfWpNiB0vrb2bwaIAhEgtVJami3XGAf705+Is7Xh
xFJhmKlgTZLfQhP9Il/+PjyW9zzxr+TZmRpYmladp3v8CQ9HO/LqYC6ZYr+u1adOqZtixW5M1owl
J+zxonT6VeUVaF4XvMoeOVLthO73X0IOjOFV530cMxQBK7XiB/mtDXxE85kUKFRCUqQfinFQgDws
tnhxKOVGjXP+Ay7a/DC0vKJzQA721dchaPKg0zOYHVTAgCUWuFFbUm1d52DubbDNdKjDCa5BPQk3
fTWGiVXw4FTb7lKp+vREVsaDoJWavjenc6clnWlOvKaeDaIfwyp2sBrpEb0ZyW1fvcdoV21NVwEj
q1FJs/LAzWElGFOMD9rrvXPbo9mAmiRHIjC++F0elC+9dWU01lkixmRgDEwPXn2VxmOwoUGVnu0+
98wgfOM6XBNeKz4XkvML7uT9NkoWw/i/L4vNgZA2XPs5rS1mdhAsgLYzacvn4117wf54ryndx+W8
q0AB4oKePQo1OOAeq1jCsxsfogJh6BJs75jzx7sOjgkY3VgUD3jgctrbBHpVdNDpTxiZT29v6sgz
dr/SyF8myTZh0FSu4e9CDeAtX7EGjAGfodwW+8zX/0QWzK82KDMhdQBnVO9StEC/0Ia+nQ8x25Qf
DFeEDWrczczVTdLJtPnSmSSMekY2TOpsplOYkkEI/8IIfYGiAUkTtxB5kbMWZPMuDy5GWbB6G5+M
FX6zGL77eK6LAQcinB8qoF2bhQr0/gKWRws2CQu6ohGkvVctgb7WPBbRHzln/TpdihutiUb4ylFn
3qk0PH1esdnfJUdI10M6FmnA67IgwD3xNZn16ZD7g1CvvHBhtkoxNk90w1i1+OTjc6VtFlL/I4vU
F96uOfGoLDXnd/y4M4DY8EDa/7Ksl6Ktsn99OO5UqnOGY0OWyPLN8hCAy58kKVZdsl+l55VeI19w
3yr5DfQ5tiMpXczIUhyVYGpzAfpYJ8IOyXdBdLpDhJUk3/D++DZeIQPakJyFLRNR3ggaBB+PV0dV
kBcEjqXbrdV4JAoCtbi447asVufehMIUMAfv0vTBwx7PNBYfH7mhC1WYv0Avmc2CpWK22hBnCAa5
jzqhYefRm25rB6/1kMgjPOwgWYLDCqCo4BoLJJEp+9PH5q9Iz4cuMcgmXmaJcZHMmfk7EU/TTvlH
YpOv3wB9dSuF2r4EraLORr+XeECY24/HMWtvwRZudpjjoHbyHfBv4uZgeKo0Ws8/+IHOXNQOQHaE
Q9g6qVyNu0vm/FK9n6kf9Gi+0cNs6vjjT4Hep1OrMR5g8Rrbj/0ZR+BaohN0D+U1ZkA7p/oUdWmy
iBi1wgg2zLHvFvgD2+rAOModz1/sixOTbkB/2+yECZbAo02tm2qxccKa79rsmm7jhiePWbOou4fq
bPR0kq1r2E5NUG7uZjgWnPpxqdLcAIMZX04gFSEU7PpC9m9Vg9ML2LoFE3qBXmz4y1t23tlcACYU
EdFif14Dj9AewXpXjSVGuZe+kiQOtGznXisaL3647ts3TFMKR2wY6Sxi5CPVgRe91nO5FMBHVMrI
HmfsGLcsd8BVoho23QExfkS+s2Z3pRB0vXwuR9F1DgVqw6H6cP9z+s3Y8sX2+XPU0GYjb7ALO5w7
g2esexMPjOL1xSfArt8S10nJpaSt9migNPatVYrlCY9SvKpSMA80K6HMzAhGF7iUx4yV/qyyuo+c
EqjZihKXMKwHXi1uKwiMCnyCzZajwq5yZIVpBrGgcFST42O0z7YsDxZM9+jMoANGFtZvfUh2Y/kh
Lajd2tkedrHoNtfpHa43G+Tuy39grWRuHhhPrN0kx+ZoPYyB4DG2VkLjSVjAH5i5zHGrRQ+1NEcW
mlfc4YOlCv9bLCpVtCvXgRSMb6BbC9prn5sT09I8VIG0decrLR0FPPkqeITSQB/tz8hqSVplf4Mb
QCuCdRczNDt0vt4ohu8JBZIuLDChEdR5RIciTmbqiKyqj2aAnRntHoOTuHvxoMwxsuQN6+GDGLMb
un84UPEDKoVD+V/t2Pvs/m5yNQtkYtlaJCLSqNpQnrhnBV0v0h1XpUytsL7Mtv4/TDvLUtIt6XLO
JzkiFwaQD1/XP71JgYaN3ZvRdK5DEyiEL9f5zxGcMZ3pRjHp2VLxNzxZyD/PAmt+ry95cXsy+n49
LaPUe9Tbr5LP5cURh4LWVljSb6QgySZIAyEywCrD7B5GvpxgeA4tzC62CAg2GLy2fHUw7E2IIGz7
iBxVQMM5Qys8pZlDGDryXaT4OsRXNJw4IPr2M9i18dpyaABtDfOm41aCx4rwZZQaJpSAp+Ldyjx6
898/IfsfQ3na9xjFV2qCEhybozOJzvtN885JLGzr0vLFOkDChmAEf4oxf0JnjBJBfor87kYzQwK2
DzCZNO3DDOQ4rZLEPwMG49xKodHSYyaSNegFeKkuHkwmqPODVYxCWpk2+oHRM5z0h5Tr6rSNvh+O
JzZ+8OtQSg8ZBGZF4KqmMgpc4+Prujn+pUBEhQG5xEZxPgT+IwF6ZqrMZsp0QO5TK5kskJCxCVNW
tT+CE5K+NawP65QCC9Ur9yTSGO5JWdRavUSbNGMh+EzHht4EbB37MB4dfqLMUkMlPnMou2FCIj/j
VlnHy3iDcnY3e6XGLwKgXMasJsB1Sy+1zKLJHGvzNaF7GDmmfb+9pUx4no0Y9EXlWNhNwjdPycir
olBZ8evsU38ZYtKb737tTMYJ3rJXQCV1cbTDgQAkwpB6d7sDLmLDgSOXbaCE858kRMLkZJSR+H5D
zYVZRgiingLzv1jZL3IUkxUiHQ4LknBiRm88S/jFrDvWjzLbNwi13xTDVxiepvlGh2rvaJkz1zg0
5+iPcN7jdAvn73EjucoeM30A3W9LQzcnXZS8JT1MYJ2/Yxqflz3hRus+aCW05dvFyMStm9MXLOJU
7sSbGtdAMV16dmdbWOQQL1b86hro0nzvk9I63T+1pwdRZtUdub2OsqNfeF08mMuW1Bgo9BJDD9vN
H2iH6JJdhVb+3H6ZlIhSQB5yHpeFtIX9B1F/xdEbAi+EpMQ97JcMw6Ue5V3YykDZRIYEJQB6IEZ1
psjI3qO0CZMB62HbCTmAV+fMswq5OXWW+W8bnXklIkVjMYNfkD0YH+Hmnfo6EDzKrOLlZ8esWOOP
pBJF3jZF14ggFj827tkHuzhj+5KVB3bvezycC8wxh5VM6fNs3wD8KFjdY4W8CCQQM7dGgwscFbnT
CEsJthH7o8QG2AaXy5LlyymXt+DUSF9BekVUUtCGOScpenxZjETOhkbjFJTuhxw5QFiCc5It3T2z
KFt+lyOXwfZdreeYhuPfM5hiX09BYR7K6TOjzyun62Qdu9XLMVFVzXxy6utePq6a7+MjEEdAuTSH
JiU1J6UGL+tXBKnd8fIrGERXLoyKi6bh+lU6oC7ykhaJYNChAsXyflk/C9md5jonqq7PCk0aHl1x
fGblknudqDl1VrplOd3DZE7NoM1MudDlhrErQDP03gw5sjJwsEJ6BVFNV7OCxWS8hXZD+sxoDchl
p9RGC94tFgM960nR+nCtvuUrfrsar9ZuJulW6P/mnKqZpi+S2S9ABFX/CCK9fzG5P0yahBSR9VTL
myMrYn+z4n3d0NRIciHxdCpjcnLd76KWA0z3mGz4BXq1LJqGX1Mj+CZkaSFeuXAbCQOJrsqG+FNo
vRf1pn4maXGAjQHvsZH+gWcC010aFb13aZP+og//ihF7Q/P727UvGxIhixNVYA2SJDVdAogbdMeH
+JThLwCXrW00rrXmXw5Pge6hqxLBemt6X7FkxpmcJjpS4VqB/RjquEZbqoToyx/dj4qezVc9lRpk
RmuMbeTldWgDYnzzaOPsN/ifrn5/nhDsmd8xMY+2RQJyK5e1NKoszQZs9216RaQDUD0RfwDmm68r
zdQFJFEDObRzhjqsXHH1ctFFLVqKRO0CoJXoOiozM7cjsl+t6LPCqIFFibxiF42vpruCDQ5lrJrx
F0o/KSMAAqvJJZxy1Q0J9inJTMn+3qXHKm6uSYm09AFDIW92qUSCo8mtMhz7F38XXfuxxn/zQJ5C
8aMwuleAy9S6+AIEVdxUaldNi/nGKY66wfq/HfW7OJM2mxwr48my1eqSBBYFv9TFPFgBIrnekP+8
wI05hxiTaVn1CLOcyVbnim6vFAHRyZGZsfegHGC0vXofcaEHoQ4OgIySPS6JTlc03eCK6lKxT7ZN
zaBaWnWa2acUcX47nKub7h6yxjZ60Z8k0FtWHIfEmVjR4Ac2aDfloiANQwTeyFQ2r5YBN4GAKxE1
yK1UWM1VkSudOLFZ+WVXRFueKh5dMbIX9Ezq5hoIcaVTm3Mdw5fbeL8El1CW2AZtCCJLKTytabCK
hyni42eTX+F1LxuSCYfOy68vQbcPyAxBDs69a2QJohDWABS/6S3EYAKxjjK+ohO6j3HPKNyyyqdW
zrQCEqc0fdQ5fIJ9+ALvFpinspxExyKs7lFlZNgO4VDW88k+D1dX/e6c771mg9PJPZH5hCSHBsl0
pzW28e7MRWKs9OX/oVwx/b2GcAN+fIrn9U4RnypO/0norG3QnWnJnmgHhKYjmRXz/y95XM6dL7lu
eTYEtSzfkGJ1FOsY+u9RuJQNdZULQz3o+VbkrB/YCXEKi/j/9a4fkbmBXqsYxN3WaCgfxmGlRxZV
dg7weNF0MHLVsA4tsMnfTMMKQTnvThiqgzr3RR0mNqFaZcW1mV6XMGhVwYt8JVvtDjtcDJ8G2YaB
RxI6apzVin7QYXUSrzp6U0YQN85QL14jAfnBpJEvGZRmaT93TXGFFCayQ6es5ZwdMUIxpiCWZBx2
7qI2xBTo5LQ+OvUGkhJvXcOJnnRT1UmSohIXTzrzDdzX7ZsNLrYQb47K2m01DmmnM2FFUnby3xhd
wvRW/p/BQ1NiGSmarMsnr/5jOqrYr2I2/s9E44tYumaeeDdaycsDX6rDai1CA2zMdrhBePHGSM5B
mepjOZJRueLrypqv8aGwQH4GFN/j8bgty7Y0GEky76OHrdyfzH4l++segNA1PZNmfBPElFVZCHeO
YhJTOykYwZwtPnDtf90ws0Jl5ApYJQcGGFaXkciCqDBRYvuMYY9PU5aBwQFKH6+dY2Tz9d84Cy4R
Z2KT5iZEI+8tTnYrhBEuhZnpFwhDMdOKEYH3iONPfBDVL15Hf32+5xStfbwNzpjCdLFwp3ik9tWB
LJIS0vnc8E5kgmlnLp2tqpaa0puAvhs65Gi+mADa+ODw6XSRHsfBbkGOV/owdbj6dM2BMPQdySrX
LLa5T+OO6lB4ho7N4ua+H/lohp22cHbsnHJigpt0uAq85XGy2bIlSKo6C/JOZOXmkbm2LPRpQpL0
5PNeze5uZ1eax5cj/Cc89jvt8fNzcmjcEeFD+UlEVrnTzJas1xXhAbuolpKBJdad1PNmDkZ15p+B
mcf2mepQDm4TA377Gu5EfCbamhOVbzyhLHguq8ooSlm5w17dxWBsv40md9XYmHriwzhhRq8HxRG5
uAFoY0IpPEhNZIWkuFd9gIMEhxjmobOn3MtGKc7L+2aH0q5kAmuI6/j9eVnQuOgsOKUjsr/mEEAd
WvfbDt/Vf02iuxgFLV2+0xiyxTw6qs7o0dL+Y6SRRH284U795cFYl8BlJioxdPbGtqCB1EyHRscD
QIJi3u3RI3257wD0O0kVuP96osk1XNIpLB/9Gv0cqfyYHaG7C6WL8mFq9YTVPb+zPnyPHkRIs2o0
Pa3fnpy0YyeP3MA04PGJMY6g7BFFh431rOBJDwtDGqR9cuY7knSGNblfnuXqLHad8IpzXnRRzhDK
EvDnTRln6SG1CrFGFM8YV6NivdgIamrH2mxTbryQlGEsbfezykRyVxsxhGM6wJKeQFIR0uFNZxbT
8ou7w1ESPow4CzAuJ+65xb8kv478HBGPr/sPSbpdqw/cEzVpiEdfi5rZOcCoE//BEiN5EQ+1II1l
Y2thOo8+zGeq55oL0Cx8YIERT2hCXJgp8mbMJZiT0CYavaCHfU1PoXuTMw2ue18w7eI+eowYAJ7q
NHLlkJG+a3mxvXRs1EgZ6DCYaczkpO40oaIQz95+XUGIcfPRaF4IqwVW+1x02kXCoF0tn/52DSN6
jVrR7tA8ZCJPJM54cx6Bhr3i3wlCp79D6AuGrByahnRI9CK2VifKYHutrDqQmd93DVI2NvNTHEOn
/QgII4qjUBFb18QoV/wO1oF81wcNW1oeUROA0yirwJMH55MO0gHuc/J+zvlGxhXX8lx63xG8rlNz
BGAGs7DK/7ZK2SR+v1pEO7b4idKZJ00EcsPzxOhV1eb8H6K+4LHOXi7aE5V3g5DSUOpni08mDHFi
6yjxVAmjzX6kNCqpqE5ni2guYahd0IG+s4uV5f2knFCauYaVNPL+C3FxlGeDi+zj2jHLlZ7jgXOZ
PP3w/qMxCxJAkt0LvsYB9qUJpYAOhY3Pbsd0xVswerirYeN8PVqCG/0cRWvwj38st0If4gow/VZD
DmOLyaIZoOuoJ847V1OTvb0/tIhpPuwHvuB8Osdt+dEMH0Pr3v97vTDAbZTnhSCz7GWB8PZWoUkD
UhUqy/iwgt5r2N+03rhnfnEy0ejhyvUotymGxLl9sbAPVUrBhfhj78l54TogWmHXlJsjRPQM6xTa
p/O5KIQcyZVM9WLoIFMDX7OQKhYCg8WLn0ty8eqf9kojE7FSAVdyj2WwjbVd6k1A4Hl3ef3+vXQa
qUdWQL29MJhJLxLzQ/2LvEC365m1hdrx+hKclAEvuxbe8Z7TxbQpmG5Ki9vkRhUakGvfo6LV5jZG
pA7maBgSgGqOFe9l7sXTPppIb8c3nsN+g2rm1rqVG9tOWzTz66uYTsOswnezCVgehHGDHn/JIYiz
CLpD/6eaKduKsbFqzBtcxlMv1YOP4qy7MxVuftkQNz/6/XSm1wWVZ97bV5JyMuTaqVlSDWCGekoY
Gx80fu9SnlcgGrPka9BPHWtzr+D/QKgH/WoWH71ecnSip8m2moBZT/aJsAjyPIXxCRmKGh6Irg/u
RYbM67Af5LmqsbumWo631R3b+p6sAPI95+XNRnoDyWoaEax9WGzZnpBJ0Wv8LhHcbQwYtOoSGVzb
chOcJ0uCuW76aaGXa/GFpgBNTjaF2gTfz+dH2G4buiCpktGyOVg6uqe0a5Pd9NdlZP3aUGv3xUwY
KCNgDP8YmjyIVO87yWLDF4ky8A3Gv7XWFX5D3/1a+qSmu9LRFfAQNYpRqxiwY037wo5PmsIvO8kp
8SJ9khGzbEBxGkJ5u2b/WghFNghxbUbQecXP/8wukwnWOOWMWbCQinYOMqemSQFV/z2RliyxlQ5B
DvkU/6wDYEqWzrfeDJCXm2LsYot/HGaIC3DLrjFjvsqrJwLoumOMAXnJLKHkiex7XLNtzVEFWdG3
/ZxeXuMlI0VQVAygC8nX5EFtIdIHAyyu/NNbY7a3W9gSEEmBeXWYUAmmSjSog8bPMd7taxslQEOX
67783+P2s9bi5/46GyABflGln8o4/ZmdwCvSFPAU7qd9eFtKsQ1jrTHoVFLCBwpaWZdvYB//gMY7
EJk1RQQZ0tn7tktbEyLAV+aAVDBHEEmpAQWUOCetR+QxD58evfNRb/8+SLPuO2jpkktLgeYwfsKO
mpfNWfWmEMoVSiTz/+xG3aISB0/yKwJ5UjJ+MUttH1nYI7kyNGYHwB7vszF2w07TfuwfTtn8n3DP
d/d0KxHZBNGNNsg4b4K5Hxh7YLzO3Sgxkc9RnJUVyMjz44awHroZVVZHwGTH4A+zkMGQTvone8ln
pR4tSWTHdd/K3Hr51G/68txqFc1H/9rEzkeV5WeJfUACnVCFS6XcyLCeaMUvtp1HnhFP6Bv/Ez2e
R2DhP2EHN8HbgPvs6vT4SznpiZEVUV0xw7uMOn/+gpNqrZhZWVsu8qREHrilpBGYAO49Cj5vUd99
TYhoJ/RdehtHg6U8MbPs1Q1PQXdhhuWoB2+9nduOqvr1nzWOFCTioK31f8F+PrP2jijOhAv0Q0Xp
3S2mzwCNFTM1RkUTdxWaHgtOBpG5HInrBavgcgHOT22J/EgO4UvoWhkpH66Idrm+hYJEGDgyHP4Q
vnw2MlVt+LWlaxXdxCZQSifp9i68righnOI5W6fw5GotVsQxAlRBxT0qtY6NDiS7LFjfp1JpCiI0
ri3SpV7DU0vJxiA1lXY1ToS4t7fdOKPmSUhxPGs4NaklbK6TkgyeNhswg5xgEoo5WMDK+vwI8PwD
YZQLXxt6PhrDlx/xkNz9uAcW2VfqfRFs5q7Qm7fACV1ixSLdWKzxH3qSyHv80DORksMDdLRppCA6
+l9qDlvObhMxYeo9JjeSSq6S7HFT5UrHE0BDEa7ZgHlMOE+Yor2azGlbbuiz0Vg3Eo57I1bEOW+B
/ATku1aze5UB57/MlAaFlsSYJ0azjjXPlVL4My9KpmHWtw+Yy/SqLCwjfffiWAopdi4HWta6AvSg
4jOfnWbZp9F6y5Nb7qbCkhBRCuEMkXHxsDE2YRxHFwpHk8YWNAdCP8hoqqwj50Yo65zbuxq8aRkN
SPdoOzBYpXiwz+zmAE9MohoQvgaXz/qRx9wcTLC8ZNDcwLFyZlPjd9/IBhtzJ6/WcOj2YcvT/y7C
GkFOOzOO2QOfY0lJ9SMoFGw58TUHSyyadBD7/SUZn5QTEWxy+ASzsVgu3xvEDpgPdoE6VZikxASj
JQLZOZaLUI9Tau49RPBW2Y7gz6ebAL9m0mCgyj421+LarMBCQRIscwdaWyfK5gZe+/1luXUFs7xh
8V5xqvTwOdhdYecyD9N3eFLYO83H2Fdm/03K7xpqhZMxygd5sPqHd1Y9SQgC3l1y55Bn8BMguMXZ
3Qr02UPoAMODcHrPoUcZiylEJHPGnX50Kf7jaOYH7QizpY+L+urVJTw8xUQzQhAhWxVgVgLJXWZD
skE0nZ95GNNllLxLYpkU3abpq27It5FuqjC1wwV0R5ZAU8ifnhVqpG1Cqdske/ZbDY1kKJej9G/a
np4r87Skv/Zt9DG0SDG0WfwE3yOm6PG4P8gyLt0rwFbZ2EUIydU/KhoKT7qT9ya+MjpOYc0DJoMy
v8WEjFgY6flDCQgdw6oMOcJ8CTce8xcUz3KEmgAJLxHOnFG5DSyAhyGdcSbiJdyCDPK754SYjgiW
HfsdWeeSoOCOM9fGpVKHMtU/FGXjlQfqe9mJG98bGZFdPDn8j1ixy/fvAavjy5yEAgbdvmM2QA2J
vGA2vwew82ONUO61D6VhzJKB/uojI5zfqX52wXQtuHrXv/XNefUzoloGlwQemTAx8Tu5dfW4ZNHb
ElPJhMMJXCpi9OBqBq3vMJnETmeBooIXpBDcqd4qtghMUT2R5Bo6j2ITQJnKQaewmoKRYPDuGwdA
fv4Kg6TggIrKx9A+Yxnm6kT0yR5w0Ig+6mJKr488hr6kSyG4xmSiteHST7MCzSOuSvELbIymVrBs
giDtlo6OxpjRV1v1mABA9v85uFHcZmJUK1BfSbXXKeSAPNfxaMrkZ01VkJrwmTnzDsZzTVFYG9mT
N3gl5e+hgbMcw8WnrNxu2YbshZlU2PgfsyVexPz6nz2FRbVmB6cbd7ZB9LEPakj60BB/jOR+XbR9
mC5PtyVXF7MGaVuejEXkRa0accdof4M7U30loO2fK8TuV72qqqYfkYRdCI8WupPZQR3awYcCLnfa
S+EK94OZaMScS2lMBUan8mM+GRetPi7MndlE/UuwZ5E4aSrMqTVAt4Wd4Z5r+k/cYf768Sw/yVb+
PDDgiSF2HgKVyhHMHqgt9clE8ygeXyDYm1zN9s8ZutozSJ/WnMDVhJ2ppy8OBKDsRVSW27Szht0n
PPRoU10hMXHHL07TvqG2LG3A0yZy67H8uI77WV0xTN+jo43tk9NC5kC0IxYZi4bXrxFNnsxDkFjy
z+8LU8vPEgsaMIezb1dBm2PO9950XySA7jp3J8Gkqjr8K7mc+V2iJbe+0ojBSWJCr4sO6UnVIet6
DZ1/c8MNOIB7RrJqT8WV73qXXOW/CG34Et6doU1Tg2yB0LDO8YvsSYBZ6N6ae2msCj+yiV5Gz3oq
MhUzg1nyuIskHn7CKjQVojTv91wnzakLlPY0wGgjumvO8PsMCru5Ia4ktRwaqiFxDgMMY3lXubcr
jHPyu8NtCM/BWfadB8hyGeSKmRR7aLH9pbWPzGD6xqg281tVqC058A0Ud9JnHIUUbGr0TBLpW9P0
Or94GOE+Lxy+TKdK1wT5iBqX/Xy7QafPgyGiFm8R4Z1Sew3rGpm2J+1+R5W26B6mPKWztRS76OhG
8PiUIRcYxZ9l/d9sOhwcSUijoxrZbVPqGFK/jgX52qdbSZN3Qo/mMcWDe/m8OhRhVuNnL6lWq6El
mkk8MpvdDXJyAxe2p0aHMt0DniBqCERTCRGvhP8OJcFJ2Kv/w8nqY88LzOF50Ozqe3B7ry4FgqZ8
4pEWcaMcNiN9K/yBu03JAkeNVh2WJRfF29kz+PXJUMUljTCKEfHdL/5Qs15ZfdtIAUKIx59P1VXo
pWfOMN/FHDnTFq2JELdWASYoydVxadBywdgqamVox5coiydT5huwsCOc18VUOJt3djZ6oOPrPCNB
oXevQb3w5ylMMdXEXaTs2PdWK5gPY80RbsTEHT7w0Qfn5FH1TrlxLAOHUStz7Acx//rd0m/cPJmT
qhyDJGf4kN/OTgX7J6gmvLAkpNMVr9yt8JQWvYKvPFOfQUN+7t0k+GcDqxfU+yAJyHavCEAUx6su
LBtn5ustPEUak+RmDxaH5hKKX2BaUJpwEdJg22+A/uS9rbFx8pKa+kZsT6H1eGCXDMJ0iracjsoM
zucoQP6uKRg6OkEPPxugPEjGoZWIF9GgcPG0ZGzsqrD5uDmL9gmK4MnwonEy67BQmhKjfVq+Z95c
e6ChxHV4nzrVgeH865vHs66xHv/ItN1wNpCJI2f0AbYV3Uh4oNA+yhhNHMnPayHPLceqbrWRen0z
a98JLLQcQEQVpTZXbrD/JuSXT9mdcSay2qw8lC8Ehfn1eMeo/XELiXvOdrcBTAOLZvRf/mRtvCE9
WjrXwe4yFp/1QLi6naQGC+ZNV2ynBxxxKkmyryHLV2p7FxfcI/2kV5tpa7bvkBy3ERoAD+eaeF/B
5CroggokHOv4UfKHfR99CnmVQYkXivrEV2h/W1XWpwf3lldmYNtqjqDYbcAsYPcE7zb5Q4TYWv94
oGJGOw9sX6wTz3x5z7UVsdXIrggb/mGPX61ZLdceMe9pc65tObSW4V8/JHqH5vHlpeSOdn8qAaBW
v/lo9J+bHov3J8T15srikxCVGQ9dMg6Eyuu13tZCl0i2ff1++kzf3Kyetvz493e13mgB73ml501F
XjsQcJEsmsXi+pZgk7F8EplSloEG78OOARrNdENsInPDQxgy/kN2t/ZhvwfnM/3gOnQ+gHRYNAZ5
BudYEqIn6hdzRXhc8pPor2E0EsdKuQVNikTzJT08cB6RhPn261hbDpeYtKVym+DhZWP3AS8MVeQr
InbMjBne6SIngCVrjLY/B4p/Y2kYw3StUugfKAI9Q+7hHIYVbQwTULU9xjw0UAZJh7AO7NCIyPSO
7ZunZdgqdadvw7EJAD6JhttJnW27KTls131u/fqbhmSVw0jbS84/uDTj47sRGbv9JZ03XYsKeQlQ
v+V5P7PfRQxa8lsQ8p8VBDoiN2ZYqbbbV8mDEY9FRgX0VAXXMJ30l9raFq4fdDahrIOScWoXse5y
TDVuct62VoMeJtzMiLDUghOMn8WHzSiPokPDr/m+0nDOzEa4cYo6pP77pcIAxwU+ovpRYJzolXq9
AZ7fs1v4hmef7vFpPcaM8XIvmmWcaVWqY92Ir3LuNYaoBZxfqXiBEcPPTiCVmblh3JJw6Q1e5jfU
nxRmzreg5DfVx0AR/5LiFlRVMdM/MLDYsM68ojNxfQ64fSRTmONHxeqyDJKz9ytKj//qfVf4HBZu
FAN3uGbP5LsPWMVL+b/JkxWQa7CQ2eo8Z6IMIg3hAEuQJDDTbJulAE2olu/QR0EXqKMbvQW9zKgV
H2G6IpbSyk4YCSAj2ClhYwW7+qqd3VQpmFEvLdwIBG4YOsgetyO0lU+G+oyyjbhJPOUlEKDgaGzn
HguajVMxyp2h73DG3DeIZXgZB7z/aA6ZujTBdAmIqqqdeAuH18Lsno6EqmeEgD7On2acF9gn77fN
w/1y6CxWNZ/N7UnNB8wQqrZ30HZCVJVqdZeQeT+VUP+KpAKyNMMer+RUoqMfnHxMdnXzDsGRtxl5
AfJSAUSwussOWH31CLXteo/+9M8ngcInT3Psyvch8Hy1dK1aSKWJ//D5YsleSPmW+pJ2koVEPsR1
JMbpmiCzIJq/4EQFkIfo66aUpL4rHLGJaaXeZbKonWomxUgPvKo0Z3euNQ69FOD2xNHVpTBQvHbW
g0gJ37L8BQ84jBdzz8Z3esomdywAXy66hVjYh6UA1obeKmE/XCAntDDUlVvYr0RZw3pLyZxpOby2
WJGLwYvomI29HBTIuIfsnlxlA38mQPvXIijvRhWH6PXspG+fwiXcwgrptB4WWcTXXGrg/7Q6xDt8
li+kDYmXDhH0OW42shoQ9qRcYsU4a5y8lcwHZn9RYXU2/E6RmDTHkaOeOcNzLuOJ5PVoeClao+RC
cut6tJcC3hR1ymHQT6/zk4QggxYCeij8aR8cprWg1abGJY33Xy44pBXZqtuAgGt2M/MHNd2hTwTx
W9rRtQB79TnDKrnxjNkdeJ/iDeueM+zHozODNsf19G5BKJq90/KldiTcZvt7YlHa9FLY4MgfXNN1
u7a1iEB3DpBoJ+0SRXpjIL/uI7qQP7EckTcNaWrJfxL2+eX7sOKK6r5DSo1LN95ah92rdkbjzVC5
Gs3cNxFV0VXqJ4kRUyNuZj7pBkU8DOuFR9kDw27N1IN7ghl6JmHoW2ZlRoFqhAQe8vBDChmlFrs7
RaYFMIy3GDZbwI54TGOlb9OKji+vy47aD1X0aDXi785NuxdsUTpMHOaVEx/qTrBMGvLodanEffPd
zlRBqp2wpRJvEBQVFohQA5H8/bnJTN3w5qHk7UPiOi0KWyvQUIovpZiebhAKRvQ87u092BWn661T
IWNdQ068QNEKFUx9jF84LbMiX7V86Sq5zLbIzOVPnuNsGYH1M6ciDYH1L+CoYYhSp5o8RiQFI7VV
sdwNs0MRKuErV7yxoQTRcG5I5Dw+aj4D+hlM64cJDAS8XXrodUdTm5VyUI+DLkMyuta/kQM50AHx
UVM4N6efbzcLg2/0559oR8DANth7Ksnq2IaUybxpdpFatGDLGTGOXiNw69qWWpH52NL1GuDLIbRr
h7XyEiJEPIeRz3csljKx3Q1oXWCgrNWhBQRKCn1A8z1rbHmv3Tgls2uRNWwpv6KyIqbVzkgDvOdY
pln1+O+qf7oheURIIIGrlEtwBJkak3uJ2+dadIZdJYzZVarXsxx3nfnhkEe0HpTnsA8CT6Ln20b7
fAweVhye/oXm28RXPoVi6P8U+CnqLAbmKeF29Ot6Cn1RXenvNxqkE5KfcZijDTdWdO0wHOgE0MbQ
h908dmyttZP+ICkVCvOLZS6Dlq6pcjKiVNPBJd4rNzQkSMbKeJwlqzZsDB9vX8pop2ceo7uEWO23
Bw5hDf0pzPaUc0T518gEnIJ9OpZBOYoIRlaJaSYbdv8HlHeGCvRbIqnU1Pdr1Ax2CSB0APu0/2dH
0yfJCexgpnTZ96MmDOLfyNMIlOu1i2PaLrEXx3+Nbm5ggJO0zvo00mbod7M5vql0NVKVYCno+m3y
xZsQVAtXTbezH0/EZG+hh/8ZoWS8zgC9AdRiu1j/WQflbCpXKjAPcoDROg+k1vGxV3N087Sh3ClB
TU72Ye5xUnXpD5dr+f3q4d+ygn4GK0/xZI9uUTikBiG6rtc8DmYV6aI20WNnI34sFt0dqPxJWHb0
K+6feglq89JSBOETDFZ0XFWIbns4cXxrSB5VDoXbpGLZtb0uSTQH3lmKQG7wbavk0VcnCXsRFiDp
nfGhi12+Aj6Cubhq4G5dMn7z6uVOUMaVHcQ6ex6RfxjngsN9riS7+cTaKbYF2RRgu9Pwf/Nthek+
4HYyhOQDI6V+QFSEol4LzssJa999KFaIeptsmf9kK7AYV0UvM/475sJBk1V0um6yDGWKoASGFDKa
R9howBs3RpAVKyyqZPhLH7pg3rQXBTMSPmKmEZIt2KqQLfeWZko8LiGZbOfXBh7klAAoRciiPZVe
e0CKN1DFXIl9BMRgd2BH9QL4O5Sq9Lo2PuF7+Noc24qg5BARo9N3zkOGg57mYUWqR9jOA7+fCUMk
AoggQ3AcRSHWWHb7P1/d2xr6p7Kmyj/TQMDHPSdmvACup6jCVdHDhY2Vf+0bi9cC0d0O83LTIQ2M
x8xJRd6FX/vK/LUzzxBvan/nYd34mSNa11TWVh4smdBn/VLBBg5Y2R1SkU47W12QnhCL1RPM/T+B
NrWdcX94flL+N3KflCBaJ8ir/B0+ZJTh1boKLPYE2vkT6d+qK/8TY50OIcXNgDcNVYdAJMTAkBuR
HdrIfCVxApYLL6hIZiWxd0Jp6nJsx/bdTtQy+SpgH4IlE2CTXIfA/LR5MPu9ZCNjlStld2JaQz6Y
FPTZFZvgyrGpwER7BudGjm3wV9ufKz6CewdjNCk8i6ox/PhsM0gY55lBl+G3apH+21ChwEAlrl3e
1NgROY7IvEu6c6gPWv28MHMojtP+Yed4maTyJUazqanwX49FfjD1JM781E6OFZ8Quda/jPAzW+K5
my8IOp6haI+xNXbgF4hggTQcUbGhrUDfwx9Pb5MEBD/0jjIKfaepwYYVlISCciQdnYetb748WvD5
hsEQBtVbYcN0An7fgxACI1z47SNANlfXei6lRcdRD9NXucJ8prV8D9KFGoYs+LliOGKd/THSZAin
Ol161gaBfZpFYUOGrG3jmfxYx5I79C3kxNsSOluByqRPvg5N3ENU3YipJmaNl1qZ5VILT3PRU4AS
IVlSKXtmEjqlR71wJLVp2LIOXGG0Z2nzabGSgeLhsygILTO0PI+k/oGtp8N/7NvYE/k7e/YWtKs0
bwfGeGmXN+PwC3i5FI7qZ6HAF0jRPCjVp4bewfd3oGVWwIcJnk/L4MsFJv4EfPc7BUQpDfhsJsEe
CBRtXT8icZmFr7aR5eJhbvECp0x1YoQ7FQQh6ff1GU0f40O/w36y1CL7jYw9rR8RZC+mTixp4TQc
Liqa+BC1LKOFmThCET345Bb/4vAK3MBmGh6/Eyw4niFxFHknvJYBSz1TmjVrBZk77XQyX7JTnQy5
dTbuK7mSijVz5L5xi7otLYRdDZwUuomzkpOre7ka/gEcCY5RSjTdH9N1p8OmbbY4O8B08nWvPbds
BJ6+sv4b1IsRP7EJwbfu+8S/HrypaVNhwxfb4ZuppkHum+TeT//5zOxOWdzZxqqfJsNqY7pJLAho
JeCC8OQ+mG6e1bGbt1SQOaD/3VA2pqkOrCEeCE5By3I6lAz5GPBbi+4GFsJ5WSJVxnRnPI6jUsGD
Td2c4FJwtLPyZWeSrpOiS2B6x3zo91phAWxMx7yKGlT45b5U6NPHJF1frFNOyVZ8aGSx1SS5bj5t
zYAzccg8yNTNPfwrT1UrZedDfkv79Ydx9EALcFCDP/d5+i3YDfyhh4RjkzGOSgKEn9u24/nKEbCt
J3fC/0M65QUH5mtFANAh2jwJ7Y1rn9GssmYwppABGpKmJEznjRG9bsaMj1xelXqxca3Z+C0pWsH0
W1xiHCMEVX2b/DimyDZuHDVgZ2C+y5+k4DZTMnmd1bXDGn7Zha9pcUkwaWKHwAm3EWLwjpkdHswH
jS1dDs0xemaHVel285xXMYhsROio2E1hlUqXy5vdP5a+/bwBwdh3d6llRuaOjRA6dlp+dxaJSbrB
YVPTIgValUQYVOakb7gy373wxz8534MRF1ExcmSqceXUiTPexTpJy290zu7MrrRtaWiclMDj4VyL
UE4gNLngmzVI42BAi16snhvXc3UCHsYFMpcpYI1O0gbnM1W3Nw0PUx8/kqxJLG1sADNV/KWuuUOq
ZEPbTt6rWUcjATbQdlOYmkzhVdn4JabBNzaIPbb78Mm0W57t/1Pg44fv/fzvqkNng9Kp7o6juUYP
v4D6poD2d4VLZ6N5ApffJtQAjmYZgngyWq1D7oYZ24jM/0IBQLXr+RTcnSoEIJZ3xhDV9xI7aKhm
sogRS2l03xbc3iAL3CQl475Y8AmwOiagDdlIj4BnECwmq8gGLHa5nE5hG8lCQU3HBauRNIqbk/50
Ny9Uv8UPjLz0UEH0c6PRtrnDQObf+zSYalzMIDKCTuYF4OU6Tgu6epW80WkYwimc+7MWr/CNIFJA
IP57dt0sziMesxGEQZI93kEXX+lCuxvh1IA5OJ2X27O90LpveHtyGCT+gOUNFdLYYfm01I2Xi6dU
prKm40CvFZHgizUGsoExg4HWJB5pxkywcTLlOl20Tjtf+KMjdT+Aw6qKThqnP1abuhBhytPQ3/cR
F/SOwxYQTX06+K6PuzBTSUHq5sRdClh/Nph7B3+85j32EWRVvHo3O/3iFNR0kvG2dQtjcr4TOS0Q
sayo0Tfjro/P2ij/JXuD6I5PUMCwgwi3pc0i1ARCCJ+iUay7eworOJZQjGHRXhDw+HTAMiKKvo5d
z105adWL0SsAQxikwqsvmoWwxQ1fxy9NnO9E9dZ/EnSe8d85kW9CgyXs7Zt8B/5Mgy0QGY2bgucm
D09BVtL9dzjZrCSQvMzWcVxPjEZj1OIkRq5vw390PL3sCekrvYfHw6oSxd7hg98/KRZgQSXEXbSB
2ZT8CcH6DpAsXgKh/YLWlRUT7URo5BSg2qpjB/YWO/Ear0BKqEuNxNuSi9JyqMh9EG2GdJfZTbEC
5s0IIeCC0z8nWsVQyN/nvi1DuE/uFxQXBpL4L3gydJ9//vcqApmcWqvjDk8a0AR+rk2tXSOd+PFP
avoaZFJyEJ0eDOJ+2eV9F7TtmMYGRqA2TrNStrwOj4Tzkjaed/vLfKOSl9FHZq5a/LCjxuQCWlBQ
KKMwdMPHArciyTNbT7ksjzOs3msZu5hP0qB9XngLk3fJAMvBoJQmfCpz71ZsixFkSgfpXqSGC//Y
Empa38XNLOOrMWd+osvv/1W72IDnR3ILdiyAyyLaxlhUZDEkjPmtnXB7fx9aNtifnyTfvmV/6Yw/
qYZK4JHrA4JxmwFfXj72J/OFDoTUoPbAWPnFWxt6ZH6xRyOh1RL/nVT1ySLnMgNkDUMLb+JepoaC
X7y/2eIhbW5I3Tpq5FoAsZOCcxhRBs3yu5urL5r0S9K6fdFxZWvsY9wWneVWr8OEx0+DIRna5gsk
wpf0nHMjGMCQ8/z2f9+lptx5kPYrtW8itcsW88WBgbErgVIHmv8q55rLVjxMTxBloT2KUWvk9L09
Jv9HNzXwAtTDdiVD6aZyrTsxEuCJ9CHoJoMsncrE8aUzgjEFuKJyR32sDI03G0Fy8Mcu97jolb1p
euW/to1T5Es1bUoaXnQuKQ7FJk+HuYGU+Xlx3SxSbAepUeEp6H8aFFDlzfrjaNizSNSkdRP8b6Oa
L5XxIuiywbpL9Dthe/x/DawEZnU40mfWWXcDnaNkLD4Uxrrls4msvMI6i4w3LklGRTT++OHvQlS2
ZI/pGwQBUmWshLvB5orNu5h1qUMEJ9XjBk4alfwfvRZr76xS2V3FbalDAoxi9YZKLCr56l+oWLFP
R9/2pZaTmLASOlUI+Xdg9ASIwdOfbPC9KvnQ/EbRrauDRUbQvvOwmCKaGFWNJyysekVEK0oJFqu8
0n84NvXaVmcLTpqcaZGfXim4FFvzgaFJ/+gsAs2LbadR8cKFT5W6gy50Tmumuxo7VHe7R4hx4xyK
p/28MXag0UEtGNlIkvrRm6Ua2uKWBDnEwYNCow2GWPNHi8pRtxtjX8QhGQ5u3xYe9Z6W6Bpy49E1
aSlomv0ChVXzx4HtcGXkyhrPjX0kDuIjm1C5o9gwXT0sFjSrGbpnSWzuMLno0whnrMSysYPKwU19
yWw9wWcaq5UIFuDC1q1gJAIxhNnk3sxEQvtl0sKgPqmCG7ssErWmcvEZ5zrBbFTw8RS7VjRsjjx1
8bSNvzi8vPSGUvDMlwrIoZYOcoW/GM/+YKHqFHP7J7NtlSIi0Nqouuu+A/7aymus7eI6YBT7LSss
hEuGb9yG0ViAdZ3IZB8Joq4AplCoMM71yMsFPI6tykCfcq3spcO0Ymoka31Dzn/LwKaVfASF+Iqa
UmG1YndjFcAm4SeXuFrDV7CMGnL+WoBszyGzFPg6yl/Sr658ki+kKg8dBt3JDygfh+udsbDWS3Jg
9OeXJDuXZ/k+HMqHzYdJ8E5gzT92ZRDXUBvZ+RxhO8bFkNhuodWvI7VUUDa3AUHQtbq0Ml11KmNP
nI4wTh5cNeOY8PBDD5DxyK0m+cBO836cGDED7XTCeId/1/e5OX38tfHO1/dc58y7oPhO2Wq1IuFi
3OafJA1pSXmBY823vNdRM/Ojxah4StERne06LBs4sOiB4xpGk4Anl3fx8zhUcmrG6KF1N7TTJM4r
BTKzDGXS6Hnc+Y4hP9n+idkF4BmhD2cs0qq8zDemej34uAzXuMFq7FZGioiwM2FxuvYpVXia1OGi
gPz960LuBWBxIwW6SD8yOiNO2usY1dSs0aAKHkzFGRK+auebi3SaMPpoSWzQ32VHGIzZmMoFZ4jR
dqxCCelBzj3EjBzZlHFPs3IsjxXGEfKHJgdKp9Q0Tf/u9xTS2VVUxFvlux64VXTsn4GGsig1rfG6
OSJrkuebF6aRHo59NsDV9fk2rCRvgQU3k7hqdB9g4tiT0MRqn/zCI6yYPvwTxkUE2TxFxxoxS5lP
Ji6KvsD2fZ3WwU9GthM8k2+BFPYnptAMB67/90i2VVPfe2bzx6kZD3FznphzRgLl5nLZv40g3fKZ
0VNkM1pRvsQnK9HWaxnkpYTQpyku1Cd/7CcrkyMVB5avdYnsZVjBpagvxsSneOVAWMp4ouRccjjo
/5YGdoiBtPhekO/DsEu6XLfYts7WppoONAKwIO/wpJuk+BwqQIVNlqCicjZBTzOjj3XkYRIdwCfg
koqpHGpaGhZwICU8tbK6itewgzNB4+hQSGZIgzPxMSkzueLB+8r4ZzYeXPN8hqKTK1jlj1vG7C6O
0+XTgEwtSAqR1FPX0MGgM0mbOB3VxyiBdM+37uUmBL7z4levT7wlq1Clz/jxg6Q+hiIsdHdoqkUg
/iyYcpKzElyum86cUTgc7jn2pzT8QZNBVM8UwfN9zbKnaVMB62JOUIdCoyBnEfzHvrhm/cVaMYdU
EI8T6t/phzuKP5zFSQrYmbygMZ871Au3AScsFZ3v+89x+iwby7RQL0I1mqi9ULJ8WvU94hIDL+kQ
Ld7LqBRAeFhT1EIJkdgP0I9PaNjLO3n+taYnqt2YdaF0faXGGRuvmsf8U8SdViZbTcMxA8i4Qvoh
vvgnDM+mFTLYovE6yET6XxFaeV/Ke2Sxyd2tg96+UN6tcf3XT9LXVhJb2w4Ok6VOcwrYQD1qglA7
fq4LsXZlOdy01ARD2Vhvp4qqXdtPj1+9k4H1MAd8ghbfR86UxLVMrnK0+70TNB/2GQjssAaDaYsS
BSx1I3tzj91+k7kNKIZqJ/0s8bY3yNJ5mH4Vj+QqWV9Np0NRPRIO8+KEPB5i+gRStmH7mJxdL87d
jbMXHIdf/wLQOXqCwuea+bYTr3KcJ9rV95mISg61nYbUyZuhmhW8CT1srVNZEr/Cm/59dbwGCO/U
AoWWeSAop17JtkPt3YhBN1KzCC+KiRqyKyqeB8ONFqPGbiEicCGVHM7obIMROTcfUJ0Pi8E09ZQF
OJ2J9kAL9fwpZepF/PkSWnDkykcTKTi6jGoyCwvYwYxcyxbojMbnTgfCuRWhx18yL9U62h4rLpUK
n106KeXA26sMgdI3fLn1GkZGyV09KHm78+25mkMKT9++I3N/ZxBk2McLMarcQyBeGYfTt6tt582I
e1wt6PmLzvKe5HWVS7w2uf84fNNBH1fWRjf5STN3MD4wTy7tJhdpB+fUoz5Z6kIv9L8Oj4K5UUIH
dntFO1HuKim0GWZGSLzKeIJc9iYfH/Ye0TQMFs3QdwkBMIf6Zy+sOHDYbcepEIcb9FTbXy+Tzqbr
4LVWWImU3yErbP5nR/ZnYi3hvmgvo69f8HLb5n2c8poO03bHolgXqkw50djFvthpWFJd6XSFWwyx
XWEIpo5f2wx60Fva1UqhZSyDvxFDGsTVWoCa/1yYpBdDkf+udctD0wNeWsU0Ya05VEQO8uwdBccQ
mwQ4lCpGkA7aqXmZDpIByASDiO4+J/5/ZFDZusWGPcrE4u/lF0QfuLOuicERdDfbpOjbHtbVl6vp
67//rVApf4xl/xKJddOnUNT1veXFaNHaraySK6p/R+MzEa+XmjclA7VmfYICU0q8sTHH39ovwXI9
x3KQn1bCs4Gn1KYjZi1pzYmZn2ywB17mF6QK6IxpiapMXMBxDEDL+suuTJoE0UXF2dR8fBtXwkcJ
BYz0U3dInrTw7kuOOsPgpQ2vkJ9HQAyAWQ9239OAnBAhJNyAQGnc8FqLmQjXh2VHEn1z3F5eP5jl
gL09YTyn4pxyhZjp0C6lJWpNxFdmopcBaLGpQWCH7mJb4Dz4HMXIz0Fmcw6DLxIZYo4jERvuTLt0
dUhJR79cFaAAyaBFIkQmzOW2vPkSMitFDNO20UdDYxHra7yIZwe4ArG7ssDhBhXVilfDiFGrsSHe
gYq22GO5+3CGsn3ycxT9xw2gQ+YFfWhApakQ5ahjD8GjL0VjGXrq8y26mkwmmCkyP2VVUfwG3yOw
n8F8FST3MUuJVxKNJUNWeiX7XWTav9tmMGL1evhXIFdUrMHmwUOpi3i0yB3ZHdv9NGnPoT/oaliz
iOX72L4dKcBX5Nh61ZjuuYmk5AEiBAOtz36+iFYUOS/BwOVHbQtgJgEMyq4JT7R38VXIZX8uI9Lj
GcdTbMSvo47jOToFhSf14nFzUzt1dXeQhHG7RSxfdQo1t0aCm2owlY9kBmSSQkM59vBL0VpQNblf
FuZk0JjUA3YZ9l7VlaVH4R7pvwxgTUkilyOS2EOYbkbnmekRqX3e+FAYJ4/jJGH5WfDkzFs3qFB8
UVTS5eh1QX8WCh2Ohp3Jbmn2TojdDky7LPHvEDu3MKhbrLdfWU+pJVx9Yut4CxJ9xiomyYk68+wF
aQrRGeb2ShpjzSWJYcjuv8gwRopkh73Q4mq5dXzk9OBAINTPrnv2NiTCxZG4SkkvU1wKXjZlJ9oQ
WjKTE6wPsiEHAlXCfkp2Gfug13z7Oc3m0qTQkt7hV0B9KYRSoOuPHbjrqZHqZlpINEwTS0PO5D8+
hZAKCRSPqtLJu4EVCVIlP3vnyA7GYATBW93T2DSx+tsuimbXOdbndglM8Ot4/40grx0OLJyUWHFA
s3vBPSDeM8Fdwgh+a6jy8pK1KTYNhxcgnJQm+GChWLI4O0C0o0ogOahgUmSyW07xbeUdcxDXODIG
L6idXg12AlnNGBdGMfcYoKODeI1ZrkcR9H3sbvykvgGpfpl+RKBmVKxwlOnSEKe5dlPlDSiZZIZ3
33iZkAAqmHwbM7SlnXctCZ5Vn8QpnoC4spNxwngjpaUbkMe3OwX/O+EVNDqpgGyRtq6HSxm5xr2a
HE6GJJ3dD37AzFXf2N84OsS0c+r+l1C9us3Y+hIkVEpro6qodu+D/bD+lGkHwrEXTbvU/xOhiXMy
DRgQooRb5CJ8knJB/hiHV7/w7/lNPJ8TLBPqjSm4C2ZO2H+FaNnPRKBX1XoPpmeW1R3arMV8ZGf+
GW/micuzLm/c4QVYqF22VV90YCjG74wpxED325HzX349vhrPUM0sN+BHMwjjCSy6JlPlZLEqiUz3
f+vHO9CW2hKYfBThE5CP+kQvBxKaHyAQWcYKYwqnMsqJtSCINlh/isQ+Uf856XdiZWeIzb/c/z3e
cKydn3hwo23xPcBFS9jdN7q+q+O9kD6RhgOtl5pZwjwKWIbG4p3gqgoHZ3jzuMGi9Vp/EgX2pkoD
GaYWr7hJk4INSejyFXUsAg3mDJNdvppL/PX4PfmieMeFW/UsNcga3qTGzB/Ey3GxZ3X4RqJcXFtP
LifAhPN/iXferlPrIWCNMyZORumTNWfAeVOUYizpmmc2k3mxCKa02dg/3fu7S8Ujyc/10SiU2kAj
E1eArzf4fSy0SfpJv+WIqDNoosLqN0eBQ7H6/oz7siLi2nSpP1Y29vcL+/EPLSvXsvHu7nvu+j0y
MUckhD6bGkcMu2vtb3ikTRAkl3oGc+oWk5yd99w33KxwhfLunNAf8VAT+4jJp/Yqx2DBXANoGyqA
9uJ3qm3phmlCyyeWqMcgeAWFvbJmWbo5ier7v3iNnAa7MaCU5Re+DkWwLfG/eaYG44XbJ9kfdTKt
fIl61pTG6/ByAdWjeEImqIG8VRV0MQCsc5V63OJOkrPif8MpCRuAxgVRIMUhgK+gB4Ks6sjx4+1U
ayESkPqrRUf3NfOYpFj1QUHQGUm7adgo2oyMABvVlgCGYKScrnibu/2lO4k2/RHs+8UlROhqJGrX
fjBPIhjDNINMM1sVa2tWRJs8YRE5T/S3cBhnUMRKiweoliyLh0c8OSYpz37PljDTKbRKnSEslLvE
8zUZzInfyDcgHPq0Ie/S7bf58grXYcB6FMw0o285vGlMhBjdWynM67AVdQaVz+DIkg76sHWIGDIa
mXAlYIRx1U2nFBcPeDMcUmijRIHL8aNzYaROWW07yAA8+vhhf7Wg8wvvafUzXw98kAcWeSiQBshT
oRhX3qiRoPuNnVnMwa56grk4cUqCi1p28n/2kkMsaFR2E8KwQAhWXSs3kDS3bvqeouveqpTky3wQ
jOHvRCaDRgQdTlL9Ejxrh+43xuTeKmKk0BJdLiLD5En+yMi7vNrWmTuSA8K8/+9Vht5T7iDJpJXm
LqGT3iQMhIXLWlh5uOLwMuKVnEZhChS7bP9sZ6hj8ShDAeXqKxObN+DOhyOLSuj2R0+pWVkG3rqx
W/7MM0rbYsHVxsOE1ANAAMh+mWIC8TZmsuoEHUzzkkXe0heRx/cFHbm81eMaJ8EXUmz1uc5S9UyH
ebPeZjlDsIO7HW95a9kBMNSVZh7No0Nxj/pFkTPxgp6vqFUL2QGP+fIEojtqoGRzHCNj9iW8JR8q
tQkFK8kjqbZ5IDnyk3bkukzCrW2+6zA5EItfsNsHli75rzzfq0UCJngL8qr6CrytI0Q5kIadLj6S
JEGu9w0XVuEbI7hp8DKdVRlRk523EFaq1RpNh1KryK03UejsgOPXRVk1qMboh0XztYwktFQLnMaw
S7DabJKJG5s5skZgiD5QHkeRp5IBFCQDAHVv1Ytayk/3XH+woxdYza637JxyPor9Ggbi0C0jvrQV
/218b9wZ5hp81QGE8al3QzyZRRHixfUpKr/Lk3gWG6fzkLCsv+0ayTKRZlg97dkHpmjUZ9VkihSx
NIuG0gu6ULEG+0+U0i+Yo+R4yPbtlbfuoC6GGRndRHCDkEusMAgj6kMyer/40fXNSS6WXAgTbHxR
UpSiUBqlU/aGhvOBMeBvUjvUOtDJuK2gYIL0XbbqL4u1xEYHyjWgW5bxDWATLpd2osCaqJMmSIO7
LOOnth8QcxwrdsrLxy335f23jYnEkoYMb4wCYTjVfNDIo4SyvWaWnwVtCIGrPd+PXOuzxI8jzWi7
PPMxGiDpGX0G/pTbfgesAP3nf3U70UStltt6a8NQNkPPXPNgYaUgWREreXTBBVdGveB45AyljFo8
0SkpvzlGsD9vSAqSB4NFSlVo+a4R7xniZGIFN3tp9QiSVCBZMSuU0IsgcHOw+QIehkeeF7nALWBb
hrlns0XN27ai5FSYd9YMjZ2Ov0w3ktdSkT+IL1jqzywiBvZiduVquNl+IgfCpAGubtDH+NEWMnoJ
71fZiaYDi6LPRk6xtdOpcNVpxJim13gXQOlnbdy66yR2jRjyOHCpeGZ7ywFgjmI+9gO2dSjRmCVd
8rNrDE6rtnDVrV4plHC7FAyg8ElfiTkV0PK7ebjclWCQUuAitLQ1k1gWyXfraALMCtPXQBVF8773
0fA7wnAu2rCGYVZyoweT5LK6R5/dNjE4DZQPkpKer3ioOy9f+5bjxFUxAKXyu0iX3c7E+9Fw7m8N
OGfFvapJ3cx8i1lykK+e2KYK1iQkQv/iKnWC3O0EstTn149rC9Nb/lgY2jT2qI1wjujIdwRBCF3B
R009tPRmhOYSL0LUoU518FbntmJkbHPt+qfRbru0qTNoYNpE+8MCDFcQaYmdOx5OkeJYsNCa3vPe
hoXP7j9lVVW6ThSY1VMj3aSEbqJhawXL84v/qus1m9ijPkdqYlsNmPGAZjUhWy+jw0ShqTAZsXlz
V0B9RJjgFKPgCMyoud1aUAcC/N4HOjg4y8ATDtliRsaml3BA4Oz0OWQGumS0TfV2fW7mczTKJ0ww
jEyR+3XGTZdcwkfrUvpw5RQx4/tJfMmyDG/adYqBGKmmFghA6cy2jJngnFhV4AmX8EDzwNkxaute
rvLl10DtXMqwGet4nCrL5bL70YW0Cbdy9KY9DhseMoqpEN8GzQRN0C3n+wlaML5qX/BU2/zPUUGk
ws45n1Nf53ueOZxIIbxqtDr7/VPfPGu8apd5DFJCj4xQwX8ni3Iutc1wBmwXTcmMT1uRJg+00OTU
gQL6Wc+PNYG6rLObtVPOArp+bw+45yrt0kzo0uT1ZnbHrCGhB8KNA+UlSWbrYek+Hxs5i4wi6Gi7
rnojkadd6/ohjBh3dnLBv1IIPFinLHNyUVWVfr+QUlySEz260hwiCRWr2smp4AwdAk0Zdj4plj/L
m4L0L3aAOB4Fc8oW/j1HbzRnVAaJ38DiVePXjNLZTzy3jGAHHMNZCA5/E+6TULeff6kLsy7W0XKD
aJVdtBdiFTASlPRvkGgkt8IdRZ/EIJDwD09HVv9g91pyUEAa4ef8OQikmOI4Od8ErL/S3AEq412W
0Boj84/ClAzzu9nY4Qc2PbzBNyJSu4uaLbxYrBdKCeQ+nj3n77+/5o1JhCjZNCAQn0IgQxTF71Ke
wZ5S1UuehJfRXc4NLGf5DRDm2LipKtG/ZMdLRs3dkXtLPlQ+6d0aqtNM9hAE97dGYofsWXzlLTVo
6M3+ZiBijM2jkRGblZN/qFVhzJPyCHXxlFVBNQuvcCLJpmzno1Ia52i4IksBdGjopMeDIKsxAdA0
8HDtgIysAUAcU0Q5sVDBkwMdT5qAyAufSQfVd6iAgyI9O+O0y0JwKz949b+5RUwf4yGwXgM+mTf0
SCRXRhFy0tZeefMtLoC4PJsHeC1jkfZcyKIACJUZ3c6frtTQEUNMGU6dyGiwPROu+ta2BQ0dtBom
Q/8tlyNGaDWR9g1bdj8JTP+k5+sjtF6/AMrJaJmqL3J48C1W5np8HtKIU2/1izH4hf+hEXy/ZIKf
LCeU9KpuCrkZhnkidw63LyKhGU5MyBQOEZtYK5N7c7ejpFtsj/kcHfMWZMbqCb1GB59e6YzXXoRG
cNMr8eSoc/Bxko3J9W+mpGVUfPBL+EzJ7f6wNSHujUBh/6D3m0JBSuFxijcsioGkONXPfs6s27iq
j9uL8ieYV7JzFjZnUom0JyewLsHCm/grHi6NPPKjry67DNz25k9q+Kbt8Xbp2gcRrvk/k8Y+UIyO
Xt78fwlNtbpkPrm53muK69N1WoeruCn9HvUnjP8I96SC9ukwFiIGCSFDBiZdN8e3E38r5++e6huJ
G4mWnxJJM2mHLgGm3hBR/IjYLb/oXuv+WVuxQzxb0il6Zf5ymPePmUMXLoUkMcvap9JfWt6Dp3o5
RaqHS0OBGQCop6blo8Sm14eTJ1bwLeUKvmpq3aIF3/hEAdYUxLA+8KWMELYw1Nqw2jKci9EOzYdL
WRVC13ipdWYuRa3kgaJsRWZIXJwe3WSGigYU9zWp6SVjxnyqKZL+9VJPySAISAerRLO3Z9O1Gt2d
4CAdzO0SyUBb27wMPd8WXM9SSLr/7jLs2c/z39T3YueSxoiaoz3xygDVAajqCKdl8gmd7Xs8bk1F
0h5LbHhT8FnzWtrInksgh1ZtYHo9HPrQloObBv9x0YtFMIJrElEKM7GS2cZLf1vMCCxQ29doK7fB
dzV6b+ET5/v1Kx7sj/rO6TJ3YiUkEQcADS1kDKVTdtNwGEFjAYTUZkjSH0OygpNfjazO+eYE0WAB
uDtgE3loaRd2oOUFAUQjWlgjAREnBCrv7xp9MmycxCc5jHhoqCyIpQhQXOow3HhLTek/AJ5IWQ3h
boriAcL58Qe0Sl7C3x66ncf35+aKyfxElXNcU+eb87aFg+tljUk+KYsZCq4dcuKMyXdf4TdUwQWw
RKXGk7AFVjIXI6ZeHuvml8EIR87kNRHPdVJHAYBXI6yoefDDvG+rWir35Mvqu+YvlsWiYg6+1Pha
XwxHcSQwtG66F4/2kG5K80cylZqhByPOZ/qoohtVSPZsi3huntvng/cigzaQkKBR1S+vLIVWoseW
N0aS3z9YYcyAcCXnCkgQ8HTuj6IsBML77/ulY472yoebXtWCf0Ka5/wyXiQnHaCyzJ/BHF/pIFof
3vCI1SOzjYgLF4cbYSebFL172pZLPRED61UPcLLrECEIET3xoBkkRiNO5QH8UPFJw0qkG9vMbAG5
dJ6ctoEdkC/Lff5cLPmTAra3LZXvMr2D654h46xnDQLw1wojGr7J1ysxJQLWzbDhhtBqPC/YqhAc
VOAWapN0UX9HB8VK7vTNLYgW+q6xT4BR7opnxyDOI66jxn+7wMof0NhnhktHzK20VQN3IUjCR06F
gZ73LChViLtTyJ0hL7B3gu5SG+6Y+ZNLAHq8brRu2Op5YY+u2Ixif8HkAf5a2b3GwYOcovFVd+3/
NAlSEWRblwB3Hdn/dSvIk2aYf3Ukp0RxmrJWIPEV90J5qs0WOJD5CGExzDMM4Z3ArWLg/pqcKw1j
t8AvQKX3Kw19/o74KWqAo4qH0STyw/YNv7BxVcxlx4fTnlRpwzpgHj7WzkuV0ZmzDS5n83bsFSXm
jvlJoqrJWJHgdFCR4y6qlrMGpYymHqbost0hVz0phV6+TGHvutXRu+MKrpRe48FK1u9qeGZm/sAH
TKPJmemIPFfj28X2YQ2j82PRuhxSKPFc9ErtraHPvbpjjRR/MErgMgq/X6o93GcDjqEADKfirerb
8HeQ5Qy9qZqFLx3b/Q6xxxuvmXt9sh9KuuvP8hHwmATVFQXYzMUbRxfo+DYpaz4e7scS5SimSZkN
ZTm9B8lp9JlJLRFWvg0loMMYdDITNSJXzcaro3H1sKD+J/4UAjAv7pcW07Jia9EOQQCu75XZSH1s
5Ar+ZW/aApN4imKQ/EVcufih43UWdYtIbzNjJKL32fjTf3142lj5tMs1B7MuxBlPW1pXOS5lnjvG
h6VjsTAoAZNplH7srIMGxdRePctKCrNSE2lRzxo4nTdbOuDShRfE4lJSgawf76C8IIpgiTuN5Jxg
voFda6er9kKzppsRupGUtjwrs1EwiNOo6uqE3ZAa2O3ohCuv70bQprupnO5KfWW/zPk8bFIBqdSd
J1simkmPYTzM0qHWprRNkQtP4zYR8xnRBbLA42HOsQZPyPRycMz1MFCde5C35n/2PnGR+O0BmVfF
7jvMIEwYA8fTw0hbnEoIvuCWOLKIFjPVLpsaxSH4+x6ptMRu3tAdFmWa0z/5Frv6fHMZfXf4gdJV
nPl9BjppITX2Fg8CRiwXEg8w6OS2ZZ62pLmwLlsJCE/7JWXw5hOdJaiwLC+/6451D5huO16HV9xl
nUuvGXomO/dxWv3cchp6zFW5YbykjM3LYcQ3tb8sXQGMUm17PzxEGAHkPbpghB+d+xFVg+Q+hS4T
zspoL66WAghr+LvCPpSKr1cXzWkSMiUyBP6DOyNqKwUpU4ZPhZuFrP0NzL0P5lbdtl0TGF1/fAN4
2eCsBEllNWPdQ+8cX4KTdsn/RyNOXmbVteirsasnO68IsPjTKsR6WipERkSpM9BDdn5BLP5ZSge2
MOXjlLWr6J0Cu00LX1KGsgKRZt9rRnsv5BirItSYeYvhkw2Cv4jhWm6MBPVKUnhs8ZDoJk96un5M
AGnvxPuZSiy/ZZgwFL//T/B6YAQI2/JRoDZCxFhCata68UWQNoSFiYaN2Xm2vIHN+boEDJnSau7S
QsCqb/TGs/yyzHuWAo5stM/toKwWIiXGKVXbPwwHGZ8bIM2c63XAxYc1eOxEWJS5axVFTODP8Ypp
0xBA6QmeLPcA/t474d5QGInqhAnNxG3ZVD6J/oR14Sd+3N2uKYY2NmOc9Kafo1PVbISJ8X5UtzrO
uKC035QSvr00b5+wRZUkwkzAWN9dOekkDzF5rGoi5A0v/CK+KWYMH8Z/6xKhuMxmAuztyy9eiIkp
FkiTmaRCj+jFIAHFu/jjyC6/2I7xR8AcuZUOZ64LyS852xEeq5cs9Y2AhwHZ3lyvfCB28JMbZxrG
1zo2Jlvvz388Abqyp956wpFPPtaGSvRxvFEvFy0qBioO6tMuWf7nt7q4sg9HbqZOllXbKOWY2Dq7
bjf7PTHPDiZrsuPCYty1dIj2xTc8meVrVqLOA52HOFpD8awGQY2IGyuFBo3Fe6RBpoj7KX42ySv8
3CnQOhhI1/I6vltrvCBAqGSUnLjrqJhU3s5NOQCYi363IlNdZtG1R9tGLyWPlfSEDPSMPFZVhZ13
6pR15pCl161vJs/xDz5+wExPgDCG2eiGcvKnGkQeJqfsQ1QPiKrqZRAn+fjkb1QtpM9/2yn3raiy
zD25nbtvMzrm9mZBy+T16i5Dxzu+EtGuObhDYPPBz1syfXPUSYyS1QJDk51CJ3kazerta1QuisMS
dwYYUWM9COmaUnnyVxZEkqrvbAxb5hqUCymuAmq4GxUDNqaN22KIlh6suovM+oJcEhniYnNDjHTR
hDl4vmS/Vw0IIKH52W/d2rCplZ+NwR4eY2mKlQo5dlqY3lGq/IJtBn8YmW74auaGDGGNf5ogZUhq
Migtbq6pqPCpn0WUopd1fdhCONblA0aTmILegIL7oxHHp+3Qz1qsw4pA1eh2/kZRoo2Dc2LbqZfv
p2PqyuuVZt3/LVp0sE5THLpQ5xUzdMi7lLS4Ewwyp+3E9aVK04psvxAxGH8zctGPRWNxM9MGpAwI
JamcENRZ2ba7t5ekhL6o2/huyxtGc4jUe9s66ew/Mh17LbIt4BFl6oZTqO8LfnGtqstXWhRwbNmy
kzSnCE4Hwn2AbAbUX1kDDP/5iuENNKACT2DEeWmTUCYtSksahAkj7Mg08oxPb6WLs6QyrlYAyWjr
Bp0vmP4Q60QyjgfNMMMgtGVpdhAjemi7Wap1DL+BT3G0cSiQs3bYbRSm7NyNN1ObvjR8TYsPT+lt
cEcVPEGp3Gqy2cw+k315x+EWXhVumE2B5lW9BdYExJW1OmFi55wY4pOgdxLLVQeR8hWy+KYDkclS
nkKZQOQv2eG2ZiulJENan1ckE65xHKR7GES1vL5TvEv8vfOcUK0povea4NA4ggBUCXWUO3eipMMA
2Q0TV4R0cTX76/xJJ/MG0XkBTP/hswJd6VEUXLotwe5eZlFWJ7OpKEgjHAv0EqDEo8AqEWH4SMgI
U4Qw6oqenYxPhIzwpd/UV/EQMl26s7eopnmsEwLVMp/mDvobi2OxMTPJbWZdANPCrK7ldzjGAGSN
o3q9OEVQqmgy13sSEV5oKYS9jVQeGFpWIdFV9aWLSCnOkwaeOFcSnQlCqLUGky9ExoUKeF22K/sB
6h00W7qZdSnBGg23mANl0ZzP4hWVf6pXhWoLs4gimHTAm5Vm/BGo7ZfFAB/Mo/DnaLlEUOTF8ejA
I8K6w5IQF3c84nbt3Fg/g2X6Ef3Ocqw9A8GaKepn6Ibc2K6TgoEoWUIUn/J+gd3iMpRASGgLGADI
0C/23eE1WvZ4ObH+cFPaP78FopufVw+VEMnXPQ9KVgdsmcp5XvNF4y5nNaKAMTT0Af9MDfeeQIG3
6Mr7GyG/5UWHCRj19M+6ujfaawowzwo+DPjnUrNd1ybIBkks9xy6UkFyQ1+ZZzyJezR0DuwZ2Vt3
1j1x1YLi7Zl4etELl5BXLUm1ZGew/A5Flju9DYnI+WPoL5xaMw2z3MD2MD0R1tBz3e3YbDcKziGs
dEH8OteH61tfSCfZhdJnKfhIh/IPC9YxzaCNJ2EL9/2WaoeOP5PRyoIdsY/b+1b3aocDL4t2SIAu
xLSXUTol0GbTGKmhjoJ/LKnLIVdm+X5GftRs2ZdwT8lfIAyHvvrMEswBdhXUOgMau/m43ZuodVa9
j2Fbp3xBz9d4c5qCVAmP+wuT99qheVzk+urkuYi6bef/BQ71PySSLTqJqonaAqvfazzI5ehoHrFP
CbQw2dx8adM2ObuxHKx1aW5sgA3S1WBZUV5JG5yt69xsgCY5+VEpmOZXyLsNQuP4r5vAcRAJ6hbj
BUkwTSAKaDS/M5+3Qk4M2kGDgWP/5NqNPosfdZNiYGoDKA4O/5TN+yhwHJM6pyvGpsdCUVNRmJfT
OFBF0OCg+XnOHOp29mjCB58Fyd4ozhSs5cwFFTt2yrgkSSQwYFdo90cfbp2mZGNLGGYAmSjI5Sr4
VQyavQbByRJjGskSBsnP8UVLePSNN18FjddW4kZXWGJkRf5TcBtVeAPYGnGsDusb9xw2rau7DG98
+OJJT4Pxu5JtyfukAFF3mt8de14gdFzv2A3CL9joseJ3BSjKqx7LQR/BIuyEiKH5fRwiRZ29wJb7
Wl54PKWzqS8uZhMLbMmBitq4uNkZeH1gYOVS2dQqutXFEpR7sUvDpw4wH4YzUpby6LDTd8K24/AB
ck5usTsT2KBWqk0XnNMTy7h+7jk5t/cay5iXfv3D7DJ/cGGqHibgmHbmJytZfNoqlWAnIr4fftKd
wQ/SQa/i0h4FiWIa4Vx76beqt0NAwyx5tIgXI/xlv017QE3R0oH7MeLhFM586WM8+ZOAyroPS4mN
2hGcKuw5fe8L7S+n5QrGjwa2dDjUkiOZj6gyNhwiAIO89HqRy3ok9MxpxreNLC2CPku9hyO/tPoT
yHCazv4PNobajwycrYbSodGqFwJHoxJjyqdiXjM9znPBFiRoFS9+pBxg92E0udrCKUw88ru9grGZ
WePANtC4uESs4bh1SBc7pYFpdvTLkWJ0q7S5tqROIr608+YpOdXu+de5exBHlW0V6fzBm5Qubn0y
YZZu+heAH7tuvbfyzQ8b3BuIcZgIdNrgtxffeFA/bFNcZYfPyiIgRAiwaVcwKY8groPB4oA0CSGM
0JBv3yZfYCsNAWoL9VCM1XHi0MCUJEKQM6kzPAeMgP+SLIduF74YGkDqIk9YpagLCc2HTKNgdAGK
OuzXCw+cIbz2JiDUrwDaJzrgLMWqtZi5ewLml8fNfdORJgLvavDqwqDP3qRTGfn6/rSxbmGUjiwQ
SJcZ+7uM8hnU8KKHnn6BdpTX6S+FEU22PL8cWJJOpvEeeYhr11BKK11GG2gy6Lj6nnmAdfo9UDNv
CdGFyXXJrIHaPy5tN0uvBouKtlRXug1+o84FE/0A4wa7Yau92vcMwq5yNWJAtyfmG9HAyBz5ablH
FcBQZAKcD37Rm3+z+x8DINMDKUVWwSFD8IoCzMYFl3yNoTL6O4tMw9KWfjSCXKS8jSvEVL9Kknne
+FVAvnzZ9U1IYmnJtCAr9GxSEkdUy8JtRqlH1Dv7eSd1XDH/s9S59pd52d0zNwA6vJmRlgGpLzAr
7vvNKafsfaDGYfAbUoq4AkCyq4OhC+Iapqy05KloYsW4GXiUU5/XIziBihqeHs3tEQKsRD4baAig
tdEGk31uUb2ARaZeiRAa5kpjxnjxmrAAC1VfgYEmhoDgiNzjE6TBLUtzvBJDGreV51Paj+C6Mimd
AfCkl6jGkVi+w2nXPx1c2xpDMwDrOL6r/9qiMN5uWA9N/jx5gsmUKTcPx3oTbMJE9sNmbFdsk4VN
b0VppfqbqAhsswmvhjFKPOrXkD6iiJLwFUKMWSoaMFAK7uwMXw2rGQYBQesRbJezHTcS/z4BHsNv
VjGRjpDvb13RHDEuIdt/4wNUviv4wgfUewrIKgcpqYdASkl6LqipGbkVRp3TH4ZqVHIWpZhYuA9y
fFi9EIvzyCQxQ4QyOFEuw8W9whvAIBqZPMF7WJXVklu/yd7yL5PWqqJ18DjhsjSrfChX7TmYfhFc
5TdNwfzZ7n7hpu3aKHU7Mj5DOA44KinzLWeE5XiT0MjngAXcEriqXN9K9CD3FU3aDXhkmmDuDGOL
ywejBIhTRDoKMcrO6dJ8q4DKzBTvOCSPjsRj9zxaw/XYj8IftwFUuvdONxdmn0qUqLhdqw7BxonK
uVg113L2rpYSuLOa8JEdSOpIvwJNBela9eq0kc0PaW2iyLT552m8asDuA30W+7pM+glsfqtYB4BA
jnTPOJejGCh/2xQBXOq8RAtPi9DXOc/maLAs8XyyujtoGjyFvdoed/pBHqTZSIJLwLECyXIkJVe/
yUWxoZsw0u1ETph2NPxUMqaKRMX8vQmvCZDuW7EInwagTE5FbyrSb+M8gJBH7TQnV/UzoEgqGYsg
FspY0/JSgsFNPDshWb/ubakJ1eY6qvxaBUmzjI6+ZbvoO7wimoQBkmdh3icAjPsL2UMQ8O/pGGlg
ufrsETOSXdvZB5Oft8IwFvHFAZkm7irtJc/E3MlMtI5/KdGMG+b/D7HQKK6c0NJCbRXYlj8rZAMv
v2CWhKGkjlc5xNZw8czcgRyjh781hnE5Bhf/zyRw/EJY7vGnO8ZdiSrBGd7lokD1jZwVvEuqIuHH
rZ2fB3Qkm7pKGjVFoamqywGULqG6mTmDUOsWcNeFHZJePENASCdmWzi6dMnKIGR/q8sUVbyaIWvC
/CeCeJ7puXLuz2WHX8QZP5Y6zVG45Ehd16r+IQHljHlNK+5OD8LwjCCEqnsS9nHydAPv5/FNtgK4
HM8ImDdOV+ZldaTYU8EYZOIOM1RCZ99ZOrZepqoKQkupM+2JwftwEiYFb85fYs0aBu5BTMZkPR7b
WKi1HBNTjAsfm/SRA04C9Fyla8FcFEo2M2UhQunXm4mc3/fmUhewJvIk3T6SUNuNNG42cVp9ozom
yIGbzSNM0GOGWotO89PjfejyRtDshIpT/VtwWStwEHVyVsgWsF5HB+3yBT6DJ8EB0tE4eb+thEvg
M/zYj7yJXhdj2bZ41sc2FyYg91xqrrr22x7NNIgdduZVHHIzuO3g2njrfLssdbMhoZCV1lL94jlD
gDx8HfzSraE65bu9kTAviXhK3vHtdgWt/pEFB9tNG+7ANYG6zW6sVkKoiZmYY9VS5nr17TGrQpTj
PulA4FVR0MHw7PI/tgAsjxCu7yv/fj8cd5oG7zINM6ynqYh0JzJoMYqZv4SFtoSysop06C+nqGPP
P6e4DMZ/IVkjso+QEqmX6vWjspuZLLEfHL6EEx98uwP1XHYIJO4SwdCqznnI/R0zLI6EmapCVuUy
HnPt6nfsyI/eTexTs7/u3wxr9vHT9lcBltI4OgDzvPH3sag4XLfXrm71p7EDaGbQ/6ROBuxOCx2E
1nDuoz1S2bqcCsiH38tHnZs5hpzHTN6P1O7L7uP7FniDF3i64tBse+wX+a+JruL1P5WlwJ4+5ZlG
xJABJY2wjOLMqAcB0bzd3/7mfXbkn3KVdEPO8bikbap4snr6fB4Mz7XSr3WKZ41lnSNYhzL7MW8y
enfSpdR3f2mh8d6py26Q0vltDGVIk1PAKSBs3NV5ZHMcmtUvtjbKgB+mE+v4cZTQ7sgXOdmlp854
Efgg1Qpyk3RkTR9j7KEJk4gH4UT7wEFkD42C6ummY8KK+fERE+GKQRXDK5IA4wO1nrW4enMf6vAM
axRH97d5c1ViweRpGv7yFkr7AfO3i+B60t74oc07nSI7+d5hBJQ6k89M95pxG1SdleleGk+fo1vp
DOSj3S2qP0oW+2CpQwZwL0FHyY5xy+EZIynWtP97iqHwqhCDJfnD3xjenKRaqh3S48sL0KxC/qEb
MOdVk97d8z148DLh1V3IBs8ECqjY51l4HSgT49rvmq8K4fIfpywA1MU/bto2f/voP/GgKgdnRot8
h5DmMQ2bUjfi0ihKZo7S2UJVSKNdo+qDMfhmqINayam2QtlxklfZvQezQjN6mC57J41CZr2/+QfJ
K1sx0cWNI+NG/aYxaJvo+1tPbff7ppY602UL9wapKQqjbGlSnv5ux6AC3ZKPL7wfWcTzHsnrNrun
PxCbh0wwTd0Z/t3XMUqNzKxHrDWNUDakaKimyNCxyp/jpTPduzl7th1QQCrJTfXtxUoyFBVKXj2r
l6qXIh4zDuQmjWKz+u9s+WScodMLHcfanMXaPpegDmsqXeRN0S/G69soVpAmYfagAFoxWO2y0Hsj
rHtwVFQTgQtHhCJ1fO/5DdyiDqCYcNB4I3XMmM0a7G8plUXoHU8nCrYmIIXwGG7iGqSjiyqSt040
e8fiAB+lGMTIzHbwBSZv4+zknjzw3KncRkt/YYyi7uxTPThwQFlsfUTyC7bHpMI9m+Fm/JnK8Oiw
/5IKjpBRYSWWzqkXfKQd44l8QzipZKLHbOrGCLYweigNd28XFEH0MPTYDftz8hN4Q+wxJh4hcViQ
XCx6DztqXTurlO9B2yxFxdXesyl6iVxQ3smpnzYryu1QZs/80TnL0zofxpbWd1hXuo32wEK+Tj2G
HKwDjoEaKLz9rDRAOZ6VX3pblUXivtu4DbLX5MSyMylt5cMvH1ro5eYVEug3xZLcgA9GSktLwAn9
uGZl3fh48THuW/1FhMdTNakkYlUuOl7UzgTPEVCBms/omXXPRTg8sx4jtIzotvxgi+vxe2W1swlr
qySyTezdgzHTeDlip2QS8ur+zG11GlKcNwhW5t+s8VCL3rSTdFMZrtFL8kp6KbGe7n7qVtzQhync
TsY+6rW9U9/yA4I4GfBMS2T4+2srMkxIlen6NiiEfinLHIBB6cDgbmRO0IxYZeeFuLxKbO3gc09/
mZCSObh6AN0q9qtCIIIfiNMuOKAy7KsKy6LpRQMNE36WtF2T5rEg/coBe1Qmo3zDReETDa0G/TDl
y9wGfLBQJuXGgoO1JdhYrkpZtT9T60A9dqj6a3tpwE+R6kF7Y3toR5KqJfZOqEwnfc9drZ3y/C+d
LEYe1qeJDVVyDdVU7QRHERrAaWaqRJ5UgVY+L5UzTngYVlRBSCW06I33haeJe1RwQ5m2T1jF2pcl
KjfrbBtCJVSnzDbyyaE0dP0sPQelgavpESpddCt/9r3UhZLXs8lWxM8ILIRCd3sWQZBMmRHbFo6x
OizxlbeABLwabNmzobSrhueec1Umih3K/SKLNk8mGzGzsYhFh8KuD3DOvF9rpovDso2O19Hj5V++
PxydbKKmWt5iPyyKwEhDn/hN27Zn2X80kI0YI2XnfA2hKafK8HMS2hJ+yVEeM4ly6nrZigaV42J7
/TJRbpkXPRpgxc35MAb9eFebEIcuYktiv0TVWJXy1jdjlWtOiNV3N2RRfyel26E6PI0Rb2nn1DQK
A3XE1gWI09I/7S3XQZAOwY4oK0cVD2vjxnx2jBoT23tFKbPgOdSeWXTkXiZKYnokpDlyA71Wjo6P
Pbpg1TItHYoOuEsl3WS8bLxpyfezVRzXJrQD3THOgdzZdOaZeC7jOI6sQWBni/1VYPZe47U/X1pb
zxEbUQimMW6auHWCuOPys7JwgeHKHBOOWm3VGnUDdO7rcHN0uLIIgHFuKyIzy7+Oo7trsTLPuohz
q5pdc9GH1A9dHiVWvrE9WPHuVAHxajo8Hnes6cQVDwImoYAjH58MsJj59GkYsuKffwsVE8XY1sfK
HzQUL37BlIjXXSXPa3VhizGxynrL9JVDOQiDd8s3qcWxmsGmB28/j3jUEhhBmwtGx2oO6sb9PbTR
ImstCgZmnmG17NCL94zcDjSYxM3njY+H7D+YpMg3ClTNW8LOVHMWtGcFG7o7wbVZ1jjX5wo1F2qf
e3qOnrzUxck5NPetcdrtOmbwaXcYYN4dVtU9SyyVgYEenExnkdRO1wpx0hullymMRteMeJ7VEAb9
SyQE9NdEBlhYO2RYGmJMGJJLsLGE4yCOUJNaCeUjr15N/1BFagWVzEhqqUY7zOjdI7kEEdkRJP4z
R/Df+uhgkRs/GuJTAQAK42eS/7wmYKoQHFaNXur5fZf8yZzo7IhLaJplXQ0FVrENZCboqviyHoKV
+TtFJOGfrK2jlLT20Ha6vFSVHYlizWVs6iH3dgkinE978plJ+hMabHkB8wGtUXTPvc936qfsU3ix
/Q4TGGN+DXbLwFQAwpwigMKIZt+GrkwALfPwxbIkizxDZdn2Jxmtrj/Sv86tf00+UxLby7VNqPXq
FUkJQnJiG4mJ2tdAdSzij7jgSjfILf1OMJGDsPXWNwYCVl0gmJibg5g3PvCNFL2LSaAXEBSNn3Vz
KFK/x/tU6KSUfHuWG61ly7fT7m3XJw/tJHraXtn9Rc4JcjObM4We5ieOH2cXdxkpPJ/HrTOGgtGY
Uxy2If8Kvqm2lEue92L4eMFV+cuWDbemY/yPEdKzGQVLacs6V1Frf624Pv1HoI1Wii/FSFaMREC6
9DMJOvqaNuNbqq2KcAziyXoH/Jhs2Xv8xlmyLcF9Kc7w1UIGfwhVRdOkvxOWf5cjBJIb/DEJyfZS
pn+jgWrAihi8d+YrkvIE6AF3U5Fl/mupM/1rtX4vZ9hJjig98oC62XEgT+t5cHjh/0xZfQfxmuoQ
srCiP3JlsVQHE4C971h5DYUNIqbmN3s4NgdDd8pqhwdhYuJFp/H+2ygRrVzf4j0fOpteSNWGlvMi
Nx1aNlZMj5Xz2LQJO2+440es+yFxn0Uhb8CXW4udLFG1CN39C67mpho0X7h954MLIxOk1FM7yDA+
tEieiAAYKkE01DAzXKQqtOXR19LXaAvWJYkZvmsA30t0T5KtX7xRlWjhCnkUa+z6/jRiWEVY6S81
s9seZ8pLuZHfEvj+yjp/+pJwUVJu6owGyOsksWV0vO+UJKBA0ciyqBG+yO/s1iJI3RTsqIXd+xZ5
5b9FD0tVIhjIAluo8gz/C0OXDjMp8LBuynmnZKQhoNDwijfpE862jtMPQXoRP/21S6qFYdGqOv0x
HWi/spnqGFRoVlbmYNwbtz04AneGSpERBDSTZYN15mp2QvygyE6NMVRJLadxIsJHbjoGd4+wgq3N
Q57ngrIyxYDPKi079Ly+nGOW+uAF8ygp/IJWwyAF74GP/SsoFk7Hn5g2pxTZgItif1gGLplcG7e6
ojslNaqrgSi3Hczy9ExnY7/BlAEZ8zqrHrgoDANjiUCwkepDOjZoqRKmuHKAc3a1EiG6OlQp1t8x
ygU9QrjNZpaUPxe/a1zx4BpRm16avwXmqYQd0xcihgbSigC/Di6tvBmRmJMzLGGcZ9kkijvp1uZz
TsVMWxLwC5dlz6cju58WD1Q+MkPsBNktQhR9OD9eVq6el4SgM70bZ0B6Q0nI3XQ5pcfxJpMyrTat
zlDTA9TzgLZ2tj8N9wlLeCyH3WQBI1F2CyU9kIqOR406D00fxJQBWZQahgE+17TfnyAkTiB+q64X
skp7sMvthRFRF8MO4cgYFGhF5e0v2Voxz95KGooJzqCDVTBzPPYVZiNGYobKbuEi1cqZB7SSG/+L
J2GkH2u7yVQGlkbO34PDjFIVJu78v3FA8m1QcFBfcbP7paFQz8eUvpZOSJw9uaaxWYX4DYGaGDJv
CWuieTp/L8qQWMPu42bkRfL/j0AV078QNpsscodjRMGErnUaYr218j2f2h5dMXNM9e02if8MIY/q
GVffqe0E7cx0A8fjyj2qPhz3Aqr1b0oyfYWLQ0YPq2jdqro7xpOaiTnkWfxkxYX0jlXkUAu1ZKiB
2j01vzqVrZVJ2kK8Cmad0CeGZDloVSbCvtgBe1kTBDLL22Tki6Q0TH59PdpjEaJNNMnzvqbBj5O8
REaKoCS29KwYubMbYlAP7LypTFnSX9Z80hzNgPrYkQpS5efd9an//JJcuw5Zq+XFom8H2p2mvrVs
tMnpBCK7f6PGcRBJMBRndJ6hVawue1XyN2dD+XBBRtd2aH9peE5S6JPiMEHs5l4dIuYXDqpxp1Ht
eJ9ekjxNzmPIJaysunq0eG0ZF/o36nGcd8ZxSioCuq52GWkb8GdshmLyvzS7+IgEQgOqPDf5HNF9
E/H+oHsHNFK/12/ZygDzlOfoZa5G62ybuhc4QHbAAoKDu0UJQNXIb2gDQ/UvnttRNY7CqHKP/pGy
ocS7+esHIWFXpl/FHo7TRRbUauU+B3olML/U+iwdb5fdgq91ZrlLhVc7TYI9yIIg/kPG6DZ6AOcz
0VYrTZg5zz/6Mju5Euku8EGNwZt2hoSOzZJPvyackhKYS3l+8fdZQrIfbVjM10a5VxJaFVdubpRo
AmYu+71EucugmUMHkIDdgcAhkpXEMSpp2vzeq9n73gi0ZT7W0GOVnIcEAOyGK8Zi/JgWkjr/E0VB
zSd1YvKUXk0eSMZ8HzZ6faByvUaG0EXrNrN97edaQA5Fy72IeNE1a5b86UBstPXHZINTxQ6AA7XQ
YRsYL/6cnzC0YH12sS77Qbx85eU4nisk2uwIvOpVHNteCdBqwxFMZYK9G0T71nEA6zQHn5rCLuqf
Z50lAnyQUwk3HWq/kwqRe/G5p0LrXpEQKIWSRqgDPbx6WAfMhZv1duitwz3sqG7+pk4mG2RGz3JC
J/C9fY6PhQdqVpVKhREhdFMm0xHu47OpRo4Ta6wZ6gq5WPgArBxTqQCleD1Vn2loGnsMord3WCaI
PbdAceCx59s6r5A/aRIbsJ0DRMVrX1GW7NIupHnBnQtYdgYI2vB7Tp+fvtl7RCrwuwsIdJdsRRgo
Tc13SWG5rtd4JdLb0sAOcPpzNYjaG7c0uo6lsEAASJKkm8ZKV2L064o1+N+SgBdJ3uS9qSbctRBj
8l08JVFP8YevAotxvSNcJBN1c0H2ub1gFuSDFcsT6y3hq1ESXColvEEDI4bT7TfhodIUjLoZeigr
AMZW1rxDcOirftLd8LoFeMVwHQXK9DnDKHvPxMsC3227Nxc2XCg5YOhga10kKTjY89PE4Fj8urL2
z9RDIDhQKm+fXmhg7xOOwReDn/XtT7COeB0MN1LIlHaMNL9dSQzHmhE7L1GoaoIXYoHO4qdZ9JUw
dOzbHsysGgozULFaYUwF72tBQfMI6Q/4uMj68FzRm1r2LzSqKIyrX4ByRWfCwU+YGOXq4kc9dmRm
C9HH2yCQ/CitKrdTKsUGnGmpiSGnusjfXDfQpwGwQExgbbtN6IULDGoTtp8zhyfkbGvchxFmrOUV
johjaH6FSQ+QvVvnzgI33n1GL2kxvHuUNbJxfb9uJs51csJI8NG63U2Ac8iu8FyLImh5LZ0XcibX
4X43RToyVNUGqOYe60NEJD0ygImJKr1eOSLqCwa++zbE204QqveE0QCtGIuMdwm54JZLLIDxyBiD
Eqk4pCaRMCP/OEFTGHOKBojEDcHYPoGRbWzaGNxtDLBGUXo8abu+FrLTJo0E2g+NxK1+N0Klu1wZ
7whWX2RIeTaBpMBDGP4yM9qdyHltNyWgkJaTRC7X6RJLFkYJhzy/UprGRDlEK17wXNN1Z7PR2UBU
E0x2a2yEo2QfD+gJvvaQ6C8GxrNlr+53HwReZhfLg5wrNniLm6kqbLPgFFH8xmUHOj9RqKuCaIo7
/EsLSgpMVE5GFlpTBoEADCyi0FdM8o3GiiNNEdUUQzBi35m7yqW897ys1e1IGjGVp7QJUJLIp4W2
yBIzdc9JoNZqPbGQMGtHFr4UQeoc4jApSprVeThBn7ojW+Wsye/wbGGDV9yVjTLEPy0zPsq9XPGA
0JS+5FfeQF7YUz+tqJUXC/83GnWVg/vA8AAsdj7SVwh4+4oi1w3heFTLGEXdAFm+Tk3CCQ1uHf9c
zIwaBGp/nxc4iuyrnW0oxjAnetDgGkZ5c3YmlB+r5Q8w4GpkhrucAlowMMP+16vLGCJS1xSJfszy
5OeDuJ6f0wBvru1tXy3oddNxhqJPSJ65s9L0IS3S26yx/cTl8PmVS2H30eEvPi50/vhAZ7g86+9k
0kHaa9ndGc0ST25pygJSsiRxy14lb4G7zscYPDZ1hlRBxrpVeAnKGBfXe2RIFJWN5LyF66j6WAqq
T6w4u5LLLvcXV4So744q6RAljGE2v4Sh2Tu6AF8DfIHvJdgKm5MzMGPPtJ98YYSIip11RAj3xAl9
7uUrb973mpyqRWUXFSvAvaxd4I3LmPZ0ipmvkoV2zp2Bf3LOHI1XGmTt9y2wCf0k/sBQXFBZVmmS
p/5RHEVhEaN2SrxeTd9ulLOQ81geDV4hkiGGY9CSj/4SHFCb2DyT+UmLyq+Q/SpBftZJM6O5UuZh
UfHmJKAdMFvWvEWgKe7CbqFV9U3FVwoi4UiDpMrfsspY3OnyQpgelox9oDVQcaZZpz/3oeMumtdZ
pbsnDNfepVw32XA11P7DYVu8SewMUplZmN8M8woDm7Qwc3e+ZMD6X4t6eFo6ImM0fLUYsjZ6rXzX
lD16hUQf8t0hbF/G6jEJVAzc2N50B1id1NtYQdGT/EI6l4iCAFPqKCew9EQ8F9ilVhnlRoCIDNKX
/2bVhsRHxsWyps8T2WJkyv91lP4oGgqeW43Zx4YsPYYKxpkFswTvjJ/gVKkHFWMnO+EK7yZ0qp8R
lNxDsPGyHUhO6YTprkMjzp2eu9PVphXb+4h/qYwsfizGomY0ZBVpC+UsI4E6Hs7lJQsr+NahO/AB
0fDRZciubG4vD193eiqycZ7EoKsuPkzCqvcW5bRFLdNjSIGlPloOjn84smDjF8LivnGa8YFqpQ+H
nixpe/AYJ3NjGDDqufmqtZYEoLpWC/mkaNadlMdLF8hhKxsTFi9nIXbp9neUgNjIIECphS+j8bkJ
SRNwtotSH/fWLDH2ETzeWdHb0aRcUD9/G0eGZYmVpzULBPSH3omX10Pp7qDa3iCmkkaI5Wkl20WD
d+/2HvjEjKB82j01feAodZFFz7F77Wedjmxc9qiHn0EB5uPiCDnlN4oYjm3Fxlj+fsR6YlCtol1T
ZgQqOZWSUONy0+Zb4EFHi4qHAuek3b0tvG5vHz2hk9C6LrUutQwuXcI/jKUbyeqitqFRnJqB0DzR
NXss1eyPGzvhmabfBGGVTw/378eiTEep/A3ezS6ayrwrhazXh3ZJX9oMkHvpK3GV4MvwNQLtv2Kb
yoMPzGlvGg4+/h5RY6trAJje3k2f5V4SktHn/2e4ULXOmNdXh+QIxTSWZC0eaDSct2/rYOiUDdIg
MAkapEMdkVNhkAhPHKtEpWlJphWsLM32BMnCANUGnF3GN8o5r1rW6//66w0OhYgtewPXkmGfuen3
EcskZfLzAmdjP4y6Qd7ZP7bfmWWmOHHnBZqX3JL1gww4lc1qPtSippyNcjnjZOsXj6cygjaP5EGq
6LxempElxgwVIVm6rbi41HIgcM/tk4DNm8XflqGcfreAhD8HgOEtNRJC3M170eZyRDs2/6UN/NWQ
Ie6og53PcKJmox6n+pr3K8lGa5AqexLgTzL3c2L04aHzFOwPzo85X64MWtTeV1lgw1UMwX6CTGFc
YUnOy5fOcuaCd3nqdW2MrUeHqqXHKgH+Ne6Lo+CIrFtKHuKxcWpUhAxFt+9+I3BZIfYjU4Uesr6T
fvIamAPbszJ1uGgY28JQnMGPa4L+U2wbYnnFMjdLYM+LEeoxBb30ylMbbh5bMh5AmsyihFDVB4uU
od6hWX5Z1FwiWzRIfS7RMQSfACcrdxrHxV7DaFxkHkUh6F3ELyOostkh3wJO7RYjAxx4tDvPnidl
UAbtcQ9e4ukkJtNlYAJct4tj60CQBjMGow3o+gqHD9xvaZJmyWMr59skep/9BNSLn6YaIXz3gafh
pOZU50ddkIk51e7QgRpAF989MfFbEo2LOX+oEIKngtH28vTe13ZA86PF2QGoDXgpDEMUjVe8C5YJ
txIqGDLhUjuPFHecGr1MnXUha2m8jfZT6cxwJT/J1DoOlYj95c7lDBu/nvSYiL21+WNzMubw+2UO
CLu1yFXfQFaVxpAbVq+KvrzLJWQbuvcv1zy7IfgiiPCcHLPKqVbfv/eFpGMSbBVp+CoLjvWIpci6
ioBzlWcIf/UaUJZrOBgHXBel2W5F5vgPn9LOk2YHfoSOcYSM8TKhs9X+VBGp4MLRlfKiiFJkvMAP
KUhxaF8l/1E1/GduXK+y/JTPQ18uJAGxjzb2e8VvelfrZe44zozHaSvCN1VD0qfVKCEgHuj9yALV
vEnmaZWygeY39hfp3ZhOwvll9frEQjSGtsXsnqxLDGRdJMr1m9WcoH7ZB1wGk6+Fi1kxxrmwljB6
muLt8uGKUojsTCIK4ucD+DULWP9SHCSkaS+95AM1dz/IyfIs9Djfv/fQiYPgbSFKjNFL2ii33xLF
etoCjR1sRviNAJ5yzO2wZFKPj3zrWaY0iTYuyebHrCYK075mvk6NUfJ18dv3KifTPMRo52CGgocl
ItM2aSJ5i0lgK+Ifhw6a8FT9yR2/KW7PWBvrEvzktFkZNQS35cwEoyroO/EeBU6pZ38spQ4/DqD4
6TdaLHwQAn9GaMbtBm+5m/q7snOqjPMTWSdrJD/YMo584rEKWjJvd3Xki9KJiQn9p+yHFlYQ6Bri
LRJki+4TJDMazI8OTJhjmQKKAew8HcLGJZm8v04zeeSoFbp95lEzaxsEbb5QxKCYfO0bkAQRjsb0
oqDn66XZsUPvImSqtUC41uGqdSTxU4mxLZKbSlQ5eGI2GODeJqZ85a3HuZMOXcpQCYddfuzDgMqn
H/PbK4MYumVrnUZqkLO8cb3aNCDeQxY3dUJVK5C653R7GjT4KXtVlQL6bq14iyzOhETg2Ny68+3k
vhzrGrfj1IVUOcPPc+FWHDnT/V95l69eknN50xN1ONN4IdnDpX61tPFWNpMfnXobQmUJR4yOPj3n
Uak/kF3e6SNZkwGABBzrgwaUBzCZKTBQLcj6dduUs07d90w4mNEuR1OkKEZsds+XzorGNrU6CWEZ
9H+si1hjoYaohVasz20zix5x0sWeCtLrmUHMOiT0pSljRLrJlBgwunXDo9X7yITF9Ny2epgHNqPK
mf8ZeKipVr4lr4hibZv62QhFsFX1EK+YABCWCulYVlBu+esv6Xel8K9hQDf2JFtgU5WSKEvkV6vH
j1RFH54M2B2ZQLML/MzzLFZdptbtvQ1Qn74Gg4wKCL46V6XD7rR4bB8+bwdWLkFgtQHky7dFf/3u
M8xAM/Gs+H5BBZLSHz10UKUWNUMnPTYBmJrO02V46pSV2ch+tLqdLHv8rMQGlR50VuVR94BR0Nqb
djUFGpXTC8dEPaQAC/pQqdMRl7RtyGLjLbG1+bC/0N6IxirOcPJkdoPewQccaBflB90o8Qsn6Qu3
azj6rImReRMxh9yw5v3akBJw8wM4LFdcKYSpm6SjN8M3OEzBchcUhIAiDLQri89bs/MQ3ze8mMa7
LWmXAmegkDmy7zwSQJb7PvH1brE44pBXDMSrqqUMnRzpUEwYZZV/7OHsLU4SqeAnByFqr9jfJ+JM
oqo140ThOPv1WI1AaybM2yecI5AEpFnYQAzEIEK4++dCge+l5q5U1AXKCAoFLapQUNok2yG0H3J0
aaY691P5xfMojgRnBBh8azpGU/3g5Iy3LecQ6yfhAFt4IIcgFelM0p8A+yya7Y2t4g6X2K7GwT8Q
iMwfTomusjPuYpBU9ek7CbEICbdi0ngBZD2cHegyCNUbvxum+QkwNtreYOlqM3y4vqaoqf+tt4U0
x/8ZT4gp2J3DzmamkeaCQIPFdp0bDD0ps2GxJila0wmJYN5e1Llt2qsVOwKs0N+SoRD1zNaIJijk
SlP5szxhObBUSiWReU5XGu9DVtyNYRwdzDv4kiLFBPI/Z0fABFKVlQSjG1smwEJQU84g8JtlE0QG
i6hC6IizOXeTUMyPm7S4xTrXJqe+UyeiWKIKE5S1JnYjhaJclLEnh3ExjQD7RPjlyqccdNpew56B
tlaN1ftrb5+fQa5xyxAtb8lpPQcud4HadFum9TfVgMgZQK9DPAQiQSWW7btny6k9+DEN9Y9mzrru
LyffKhnGNwbhGiqKajlvcpumF52Dh1GNobfYOhfAL2ik8men3ObPtaZkK7agipD5hvD0vNv6iZbq
NpAhvJnWiXYyrbqSwGQWwvH1MBczUkmQjBOwq67yDy9U26FxcQ8W8OrB14Ztsmo3JL63DNW4FSE5
iDQncPssysBAtOSwgy1q7CtJ7/6U2feiBJyv53oQEzck0AKFYiRV2EQOm+g2I1a9YrIW+WKZiHgG
NRz5uEScbSOwZaIcEb91W+gAu9wbNzxquwsHUG9H+hEdWIP7tKJmOddAmMATZwSOjyuWr2Ha+lhr
uHt6EMWhajCDLWe+hIH7HYNJduE1kIWWOMnnmoEWMdcNyaZGPQvtm1nZaC2amIXHLyCQ9PixQQvX
PHiSPeNlnIRur5sjBXDwOWskPB3E3h54kbdfF3/QA0Zby/7j90jD8U0QypYr9sRBuKMcXWFb9K8a
NcumZw+Gfsx+RYY8uN/aD8a3Pybocf7mIw3s7VpvaCictLDizPQVM8NI8bYG1RcHr5DOunCfv8f6
8KPIL5rS3JNIuDMOGU5mPh3AIBf6ZXCqoldXzu/n0swnXO/G66JbUVMat0pDQhPdVnJXFjbHPzcl
0wQfTn+/zhFZayyPLT7adwJDg25vU5+hricfbuW+/df6mIoDpCLOPqSPHLGKmAddm9eb8uERC9nT
gDMFnPZFr/352Zm7c67C6RCCbGj8tMitvnKxKbnnfy1AyNrO28IATeBV53zXoqicks3NWpmLwFZZ
nzQnqacGj6TCW0rHyAmJrTV4nvVy8xDGvStEis2V2rMmoxgp3x81Nh75ZAtFY+IZfbAl54gRWq2x
BWLjt7KOvjtOd0bj466T4kuwDV2ZZxg8/24ZXeoE4G4FC25/d2ljLVx032b5hr6SRFgBetrmojnF
e+K52lMfSqMGBf66jxX85GVS/p9CliWo4ehMlPTFd1qV1XvClVFVoblzMWvPqYtortAc2/0EFx4k
CrnM/GzVv7eQVuEmek+Yau21YjHDtdQqqJXm8Eb6I5Xw4oc5uzPx1AQks/v0D1aqaAKiq9/DR52J
elyAkLv/V5t15rjPwDEcGT8mvUnIYEPOhgsLJEOLL0OsNMZh9Lyg9vpAX8uA46cAo3w7q1wdHolI
txXXAsXPdwLoxrTejyK50TVT2TqgoqXF7Q2In1nkgL8+8DMjlHcUYE/OGPxFZzOvVxqPpCjxxwtX
aDLDprsiWEy2t/9//7pj+euQUsQWGINnGd31h4HeyvQ2r/i5SUvPdCQjt3oFeUdXMsPcLPf6Iwwa
Z/QNOawbfECQGiMxymyexIA7+LK2Ib4cVs5avmszfpXAar3Gz98Vo77Eywy7frnEKjgN02pZ5ET1
4FlcgXpR5f8x3velv8Xq3kr6azSfxNLPae+eNfIYeL78O6wewkRDxKhMylAV6o6gZUe+lVSSgQEg
ffCcbfesYqqyktGyLHCZw3C3yOaU1WY2G/jYjV/w9kSmDFL9xDJDL3JEYLaLChOqlVZKzmU2FZ6L
CxqXCewziIikpJ3Y+EKomN3InXkcbQOIhOHWIyBXpYmnG41n/YHsPzsj+rRhTCKN99e/FOcEWHaM
DdzypIlz+0Q5Q+Us9avhQbxH0t8z20EFe/5FtCc6++GiHvLSGT31xBaqvra5medjCaVRNc6xXf/a
uoS70WP2Nv7JiBWn3Nt6zWeLnupOcAgOFy3+ZeikfYawdDUlAUryGw3mz6e94LWmi0Pa0YzElzNd
zut0HL9Nkoj+0EewB7SjdnBA7tK4RuttV3NW1iqgW85xE2gOx1gS77BmVegBA5R5PgowX4GD4ZO+
Pnv/2dO9m6EmBtvfhOVslFcCHG0P4Cxco+hkJkcul1OQi71XTsiBCTUohePuhdtnoRxwAHf2eUAt
RFOM1sB7iOFd8aqFaIWTNWVekwl0k15MRds7Qik++hXIY+RxLXMguBSKM0ip1qQzXCYVK0CyNsTc
/VG+EAEBFyk/d5do8rUBYakO2FdEb0b+ifQMH6BnVWtPBC2P1sO/B9akTUDZfOEbbs3TpjCbQw5o
SrcOno7UPsNmRPg/O5TR8Yb6cCgRLgh4eBk2VLH7PQtWxnopVSiZ88BaQV4qpRuFxoXW3vWHoY4g
GJBBuvR/lE43bEfHDTXj16x/6OF+YDMXnFSsRa/nxkPGhd80g/XrEveqBcl669hgRVdc7tdBpHKy
XsckmdF40zQrGHz1JKqICgBUhbHAOS0boK/3r5k8WWpekt9/HwdDgTzxxiNSYGGa+dYgVnmqcJ9e
Cye/XIC+JVRHbmJApaekLcF4rdn3jOw+CtoPFRdSEJ+SIcXSJuGK0mThU+cZeds2T5lYm0h8LJT3
e3RpeEDp9oVB1WbacQwxKl0o9pxpBYOE96NWItr6iqWMwgS/cdmpeuGt1Zv/RO4jnHe3rKYqS9AL
zjGLTbAop+anBTyGmchXIzvsNDZSuOIY8LZvj/u/aaFyHSC7ILXPbt4TjAe+sM9bxAq0t845I+zj
iY/zfvnPTMwmDMyR82sAi5IjQLsw+uyYR0kaLjR1jBbspYjr/ez4b8v9yACM5SCOZIp1JSZdAN8Y
/tyq9CQUSy/VFXE884xoQuIt3IanzTRAnm1YA17+YBV9ievDnjBLMZSsqkiBxFeXKXwwlkStTvbc
spBGKrQAspFLwnB68Pgfoaj3ChI+Md9HdWoFkpdjOlQuvRN/ptuQQ85IraY3JypQOlm/xT6rAhsU
gURXLXVElsL7kKBFcztILq38Ss61tTSfgaqi3eHU4HKGXOVARjFMufRguKs72qkEeYFG5BMQ9yzI
kn4S1EjaN+/wfuyExVsXnV3tcZ96hjLir4eTZiUp2fOL5/EQqbRRJLgyLdq85sfR6kfcZrETXGPK
ExbHk7IHLzymACJVoKjOEWvKnJmuccl1xlMNJpZWsELFn2lUoqBaQ+nGOCwt2fT1KulqCVCanMFH
MiI6T1WtThq/bTI20G0BIEV6+l3TI+/JtAycjseLyJIGo06Py9dtXMOOd4ckjNBIC004hF3oQKri
EmsFaJtm4LENZ8lbZcg3ETaMjo9LJDUTUHUVD+j6mWV7mRXXfFMpbm8PR90OBBzbp7r6+vMBU6Xv
jCDfIIJuq7j6rwie2TPGPG8mumxfhcgvAw3Hib5qIvB4YKyYCNrM4zEwcaxKlSGj/y3ryaSlj16N
9Yh1/+0Na+1/U9N4itxXN9zuHkcLAkJFvC79D/MbEP2egYDU6jIv3/rcG5ik8cD6FIS0KnO97WLk
xBM5moCT8llCYKrI9nPi/VTfZOofZa4l9IuuwQ/747znJSl00pkcceq1FJ15Q28nXWSUHRnBTTrw
cImMvmHEskO7smpMeBisO8EXgcBRB+GCiyyrONeKIATnu9IJRFd3xAi9u5N0Vu0thjqdDxrVngjO
cAQ4SvAFV2FSHoQCWUoEQZd7bWuz/WanCiiyARvlAJyvNgigjEUQxom+GJ4qfCYER5joNm/5ko/W
3kqoWJtcmXg0hpYNpaYJbE6dongYJVUnXxTDQuEBneuuBUzdLHytM2umUP2FFLuK0Fkw1FtIzdOa
nt6UKmSsVUoWdFmT0NUViBTWJiPnpQhMOVPuMQsy50hz5hX/NYUtNNbNMxwY1kduS+XyttRODcEF
ZDUZCHS+KCYeYDjYuNzOOxJySg9eOvt+v7E1DyxfU3NoYdH5iVc2vsG6H2q78+6hQYNZrf9Lr9o0
GHzFACs111yTy6T5ezrSUvyq4SPumRryArR5hM3jU/UZ2EUEU0X1JSZiDkmUHnZgIoo32nshAweF
9QaU04WLFouDs5UXlD12SkS4SDkmkbZTd/kx1KGfacK1qUrlVbWJ4AbTyVlaNLr/thI7gvwfYbhV
nAmUA8mdgb5HLL9PDnyvHXWMb2vLInX2HF1iN0p15F+OqNtYI1qj5Es38z96gvng8e6LvbWCOU9S
2JQs0uEY0cl0w2vx1LW3lxe3nd9QTas69NOnRuVqxLCHlfcRWndFSCpOB8hdk/1q4yPlxTqR8yDr
3aQpPV2O4lcr5EyPFprxGdudzpV4YUI0HJ8ta2Ikr3mXPRY9Pv/bKBf5H4YeIJbGUfrATD+ifaMd
V9hKhrbx8OXah87sEnMn0ocsCKZZEhNL5S1N97l7RJMLIZ30ioFKHv0pahIphUU2dwWBu0EnRwp8
KNjhTflYouqVvmb/EdZVqccLnGbeTwkmTGP5Clihwphm93lqxfmi9rpd+w7VBPHXn8RnCmyomsjy
jdTsA1o8T4QUbrqoucrzvW//xdrwZhp3J1n2wLXcGNxY0NigV3a0DlB2Bd3DJ5mw36dtH9CM/fwi
FnKRR7sYHqyzAhZe6iyPHFXOyLs9gyaQ6RACaO6pbQmvbxkfvc5Nz/YyBf6N1Qb2qSWvgH0++TCU
sJmDH1xfqGPf9s7Z8paAPLhB846mXWsYNc7HzJTvvps0Bvk5yFv3DZn+rIOuHEYwklYHZZHKP84P
qwUhdEO5P+OyHx6iyJdFo3AZH6qYjzBIhbwgQDOWr6PC827OqNZFrTDscEjcyAw9uhBfrFs3BoWU
FIW+vttMnwKj7UA/AvnVVd9BnfaRRCPmMs4G23lLGaDO40U9NQ3o4LbzgMAgLNo3kdB8WJ9SokNv
dnxIFIzSvs5Av5jIUzI1l5/Cd4fxhCA5PUHT8zad47WmzdHF5KMb2PeSt3WlDmAWO13Nxc7pL59T
kFMnhV7fs3Ny2MB3pL0EJi8xBXYaA/3uDHMyS8ZoWkSBSDyHIa9cjZnTWcaevwl05ywNvYKkO9dg
P0G83ro+uIA2CbBItMOSgUkgy8tWP43+PAB2OXzu73CLS0SJEabiWEky0QCPZWE+ryAAwSIauhX3
utrXKkSOqP0Xu/Nkqxk9cJlmsFaQ8wUyT3OOrtNKYkuApR8/E0aCz6CmbFtHBjMHvPfWYPVvivrW
n6/unkhtoMbsMhMPeXqnH9stlhzIfh1F7byhP9ceTq/5wEbeP43Db60vJxtXSlaMTQNQsbTaRrkZ
7fGJAMLOpWXpA2+KeD2ui/FQNIUbc2pkpSoMTIYiBY64Ap7m9J2rtymvyvPcA0095Kz8IE0wDSct
RPee7mUBB0R44/X8p2jmnYs1HD+vzE/M0NM4VZg8j2MLW/+a4dfNfSfV+bME58hb++nHFSHminoQ
lRMmMvJX4t9K4PtY62aRXMDSqTxq0JVxfRfadIejzVW0eROs/VYX/p0wJnAbXewNyevqHwfYacgy
DAPnsislhnDRLxHy9icozuVvBV8KhCRuHuBWuHmBb16ajLyReNKt1Z3YKDy3WhXKAcFApSFYY1Ku
VcA+/K+DoFElAv2LpeQm1iMHI0d1L5MuWqNA9VYwoZ0jJvE8SNXbc0OlE6+DCTSg5Z1IsfBhoQDm
ZJEwT4rojjGmRS/xWfsLXO6ihzmDNLIJfoR36Spro4lRX3TdxYsP/bmEs+yV3KUJ2914QnuMGbk+
5OsKCkLxWYR4oAMZ0XvOB2UOfeELJM3LJ4HpdrpdcBiFU0UYGAgla2Vb2lJCYvZ6lxHnlP6cv+w5
tPdR3ycM1mdkbYqpoSSGCpEyVI/qMIKCZxITcODkN4TG2s/5nXdvboTlRkgZOgCdo8cl0YX9EG8J
Y899CFFCa7NPkIbIOZk+OAp49o7NRmxHC8vEwbInkFWu0rlPIw1HN0BvfXFgYJN5YyyPgiho6ACt
J5L49Yl28fFf310B+187lBjBjBdZikYlfcY6sOXwVpH8cZ8V0sCDQAJXPLiCZ/dfKRtMuZtDaVzv
khlXpI9DNaIpjiUtvTaLjYhLtl13sSWCU0AOI99o4QCE6jAPJhDJjZkeKRNhdR6gjONxjYUIUEw4
D2ZYY6DtuSB8SOV5B1Whkf/cTBHCbfAsbo/TGdramgyknYNL0er/Wr82Y2k5bC2h09XBCriQ8klP
63OL3S5GNewJ9EGOudTItG/BW8U6RBGp6VxVLKSFDH43m9Wkrwc4Wt9ArkgpOH8pLu7ZEKclFuq/
bd+/1Uaw09OroQhYsRrmVOH/UEzXSliNuc1A0Mw9K1S9jPgvVcglbIU/AeBLPthdzB5Yta+2Q+6H
Cw5oBeZp9N2uVs358qEF/OMSR4viVyCGk8/jYHcdAKzWxNRYjsgYvPPRJA5APtrw+McwNZESVLSS
sO1+3z8U6Om2TD4CEK4hrvH4I+EhXxvSf/nmviQ+CmpNCwj6EPmh6DFAUeW+Fsfqr7VAhsWOr/N4
XDkxKrr1czXDJRDvGi8reC8cElTN4BseLgJ11SDyrZUvf4e1rospAFzUxbt085vXeBHAumzKqqsn
hpwuK2eJoHyEO2gLx3RllSh2G+DHWQZKf4zUmWgtTomoOl4Zj3AUhqpSx0ZXE3GfIpLVAcT+cReY
jTlcseSzrG/q9Sq3JG450/JGulAjNRNgk2bBqgatwyklY1JOEDzSjWFKe1Dppr++rqS8fWHtuKjJ
+x+0eq1oVwgd7tHyC7tQJyXPx3ryAG2IoVu11cyf4JFcFKw2uSLOoEswyG5l6qF4yuR4BG2SLa53
AmblAz1HEUMO3wvRk72LMuOMhgmxfBnkBxyRURl+cSd8bRPRk2RiERitpX3MpsM2F3RKfGJJ/02T
I6CXbdQBi3cuSbXCaVRU1Y3uyhYLDxoklgflhsmkuvXbwEMPDTrm6Pf9o9pB4OQk+SaNpNzqd2I8
j7WQQ0VG/Z6Y9a7KC5+kj/vt3ZvenEMSl/Zux4foGxtsYEejDbSD5WyGMQ06vAzsaA8rLcdXgnRu
Arkgdo52uYM2klLuAYc5m9Qcmp6jgL+xdNt3dex/Dhk+o+AJXq7Zxq4JsEtzIyIq8ABjb03KeAf+
NR7OY0iRqlcgxIUOC3K8M/7KQtx7XF4DBu9RWUy2oJ4HvheV3YJMp6k5fzSmUIFUTazarb5V0Qdk
BwZR+lxCeawB+UR1QafHMVNWg7N2q3s3FYAZAabuOLzl/SYqzHhmHC+SHV1gFtZjNv7u+oM4TBnq
OjxBzHrGVdpStx8QjooLbieZyJoJN+Gb1hio8fdW47gu7LbuaAKouAaPEtPTUuZSQ0YuRvjshTB9
bSVHmKQ9dpiZj+i/1cmiiELY3ZJaXMeyByF175M2tTbHkCX4YkRits2LOaXKSZV1sQKtg3Hk3wvc
E0c2AxdDx8UPTHSeiV71k7cxNgialN2mZU24hu1i0ChSJXOEpVQaJLqQbZHAQwMRseMktwQRmYTA
TnhJxyVhE4xAY5JFJZUPzV7r5NcKXywbdzJbtoL+3fARMRA+hZrhgctF1TT71HqqetTCKo1CjrTK
kbPR41fLjzKVaDeIBtALBahLHngyt6UCGbnXy9h3g62CIovVMcz3RWUzlIM27+1GqzRITpDb2UO9
01C+MNu56pb9hWkEcM+6PoUMTBl91WbYRTjbvcAsTwobpqaV+riteT1vdNKJ8zLdDK2bemAYoN7x
6G1XlwO5dxsTTAKD4qHtAcceKVcxOrS7AwkrUfH4kckavqwvBqUdf4HYbbjxsBTL+wHou4ufSbgn
Ph833HTPNVz1CyfO3i4DpcJXkbA6S3VV+EBADzla+Z73LCEat8d3AMMJJ7nkJseDEae2RsZ1WaPx
jlJlG3F4JojBECklwcXsIFNpMx133QbFPZ3j+xqsm/0cUnPuJsAhTmmUh3apcGeKJzDPj7qOfwG4
dVtenXy1kXATs88Euv/p14Wa6sM137wbHJCqWNsyNNQUzL7EFnfyswGeXnU8mXJ+Sl64Lnuwmzgn
Rkdy/0d4KwcAkcJ6aWx8I4q2G0oC0MVeR8UEjPiZl0Yf/sWDJiOM7tfwuubfTmdm6qDQZSS2j/+F
b1d+vZ6Eq+/13KLYecePk9hwk5aDosz2Fhxg5Pcs0O2UNuVPaVHi90S7fC1vY5eVCB9P6xKFgLjM
1N70b/OSimOULGyLdC3FVClHQKR+k8D8kmmaudTe/VFM5MprFFy3NIrqYCV5l1ja6w6nFq/D4ZEf
+Nx4jO886WratQ5KCHe1JZc74cxx6USf0Kf6sRgbgy4vedyIEY/MfEGslPqzzruecCDFQFhh7wpm
w+7f+Zm30ghBPh2RwN5dcxnCT9nuNLR7jnZdmEaKdtjS0f8UyVMZBQOx9k9P8eS4CIP/1Z/E5Q9H
amg33sNpOJRek5xQ02g9ZDy3ObHXp0dYtvBGrHJQ5VG2C0xrHnpvkjmVW9aw8z4z8ukTKD+Hdq4O
ijhcsR+lv/wjzoXDtSa5FxJ9v83zfzd7pM6xLhp2HWG03/wtHb2PiW2ygTrbWQ9sLWSFB0THhkz0
RafxRaU6umtmWcgH8V1oxOUui/wyG2UTOEsY4XoGbXMP2eaAOD5/sgbwAbEcqy07wHVvyKtvUhLs
e1Ktk4eSlvGnerbOUpPkcpx6/A8yVZOKHp4xKzcYlAxIbAD6ja3xi1lNF96Ca4L2I9LIY0Q3WB4d
KSlzzG2/OXVP9bPVMeyR77Y3PRkYJzN5FqgfAiCpzd6nnkIghgMUmTUeZjn5bbxcg2Jo0Fi10vvA
ZvpD/yN8Lk2YkyWdiQsGWb6vhMLXEqjW56VCq0shDOorKNg+ntztJch9l7ACUxhdBNA96XRCo5RU
3XosxD6g/elHJsrOt5WEour8nLEfybKqZR50AFl8WWNCaMyf4qJ3V0opqgKlD5iRS/C6pRYG1Lvj
1scPaQUueh/qgi4ts2ch8eM8JBFJ+EUDIB3MJc+Mkj01ackbf6Z0E1UGkWYefNRyAl5R5E1wEv6s
2f55XEG/EKMclJW+d/1Q/nqiUTHysBdM0MmnEhmtUqh8b0H2ZF6eI/ruJKf2T/X7mip5xtv+zN9d
5yitfUNkPhXFOnG4KxOHFOmuwCGnoa2qwN8LaIcGrVLCd+Bqdhe78MUDgEz5QP1h9DqOxIe/RGv+
et6sS62LT3shrfxnjWl1pMldGL7/P6TqxHS4hu3x/D+D2oOqrjV5gAADpwuiJkKE32dsdXoGmYuY
1Mzy49Ukj3xwFVRuVQwq+7Stf+rTzRYKMqXf6lsYstvZ5uIINMW8rF+2597Mf3CqCJ2b8zL2tYUY
lUyBQV9qrGgOEtBkE9pRW1HSZOWPsRHVOuAJ6PYiC+d8TcXDDxpSTDzzNqkcLWjftAGdFiGsjkw8
sna3vK/+NodmJiJU2UMqGJ0cUQRacsb18qlfhQPt3cejBLaZtzjbEtN7PRZq3GiL3q752w9lOu5a
me/XTP6kdkqblcibFxnaOLIhr68FqGwwjp25kTSUfTeAybJsLNL+wV/VHP/BfugDH37auj6t8cgs
wo+HLz7cL1K/AbzAlJ1zAixDZmkgPzvePKN1j5MJr9P6GHSli/CQN+CTR+aNX0dxtmPbVjPJtxAt
neyq6ryavw+oqIObFTY0jxJxrX8E7DPLofmQYKoRnfZ5HXZfsYB8uDw0AhDzSb9O8Rfe2VBZ0tJX
lne2+dBvQJeNofpr4AhjZgCgGuD9Lo6X9TcZ60w5yWJq6g2v5XZBHZjd6ACTEwDs4Y7xtmkKtoGM
q+InLtjwCSXTNCsE9bGWN/D+mUAJq0HWSHLjpsqIJ1H3acDHfMAd8UsdrqO82CwEvTnd8LsoZcS4
Ed2Hel6dWs8rsEiuF11xtqXC9SpNH3lfyE0ZWm53+3VgcizgoF+82L4ys3oBPMVTSaogQy7Axp6L
fTWblSeMvIGvRh6kklx6I4ih716oL+FgTrxBt9+HyAnBdSekjUCj0g6Sy141tVqoVV1Zn8OL52v+
nE/5QS9vHOGubGAC2x52sr5POKP11ZwOsUGBS/TApEgG1E9rT8a+Ws1o4m8Pz5RhM+08kX/6Z8Uj
orCOPOBQ678WQoCVbZ0+kd5VEWjnBwFYmV8Pn6SqHp3p29oA38QjV0bW8vcKK8dwyxsBZl9T/l+C
+9QhDTyGVfxf1onzNtwTRJ++7jTeq4VGq7r5pwvQqiTG5Mpfbu0J9azgu7dQUjWarPS1if2b1W6V
/hW1kgF7pe5YVbVIDFuxd1gHVTczi6e5jD06/Kfk17RYcKfU/xHDDCKVLODjf2yPJmZiS6oW7O/2
ONvdsSIA3FoPj0kkZV8ZsgJTZGm+vE8mw1yUk1ULcrwNEc6an3RY1PHSzgxgYb9eJEKNATgLLJX4
M08W/oyy++PtWBmJBVfC+uMDrch4ics3i7CpYloEik3FsNd2x8sRcSMTEbLbQoIp8QI4/F1uQWqz
N9GVw3mK6h6phm5bYJwmDUrAk7TaaqttoZyi0f1rvCdu9NJ833zOsDXQJSPXBTYVCqBnaXBh1PZy
uFQiBCiptxhUiqaLLl5MVYJzR1omGBNFdYgVAGZk4cWwfT75jvuTVQ9x9J5GiG3dPhsVrpJRrpmS
kg7m9LRJyMpWyrTt8gs94xH7tGtLtwkGOzsLS6sDhoVjlFny57SCTWuFys0kGp/LFitYlYBz6fqC
ymv3+1xaGvSZ7udLeZSF38yAnkLXLdJBvncLLn34apDJYeWEJwUsw268QMPP7m37R6JkU3xBOKsT
ViGr91tQlFsR1wLRA0drvi7XsN7hEz6gtMMhIj6U8FoEF81g+sCJSnIwpLQmoPECjr04+kwj37fs
CIBXxGq807/dMGod/67aqPSomxieR/OuqfucV2JPmDJT+DJrGsuspXldWVxCogCXfB3msgZUE3/b
boHV2+rebLxZfB5nYtGSLferVJoJ316gol52BGs8mcZnzMFSLOV86jpFxzZzCq9C+f+d2wtOAklK
EcidXncC4bwEXqr29GcI7dKeVSI0HWVuQxMBb8QsVRd0KsabhUE+3MWDKEJeQiOGAXBroZqh5Xud
GfsGB/5oAGkjLXs81XaAwYvCTRbMbaTYUsgRJDA49m1JfdY05lNcy1egFYVf8Gav4On6eDTnXyAj
79GB+Le6+SjTdt89RZyo26ydSx1K5J+/DmwhSEPomnJCsYNlyaaLSTLXiFZfGt++PvcYqtmvr5Bm
NPDQgW0TYDF2HVI9sIG464S6ZRRHmIOS3KcjDsb0YRmNqxQHVGGQqnT+ehnJ/OXwAN2Eof0i1wIq
D8A/BBr8YMxjNTXPPRZk0SJw1rbQRwLEEFNudHzJT3t80+9ipMzruZdckWrV80t5ceOHnLvlvuU3
t5T88Px/6d3SFUxdiMpKdJwI50FguKwWjSTWBPfBHZYKyJNpYcX1uaqKNC0bPj8KpvPFlT/7azvk
tGGKZu3hYp0D3JIQeYDsEklg5NEUoCwhMTuCczyhfpG/KY5q2XZ/UvFDaam+OBvzRoSOI34YSNrU
MEPxNZxwX7wEeJJf5eckT1kTRarwlLvwMOsQHUiTGN9OMyJagLglJJrbRs7dVReAc4phLps0pb+I
4UpocyZlENAuRag1ukltsKvVdfL/VOP1j/5lbtRZ+APGRzqOiFLMr4S9a2uMIMalapff2aOpVX4Z
ite9ndaBd7e7Ijss0GweDa/I39UR/t+d8eEOL/EU7nUn7o7mtmgHeR9GJ4jI0NUqP8iLqeDPLE6i
SycCSeCjI5Dllpp86AwPFi7APXrk0AJYzB5WJN+nC+5Ob9PWXbBFXONNhZ26QhO1r1UL2Z+rahB/
FMbzSeSvX76pijh8AnEqIsmwlaM1ztVydV5KAtHwr8I9Uc/BrhjFtSgl+yjuMq6G7POwDAFJqF9S
kKKv74zctAwuGHFXKm5cR8Yik7cVNnvy3vnI89YNCtOvqc19dBxtB8zBsFd3YmQZ6iAvdTMo5DwE
NJHMdzgJvjXrJo+uqhhld4iiH79jg4xL7QQ5WXynk0HRdkSzf2hEJSqCJhPO5HSE1ioY5O/WvYEG
h0BEuQPZefftYac+2d7EV2O8ajZcngx6lINT+i0wLXbUaEqRTcGsnMoNWGvHkQ6bRZunyfB2E8PW
qy2V/Sulp1axqriQnQsKSEzZxgxpx7Zb6UaSTl7yFFn0NrMqM1oURh/x2DbuNpIubhnat9aI/6v3
Gm91etJDFmpv63pG3a6+4TIRijVq1BictLlX6Gcs80SyKiWKVrFHE+3zIkoBkZt04JNoXvyXeF6P
wBNFFgaqnugLWELCpwg8S1Br5I/urRPBcnOABPNY0h3b6r4rXiQdXtYuSe5+rTWrli7yyGO95a4H
IPxIvOKWHMiBjpXh5kKH0hCCepbZB1sRobR9p1wYtnk05b1AaNDUSTJ6+B6MCYlDgGcG1APAinXl
JTkv9Y0RYeNNb+JwDbV8sDZ6DlAsHbYEllapiM+nWlszrXK7s/ePI6KncwTS8BeXgQl/TkO7J1mZ
oYDb6vxlHklUtSLBm3GhVgXUWc+yxPl0ZLO22oStUv5w3d3jyU4P6Wgxdgmhh250zPxt1Yh+qpMh
F0G7CwjqIItrt5ioUAb7V8r7j2zRwkJRoXz4GOnCVyr/j9ab7KlNZNHnhqMpN95TSLXeZHMpHcNd
3fuu/ceBtQfCtZuqLe8NGsncwObo7vsLYmF2ttKtoefKT/P0EemA/t32rwNwbS9wBdNvRhYSW7D1
v4Nz48YTXLRwvQSAsZy9OwR/mc6WbH0IDu+UbcW8CZNZlx7HDRgl15wmS5KuMwGhv2zRBHGde75f
5/oQxc4Mpq1wQU9aKmVbrFHwIP42FEYibs5wi+UoW61hCXlsYPEKnjP20njAUUI4cSMbPKp668sH
LlWhqmPHHtN7ewXrE3GTv4t+IzHnoRPW3izYciazmkrS4bmkovkk7U0KicIZXcHkE/zzElv4koqn
wO3uJ/C3kq+vRmVdp4+XJCdFdUYsMZcCYXAANz3qGK5zZGq5GGsx9+CzRw7/X3KNXN/z7lgoIcoh
uXVxUxQ8KI2pu8ONqa37a7U7DvwJSkX+xs3+fxDa1rSkBZ/HWVEbvsO7zZWc+omNv0eKgLPtZPT1
M1hOwEf/sDW7xeLCKvAURntH+eo5FSAUsXvMHq1rSDCqzFaqOwBZ7sXh+EekLMy0VIa2cN8rBBi8
KZYxkltd/NGpjOsXFWipJ/CTUF4vmuhm5xtWoy2c8pi/JnGvMMm8lRTSQfgZtimRFFAO92amrdmm
BZW3UgaARiWZVBYbKjkpE3+6f1J6laoNE5q4uxPWYcRTrpldsNtUSy/ZERa28JAG1WKtvi7X9t4I
3Ma06TBsZ1T9XnqVsRp1dzUmDHNPVQuEzfESurGTr3YHCTHl6PTBP47/3mIIP95ApJF+KEKGlsbD
afcItjGp8LwCYF3lvYgWOvmk7z1G6tLej4FfmbDRGwIrqcYmkFCELSb0ubRJ1JYsXDiYV8FfnQRS
L32i0g8jjjTPkJCjyYJWIRaj6eB+SncmqAHPHGYRXH0UvOAi89P11tSYX3UeZPJadmaQtuJ8HCMJ
UvyqR/fgdCw9+u9FCOVaHenEIKkqFmdy5jPz50hHOwztWlRLo/AfypVrsbxvhZVENIRyqdW7wLxI
BIisiTsXNhTXo9ER0Ihhh+cnZUZUn4WB6c1PzM8s14EjDL66px5oF3tu2pzxlBh6T/a28sKng/+u
1zfl8qqySYTB2k+EylICGvkRQDRGZGx6JuTHcBWL5ibB9OCAODNANz3gZdL3fcZKk7XR9iVONS7P
jbl0+fIHW44ne8GRCRSQMR2nnqwf9S0Zl2UeUgsLK/CGxyQaN7YH51ctNjIyvmvknXX6XKXPeLMV
LZI/LcLzXrlJOCX3lUVI3Kzn4WZBcAZ4E2FU3AZ1nWbKzcVeReiW9WSzRcr0dX7PRqYFzANy6uXA
zpD1W4JJ0eOryCd5d1/nstCEoUEi4NF8NSclGoiW+K4vaLUWz6tbCz9D186uCMxIeW4P9JUEeJVb
DM6vnYCOz+g9I+xPb1u/xzzbqmVumcwKeQhHLfBXiF3K2r9bahdOL8V9/hJxLWInCfKXHKsT3zit
0OHW7qfluIGdvSwtFuZoKQbuFK6lhiBrBxTHA97Yl4SXvcbZcKyTSmP4i3W+JRRf42QQ6VNpAikm
YPax9UOrGpfAJAsnEhjco6vicxNcknBZTFzI5sg9I963nx4WtorL9ohL/PeRj3iOxUoM/k9Yex7f
gxqCpS0r43/tU20KLT0zgx8voLSma3lKj3XsO5d07iNcAiaedo9Yj4x5xX/WIC3AC34L9z1P3f+3
h52hHTDg9WBIKTVhSTBtFJq6DljUSSSQXpmafbx2ZAXleNMd9j1Fd6/7P0cHCuFXcu9zn4GIw+9C
paeZ14Kv7IF0IxJ8aRmOww4/i4ubVY5Njj8Uxh9Udto4blRUzvHQR9CXjVLveA5Jt0KLmG5wE4WB
ycYeuyAufKZmJoKvSbKRUNzNzD6Ry5+910zLsHgzXl7/cJsOwLGTNmbUR0G2VmX92hvIA4YpRooB
qBkb6yCx3dXlGgXHBmrlI3tXI8Lzg8rSFgNE4usTOIpmtgzYUX/ArQd3n5kuYgaqiWeSuA7o6njA
+XKMCEcBRyIbZ4BbmKVyd8tw4GKQhTzXnmcQ0Iu/q59ETONFS5spbj4odB6KI6abiqB5Vga/ZMNo
pkzMY18P6ThG6N94JpmvzHtkxW7GchCpZcpQzJcQBRezoTF05lKwySSu9tSzJItkAq6VFrK2fyfd
JPfxjg7VF/Ov3MFwjFTlDAugQ+InXd+Zz0zM/lI18UjUshR8vDddhu+6SR3vS2V1TsFV4RRUsB9R
lOFk/cNOH7qByNmdaWZQa3EHWD0UoxfK/tmUuFPM16NUxe0N/2q/RE/X0TlB7QslIFB40dnmX2wJ
J1DIbMoODJ6FHr9NRKYsA/oYTVbBoWgQ7CKC+vNXIDEyTFFKNUyFmONvYhkdsxH8/bYEcOEbClQ6
V40AVnZs0tW/GaTYyCxqJ+htFirtIAYY7R1KFdMGt26jyCA0l7PtBDo0rBwCCG/zABDGDjrvAWoc
9NUmlLMu7xqmWPRHTZ/6Chil2uGzJUcTSJsL1etmrvr8d7ux6UqHMeYaDrhaLOGoLN5EQAgyVlWg
XANRQgYYFlRDqK6mWW91dCyEPho2MbeMkLg6cdCYbZv+l8RrZwg97uhuMAL9IOpFmIoDzlleKzME
4LCoPFwAliZE8c932NoSlntezYKMtQGx6HT194wSM/EhabU4fSCzPuATyCuloAnvTHWd3LT6iMwV
cCh7Vh4RA2nauSSQcY4CGnbM28dSO5rkH31FW93doXd5AEWqdDni+umacamy45BCWNl3jqWV1XOY
dZBizFezwM3/kXgu3KWA7HKw1IL9x0MHUFQOJaVIVc91Dqq4XxYPs5A8G6LsdDZ0C4Ne3RD2yyUO
DzpYXzolhF5jYSXVUI1WQUn39HZgkgDwGAbwrTFl1WEhWvm2Wr9Z+mMGpMm/SJA7dLIkQ3KCLy9D
k5iSnTyCmJ6DJkF6rgWQ13YIvT4zDJljbs/iFaskDlt9mVJnf4Xw9VoTlOt1+S5cTNB7XHzJF9A+
6bCoTPgmv76tIvuOzn5Fahdd+P640wlLSqwG5n7qJ8tLsfMFCZLcZRd7yLrSQt9RgKk+bYsdSdY3
dCXhw9YAJuIHVlFC8n2n/66Qv7mgyVSWeKcJjdrehBf8uHuCeX+5EkEOwpSgtz3vKP+8OJmAfflW
765VN7F7jOlp3CvPvYEhRmT7bQPvA6lbbwVf6hcIJsvrrvMAVzO/Pt9pcI1fd2NdMX5pioMpoCwY
TdaefpNJL7BvGZYx+U4LD1qaPMYKfBnKty4OuOT0L20IZdH+uPe3V7MSHiYipFWtFwZX3YgfRGqI
OtVmIjG2tvuhQWOQqY6n5aaDuXOTDZVs7EZhDLc4Egolk0wmU4WC13E3xANy/z8UpGay8MvSZCGx
DMil+aQ0gVUwaR066t0+uT5z6CF8jMcNBjnyIPYdwmT0O56WCbQxhv5BjFifJELI3pcCp5+i3zrx
f6oOhUop2cMjGGSLR4Ve7WKSmbxcpcq0vlO8rHWSvctT8iS2/D7O21BcQCR01h39uW3W/7hLLOsj
LfWCBy11L9ot+llgVKvHlcSoVtKFRyuwEN2dHSeeocqheaMGgaDmw5PYL+rKI4hMhg0JbWpBbxO6
+uU7gWtn8QE5z49/TiE1tTHPE7eYAvTmOf7L7KxNf+w2vJPBoXTCdxdBPMLgN+/ZIZyS4G1OQotc
sSmYA8gF2NB7a7w7Kl5RTkzl3+pcFCWv2X8q7LehW5BkBbsbQnnZxMaeTkqSZpfTREsT3+8pmQGh
3ZS+eTffxtQjl5z8KaWw+iC+erLgy4MMg4aDj8asF3XIRRHs98QFpRW5v6QTfcjGh+gSqU6pIIrA
SDCm3Bht9PlO5aM3FsUJ/W9LNnaOY+5TSiQBJHbzAz8uUxqtXfKPG3i/SPab5QgyH2OuiD0sfKtt
v+1FJpBDfaRuArsH10MjbqjZx6GsVsHXLBveERC+hNkPi1EFcwyI2bpH18xeI3x9dsxEPn1u5vD+
l1gP77qkGVYC6crCCrSGqldSJfT/1Lt6NtHGpzd5/WjhGNZBdWPUVEVeU8wIWlnIHoqnCE62CRJJ
ZFLDBIX6C9tPPZPIrBOqqgphfox5G9ITy6oL/RQwFZM2bJcPyxgGkD+bi3yjIGpDSb1c4NxjwM0u
LrFXvtDC7SokI71I4aEnCjCao0GCfyR9MEu1ZAjsqW7ypzMim3Vm1rdPaGrI5xBpMLuDa04cTaOT
DDSL0lyJrXl9B7bjoHbebFmQL7xwvjd0Lndi+9woMXEbUzF5SkRWw4EC9qGBJaEBl44qVTALzKiv
MWndaAf3XTFbHoNsM5mPRcd2TaX5hlZa23s4Bgblt90crepl1IFmnjyfxVPY1os1op487kdELJin
XezJ/3NA3pOwKq+UguHEOztBpo+6xgDPj8eAzdhNvfhfJPU7GkDv9hBTdhPeGOhOKindnD0aRRF+
JwP3LRJXwMk53XAqBHLaXpRQTcz7heJUS5XrdpbTe4P3Wxk5ACLfcsj0QSR95J33T3ZreRErl8zO
nOozH0+VTAfEDCDZ22Y2Kc01+SF6UrkIn7+9IXQcLgz/xON9+zBiq2PcQx4IHH3amZxYwuz0qFBZ
aPKeMEnZHGgobaoaa7aOP497MQPMhrcIEe1DmEErGS9wGeuStFAKOSCaGZvbTnkJWL7WQr93wA5q
BWCkAVJIFWXXLkQKBfKyKAOJPEldXyxrikqKxs1kqrbyGYXoiLyzCsUMUfLswMjS+QBYOJkVkH2S
gwvkMhZiQctAfU/mIaoDjS6zRpm6fal9VEmF/Wty3RzLUQT3rlfncrtg7m35gmLgMEl1ibvspFwB
xg5gJymb8+7222bVTaNyvFI8V6m2rdgwN2YU9cnp+GuMYsBsRAw7JWxSoq//qYxF2vdbNUdif2at
LpEYeLe/0CEfNMR8kYXE1YZG7UV7SUswNS40beLHs85PrA+S50XObs9iEUWdieLPERfbmm3Hbi6C
Z9ywUyCWJfmRqVIzHvDLZiwjjFBA944TKsyNsf+WCS0gysc6FfWg4eeWcHJ+mGZkIRKo1bpOvle+
IcAeVv0TAdUIbKO3jYz8MBRmwlxkxY6eU0dW+N0/1PNJLEvI9ZLLUtoGmn8RZl6MiQPf5DpGrUJV
a34xAYIaVON6r7EAwTcSJfVQ8cTG748iBbdG8Rp2YYMlmAdou+VxswBI6Il5ZSLnXANqoOVIYgC9
ernS9O4CxPlp7FdxbTEAGrgApA9KTCAosTJxcG+96UiOTJ1cYL4FdMENwF8IisqAGzlVoII1O9uW
pVWMDl4nXcRPQ1Jw/9V3ja85+tP+/H2yrHhTMHaK3XqtxLK6v9nIMz0FhU/Cq7+8TZwsidDCuJvz
tyuQtgMJoUw/u725ONqDK7vUHDx/9F2JbiYYbuoXbIJc2DWLkpUTqBFmTEJ6da8LigXVNBjPU4s/
QSz/7BEDCtPz7jQfuINIlEIVcDkDz7kyBpvMmQ612p+6gp7NqBNK4F/WZvQ/FCmv6XFPNZQl8j5K
6NxAPEmPXSZI/Wvse/R4nDv/p3i2vkBjl7Li5wZ3A32iCczNJx/Q9tHzluHgfohMiK/wrqJHUBVy
1hW5X4kKVGBHstEo+0j/NLX3hSoQwOcoxyBLvcqonZC0xfho2SbluhoVx+PkSjwx0xdLkoghzAC7
wjv/3faD41Gr5yA289KkOeJoX7R2zLt+5iZqAZ7kfrGU4aM+RXu0vXzIWfLycv14bRyYvh8xZ4f/
ohV5A24RC1Vwbcgp97geFBQBX9NgG44Xn6Mz5Kouku8TxKkjBPw2e4GtSF0FxKQ4G8Hn1P2Ttjds
54sTwc74zeG20rM94ArfvMX9k4cE44HTsE/ryv8Ze/SaUa8IdMpg5eH2Caw4CjKRm0WbdsRnFeA3
pTGpmXARhlKpp2b5nqbkatPWU7UaYWJYBq9sTOHCrIeHILNYWu4JgSKnjtQyepglfbAR/2y1vw9d
kylYtqnHIPtS2QmntjU+bduQbuU6p6Kyybbqj6WM2c5B9dkjdFFb+eU0HpnFiI6TkzL2MGyfx528
KYAdMnUA9JhE7Lxndd0WhdbZTgQACaMzDMBMQI2XgQzHeoWcUKHUxT0TqJnp09TbRy7B1g3Jz6p1
LEsy5SK/ZijSSQdFIjXIcLoXIHU2NYj32MQ9MRQBvBWTSsxhs5obJvY4JZezBoWbpHxjZdHctCFO
Ux1XLYyGFK7akmCRW1KOmCCB8jVt+TMPvnMBW+k0RKFaUOxxI9UrQI1Ctgwnvg6pZ+PheuOBUf9o
KEYbli9BfIe1Dk9kptV63yp3UYbEOACK5Mptl6dIgjGKjJX4QfE4bUoSa75uBqTSMbLDdEeWFOkk
h7pTV2FlnmNsYwQybFdAM8yWiyPa8elia4l/XGzRxZ3Xw3D6isblDi96hY5SuHsCLKcVPJrF+T2W
nwVKmhlG96+dB//i8yMiVIAphcA3mVlgbjQjEK17+5ywyo7qYSqunwrU37qCFddfBj4+IXPhjwu8
nZFCwWddiODRuoRn3P6SmL8K+npn+mX0C5r4iu/+CvvfGmTpknsdnPxMRP14smYT7PvxlH3v4Dme
BJsExb4XaxLhyepGYNsqIet3nMMFbxETMomA84Xo9Yay31ebFJWBeb9ZopDpae87aH4gjyiRGPdD
RlR6o101KEjpWk14+Gi9mzHb2MzAAV/oQoJkp92UWG1A84eN8ajxa/W8GbPME0GwQa2ppwXk2W91
xu8EqzXosxYaFDi2ztus4qTZDGoDnd9p+LLGJ/Um3l35Z3ZCpK0FKhmXOsg/f80RRxxPcNBKERpv
yU4pXAm+0pw4SkfDsH8UdLgAZzqjQWDCM0zralbbJegmr4o/Qsr2OkwdXlT/mq6rHZVxiXCGztgD
WeWBMV5ZFU5qJFIs4bCIVVZCmjAM6WoH/1CFL5ymnjisZ/GdpgIHyxewg5PPdpNvlJfQDo5GFDKo
jztYMumKHxqxeatO4mqjJWttkKLQli6XrVwXPP/nxtV+1qnWwuhNXSasWgKZfIbgq+ncwinWpLYj
QIA7f/Fi/lDLUcFOEVG17AS3NlH008nq6jKgOgoDAdkkO6efEl36qr2/K6UwpZI3BtnuS9YbHWaH
w7xy3bwPnGoKzV+gojs2LktFPhDKVDju1eFYFZahstPv+B2miRvYtaSA2p49a44G4k4ZrBD6wiGu
iiyVf9SQ3cA7Uvs3PhsG2LSF9jPWEvKq1z5Oxf2ncs3ajUiX3RNOuxBVDDwCzaULG7ZVqAMCke0G
pTm5agKTjn++OUX2F1cmXyAOvamkXpq/Fk7mOjrlA5/h0syhkjobqf0hjBkT3LJdt78yCHpny/Yf
dNR9ZV3rletTcqfmKTW+nOGxhovOxfAHmKUhQQq2D7oK4WEyeG/EN/2JPkUYgefNmzb9OKmaTV3H
esmi6TzqHNHTqfU8RJAt2vZYBVJqPXVpBWiB7wG7rTKasQkf/DPNg3UHnDlDbN9qTg2u+Tt7eMpb
SlTZujkLB9yAvpwOnOTz/APCct9c9JUEQIX1yp+q3w6Ug7mxvykknmedhwiwjr1PvyfjPlEaee1H
kBTvz/MnUg/eU1d2PRUwGKBuK/hVNybtlcgnTMKwpP9tRnkov5KcYk9r2ArEuoBpu4idzsAK4jck
IqkYbCvTNaAW/GcBAwwLvAC4vA/3Us8WcqT51TEjiC2ncVkAJzZGqBMmhH38XRiaAkC2cmifOpGr
HYUuaWQj/ckmbuRiqXVUrMo/QS41IlVThNkON9YyHKHYQC9fOl/3aohk3rzaoWlxtpxrS8gc1SWF
kvEw40iPy83/4FDdKq/hDCOzkQCo8oDCCoYi6f06MW1lCcgOVDnxZL4MquKLbI9tsAeKw7FN7yT9
dtZilsMX3JvRBYU6AiHSEP4H0zD3ysxsUb6YIc36X/KtgOeK1rYhyTWVf7vHvlnR5V34KZFedmED
g8byPwQTeesB3wL5tXieoMmgZO5FkNGl+vbyr6QiJR6azepUyRW53XBk88fMXdWDq8/SKnXhpJEv
ZAqH/RNdZy60X3hGqaxAREqy+QOgoiLM0C8bif6Jdc7a8E6hR05bIn0rA2DvhvuWaWB01Bs/Pt+U
/l2Z+7Tw3BEfWoLDa6D9Z5dpA0qIUZn2NqE287l4H1CD3uzh+gVKPKuQz01QBse7dbhTz4rphnah
nkWCd/XAsJlj76eo8BSjCn1lX+g1S6MJLYsR7/t3NvbgkzXtjQF47kYXqbGsJkUI2vBpKxqEhmP/
K5IfEbHNLTUM0+EbRNmAoo0/ofu1AAdLhyGQGL190eWya0hC19G+2RarNWHDWMwh9DpIdTnfRA+c
I2HewQ/QdG+O6eFe1eQLuHIaQuDsplwc8K1Aw8LA7aqcpsArRczgo9D2PXY1WMKuopuvskkfEYHP
8cM+FE+/ridYYqwDYeydmuUgb8tInaTnqMGyn/DfJc1nSX9H3R7Oyj1ClNNY/B8CXvlpdpwuj86l
tmLClrb+gPlDg8mqj878OYUN3RGvh0R55O/XLMUrthdr9D6yO6Tf571bCDvaR+pdragd5RqvzZ9e
mrmZQ9QZGaxMwLUwuwrWDFrMk/j9w494lWy3829IxL7TE2yxO+//PMFho/e9xa7EQWSPVaw/ULBk
moON1wpxyUmRFqM6pC7hFfo3a60b8KfTwOm//oxThVEm51DkBEOCxJ6cqiS2vQRydP3mr4a7VjEr
QpAQgT6zGSZbHdNDA1pVEqRYCUCTo2NhnWG265Q30KEdoswGn7mGcaABZmpgDAdHCsoGbKR6t22U
1Av5YeZpbEy7D921YJZpTPbhVmHsXMtemI1ok9Mycgwm2B9EVY1NDpS/kub8lgAZaZxWSSMsy36r
+ADbdS3K+YaaXkFWai3jITy7IQW7sMDi5hewW8sHsmlSu1XNvhY0Q6M4mUcOzfweao1lJGb23vr0
yknIccVOeXQE+UsaVl8cQ/T6w4z4z3zCzxwMUBhx9knCrkGj2OGMj55NoQXae6ycYxpMJDQG2t9u
LQX+WHCVm63feICnhggUyYJvbqBC779vTlOcTpXzPchb88OaDV156nGZrjjo65iLSpal2r71fIE2
ZEWzgBmkUv9P1Hr0XJXorJKOz2LQuKEPcRPY0VsA5O1ENU9KObRfhOmApBIJgChi6H1GZejgQTTS
IGegSEWv3Yw8C6Dc+GWwVncfUR0I9Hy/vzW2Y+jNDDFJRqoasBAagoIQ7Tx5tnMe82L64kFIuE8t
LhlaVog4KgFjNyQHXnBt8wlhnVjlC6mgJB2vle3lzMB/pn3sW3ak4gjb+H0o1+25eEw+JDVs2wzG
dI/hik7V8Koe7fQoi1wBI3viiWDdW6WKa9dC1QcT+hQ5E+0abna1ychX77e/hUdKvrcMGIRIxAo4
SaOG4vx4GlKHKV5/1QeUyo2laP0L/hUf6PNJ/IQNURTaUcDZmG6fpHXiX4zGSiqFwMC9ihq6wgdk
iGaRNtCQ04KZ7I41WuI1hESwdhWJp14i7CFxHD94hakf+1prT1R5gZRrJgjrFenKUOrPOiDTvGsF
vnHhMrqICg9Ldt+3/Imv/IinXvs1xBvfBoWOK25xlc/YQLa1+vQHPKLgwgrVqGUXBmPD8H76FEaT
Zt0KA8A9n8wkGYtgL3weaJWYGAPL1bB252dtsfJomV7jhqJVe81AwTzZomUaUBE5QNvnpWlxELm/
IxNZiF2HZxF9GWn414YKlkjTqqm9RfN3bWxsI6Vx2qTmhyHNXOIqs+x4i/uBOL4gAVllzu2YZPHi
B+k927armdzloqpv/0Xf3n9ZQbcClnNyoNv4Li/g+lKz8GWsUkPljF2PTWtvZ0QfRvj5UUGPCdMw
KOappOExM7+zGuz53piU04ge8BUAcEiU0zTIZQLYBSZ8L2bsKG6bb/gIo5mW63Cv3iyBxJGGt2oy
/ZOty3oeNwd+B7by2xmFUcc6vOZUKTyp66T5AHClB3P57N+ZpGXlwvku5Qnaar3PBkkDBuWHJIQ/
UQz4VzJdV7CXhMCOjlGFN47z5VnMcKzvkASv5Y5iVyQDvHtC9wL2ijVtiilyCJo9I1Hztj0bo9lF
uFfXAoobyPGJa4o2t2DToBBe54R3fs+7FtqAw4KEy2jk9lcZG8xDqZou5mXsANQiXvZEM7rK+Be0
y0DkLYTfEVe6MUHfthOhVfWPXXOie4BDcA622lLGK6iR4TelztDwG0uIkWqZLxAnXsQzRB9MGHCI
YJx0AdBdvgmmFOvk0PtOujLK8pJ3hxQR5U3g5XLlRxwNTiqJgKoFuemSWcb0jnBNgQXyYqF1Doyq
/CTleAAwsMprkShgVML5xJS5qdvMTzPBes7sCNnBjA+1y0nbcBthw4BbXfW3YVp8SCBUl5CZjYg+
X+rcOe2Cnf+0wod2SqvJZVLu8B30hfq4d5hLjEO72Y2FQD+zYsR5wSEqqHWpZhxJIt9eawpXNoif
OvPzb+vEy7QCjlDGcww5xfuzjN/H/5+5M1O6jH3CiLkWJS5F13bEcrDr4Gd+JCv8LA4aRhAoXr8R
IIgXquUu2Q5XuacMnh+KHen9zhOjCsKjytQB5A/CbNLSmJgaEYTeI7WNXHHlkNPI+moH8fpmVkQ/
oZovgRbzdvXCKPj2lwh7RC8nVUF80wDTJo2WsVdx92IcilmBvB3uQ0fuMWg8lZQqZFuKUWfKWma7
yxf3hRVLSmssTQMTuv/I0+pdPsl/+bda54R4VmmFkDqO+7elbzgeH6jkXR48ABMs8lsck7Is9dgj
xvuUstSHUHxtk6pUC0dq1ZVgHaass+l0xKzonEOVTCxOr1bayO778LTj7WszFKrgj265OL4B+iDy
LWHkkD6G5UUghWyMX0pEwGuNHbyBn4H6E2thiuE1jHYypUjUwjv5ZUEXBWiup6pz5vlYLMh+1/DS
4YIbKUyMmnfmYQUtMOox5Qpgb6vXhIdbTFhK+8RHf4CILGkWVWpRAlm3yE17w6iEv3C2WdVKr+LT
w6Dj8IZk+ElWrO93bEVjAHdBXHruiwLWYCJrHQEpZecC5MGPu4y0d+44rwc86rCOQQc7QBqh19cy
/7HLXsM30/Vd0Cc29ZzEUZYNB45xktRl3eNaWfzTwpMwGidmKvLH4DmxZws20tfy3gSIHIs+05/F
i6LNRH1JhsS1kYdD9aGDqNrWpKsgJ5NfendpRSiz0kA1XxLQceq43el2IrlwjEIJv3c/cJlGPEku
r8vqy13MYVNuuUkUal/hZlgHKddZ9y8nh+K6va/epJpW9C1AOv3vZHHSteZN8g0DUbjPGhNyI7Rr
nX4h9AxfiY/n1O11Ohi1EUN4PC1AJCNqkP3ObRhb6+R3+NCrk5MKDFndXmI9csIc6ZQU7OJ3XQcU
GQ5R27z4iH33pNbAF2R38Nthv20ElRUUGyTAUpo1VTI8t0zrOvg29yKKgAc83+PYTKRM8m/7bbms
14RjqTOePUdUUWpVI6cd4E7fX88OuU+E46mNmh8TOCbeGLnSiU+0YfxEWY+gBCqAGOVe10IQPFys
sU/QAxucza0FAPT4c4gBmCIzIkaCrjhvsuvr1XlEoTv1X3gnAQWBlgZLJjCjt0kE6DLTqSNwegAr
Qu99wnsBAfsb0arH7T+Nn8pU8wVfQtpAPitC9+97wHrVkJgkdornFID37v0ypdtWL11pJcPFHQIH
RYmTJqFlbaAb54OigAOU/6Ky/Z38MvBYgUk9QKBLThvSleNwtG4Iksi1x6D/i16O8cVhLVL12MyW
YR3nw36mLHxn1U0C7NeDn+OvgWUKlTumP94pDVRvDisvX1nJ5Cz4gMMxfVZkyUxFxski2IQn8i7J
6MuhRfPOXQCJthBnogFqlwOXNlX4N45tMSGiNjdlwxlA0eFqZcNJaaRwBc39HTs77g2LQ21H28nH
BgOLs94zbWemEXGqGD2BrNG5YKIDBjiCkrQY7Y3b6zWkS2qHx2Q3dfjiDY8RUeW0vNyF2IsZhAAb
5N2PCP50gmZBUAzPmLpSWBVfh2sTwHy8lkQqxpJ/HofqOT3oUlINL7cjNNtmJCBwa42l2aW8uZ4r
U28nbHtpHgGWESq6XiZhXa0NU4cD6Ny6dfj/ZrTMmkSo4CGb+KUN7bKEWINSmnOyKWP251OchkVH
nnU2V7Ww6ISCPBqgZ0DeuwJ4V+EIEswt+V9ioZC+rELNOYIagdhpViFJWc6SFaeh5BOfoD0TlkoV
j+2LStaK7VXsdfTMHnMzd0274YarMzyTSz3jGsemF7hBbK0Go+MQaSfG16vxiXCPtCR/nLX1O4DY
9DHCH7LAxOlFJPANsIzPvNbprwmwAg+mW/+ihUnNwAelLSrZsTJsjnskKsIps3TM8ei69bMrAiW1
sZgdBqWu/hfbwUGdFj+ehsByBT6pRtgUSCD4kpdQmIV21tKAWM7SIP6H40NVoLVtsoJDbmp5JxG3
IAjK1bEbqDUe2m9F3PdHzg822hQEwvusj84CHuoMy7PWYSu/dpw5Go5mcE1r/qo/qv9FGQpgVe5T
6DmRccPYhBIfUWQnEgmoysLzN4G925tW83L/gNQbN4IFvlGKdJYKU2bg5XV8FSUrUk9JRS/P9g14
fC05Q/5jSdH5Gcs04pkJ3o6e6NXYxeehxHdIodGh3Z0qS303Op4WKlqd/tQOt+wNqXF+WtpwoDAr
5zM785zhI5dbuPAZgE8bm1IKi4314BqZ9M5hqvWTKOLtG0/R2+3hOkGWAsJpzwEAdw5nBg5/lvt4
Yo7znh0b97HWlxnU5PmhLrYSndR6HrayZOBtrYKIlsNmL23Vj72ayWpsc2Bok6eVbMvmv6AQP8uA
cwaZJS5xGtZsbvS5zc5E9GuX1erwJ1H7QvfWJCFn+VPYQI8XdmhxiZdA97Mbdqsa+MqstwuUp5PY
SYEBOMCiyXIIlAfha168vRBC5iTdjciyQla1kSp8+oKJYcjKEf4fCkb/Yf+xoBq5cHwcK16lakOH
ODAeH+8AXsr+dU9YcO11C9bCQZittvF9zCoTHvWZsrDIRIBBdq48Fme1MXFiUcQmvJk3SDRmqJFQ
n6fSWEtyt+aIgPIM9pgc9Af7SUygynQikTFLTcXUSVhwYv2dLRItOhIgZFyVPGqz9M8mHlJXe0tw
YMNTnxRhAkqoYCifr3GndyjpYC7gH0jw0zSgSsmlqkYZGJatXyH53as9gYQkJaQ7ssI8IIXUTwv3
3zS/HkAXvPStMNXY3UrD26U1fpLErLDZzy/6FNeZHBVojaREfda/FPP3TS2x8maApiL9CjeWlal9
Up7bWnQhA/jQ8VQ2ed1hNpiA9Sn3tnP4ur6VwHFTHU4x+yYnOb7+MfW8atuPYz1BDogCNJXNtKi4
eAAgUNvAgA71AcMBm88BW4ZUBEQ3YhedmQY0hEjngqeyhADmdf3EybvPooCjEcE4zWTh0QDjQnaX
u+KRA5Ufu5xjBh43hf6vGvoij77LtiD5Z74HhsTDtM5BeK5L2K+X/a4PfMdlyxfRRYdHp0JkXEe7
Xt79/3u6TDWaXaCKc1WC9SNgr1k87NBeLsUPrpzdgQE3T1tPYa0smNqSSy1XjKpiEUz9+hB01oOD
tfI+QIJuBn5ehMm+iyNrpNP+9PvqzWDfEtm/F+Pn0z+k58FJTYEnJjJ7i9egmsSoQUrys9/26nkl
LkYFaT7qEDKc+fjkAkSY2OIbYGFV+b6AL1M8CWgoOpX2o6bFYkEBwtUuj3TBz1OhLg4lTdgt5/Ns
lxG1stHdZTMGZcbLsyVJg52crlhGG8Y7ajTJ3wrhzIC9wYeypa/9GVaCSUlTOW9a3JpjvkB6+D0L
VGaNSMk+Me3S7ssv5KakNWlFBmr50nXnheIwcz1SGAx/zR3IWRTdmL2VyKGNCBetcaC2/UjiUPe2
kSIXKi2evZhjoJya5Oyl5rd1Tjm70SMUQQ5bNT91dBOTQjtoR5//nr1MbIKt6lvewVSwKFvwHq9Y
ct/8CxFk+lbtoppdDr2smXF/wd/jcNTRCRXtRdnQif/vPcI/lgPP3sK+gASTqm/lc92xGuhfHK2m
cSlwGkk7/hMWBmgEgKiX3+sQjxAVuDVPeYQypQVTC6iQK2Mx83AZMIIQHh50VjxxoCCXn0HkBR0H
K7pW863vAEYUPFZXvezMQiFa8Cx9zIBwKbPqqfwdD2YStE8g4uraUEkvWecbIy4sLIRUn9WjMFqC
wBppfV0sqpkU1r82C/5MREnjvDQ6PGn++unGRRhQK8NXdOLJx0bWxK2yS5kxevztN3yYGCuiL8ri
/pJ8iTTHaRZZNz8AM1+OyjPTsVcbHmF66my43xEfrf2mpF87JtFHv2utqS/tKR5NlDkbGFi6Zy6j
Y+KeMEK2UvRYIF2wT9tVyVni9+lzM+B8qQxhq9+VReKqw98uHzAj6xJnRM46BBQDlXqf++YKZmzi
i2GR1r/pweFgCK9FiHU6n97m5yS5gl8ak4NtQsoJv3qPHBcQK4mPHEFMn2GoSmxcno+FTSALHyhE
ywZwwjgPIof8ppdTZAbL9zQoWLXalO/Xh2EE9Bsogh7H3IYFLmEVQohvDejmv+pobjXQ5HojGPIj
ufhWl20m3MwBL2CFZaG46MOyqz9v1S/V1p/FyaFRmdQSiNJodVea3KgQyway4CBT5RSTY8Vqzu8w
yihoYkllk7lN+zP7uscTcioR3onq46fkJv2J5ydOCoOY7wnQB0i4uhqbPmYdfskdyxQZof/Wdp8m
SrkpBGMO7uTJjiNb5FwpZJUJba3/r7S4d4Ywmd4m07bPQboyXubtdbEGz7HBx4BmevRF3/4EZ2lm
IIe3L44T6p+QvegluwhL4M8PwXyDcQZ5AVPdAIvkSb9HtKrvIJPeByk+321nAjvdT1RlEx1iMAFC
KCcvuSLMA/3C8gX0bsPZKkTMHHR4Ewyi2BaEytb0kxpidVSXJxlZ6LANr3T6+LIRcgUMNFVPeUhs
vp6ZACuMNReW/i+m0ppkEWRepcbYnxWeuf+joNSjp4UhymuymZX05ASvHb6E8nYPwvKKUgy5iH+x
2tMZq1yYDG+c+6neyVF8qe9hiOBNZVVGZ/Bcv2ZI/0nW9MnT068Cex4LO1Pd7sOyRd2ko3vXwPIx
j4ksoRpEwA8C6v3+wLvKIMPjyg/qwX/0LSrBNkISQSeOyrUQlxI7vT6IG5etmNtrEZnR1wNMDgym
0FG9tM7pvsgqAgfXAp+gQhRix641ugnEraOqs8mD0fFQKNc4fycBi7j0sbmLrVe7blphT8M1wSet
nG5DSzkiXQplAwCT4vHgu4XuOkxCA+nOXBA4D9HGq1Zju7D7BjqyDhWvXaraUnBHVUilPfB5jDmS
nAH+56GYpICQJ6xywUD8GCNLfes35ndAL5OMP1eKbLHi+zWPCEuTwxYvre3XOQ5SGL+TMtCy2m69
TdJj4hmJPRMfc3s16rAOgojP0PIsp41hy3VeFkSvfU3xa2eYKiCSk2O1UEmLOsUL/6eTDF+FFlAu
NakHFqWQYKsWIk7CYv8AvbF8IxnUyT6uW8B+ZZ/AsNic/akAVU1F4aK0QFpDZzJcQ2fTn0xN74OW
yr/j8DDRxQp4UklDTddfgzy8ipr45S7LMmPSikxlHyS6MRguzWc4rvEJVqX+13N/aktti5+r72Yz
OHuEurtsVm7nIPkrCJSKTDfmIbbwG3wyQVdGZfD8d/yVbjCtyrh5afhLqTCUz+vxG5/pHxlUV4Bs
uBrTnUyw2qrHv40U2x2XsrMnIUwyDJQQP2Lgf5UavhjL+giBVlYAueqIieBjbTMgrFOeHvLR4iFD
WMZPTDSls22k3EmgGeXJ6F8F7IpWtkOlzKiZ/6xlvBV1IfXGRSlrk7ubq757p8/mpyiI+7bg/WHa
WiMmndS8ZbyB1SPkFWdL6O9OrAqURHnXT8zFvf53TBnaOA43U3faBCO672QN2Tfi3umGApXXxMHp
e3nDQQm+PjdOSiYpJ+wD4C9lUuj3u2nCFMSC3Bwz1YLdkKtpIB3VkGrMOTDNThPgQpQrkpX/Qdzr
byNrESuACNs8nmKzlYgA7mGMzLMHxh0VFbZj9ng0C4CNtHEJ/XE11DjkbEfFkFU3cQ+S8VO4ehYR
SWdL2X4Z4ukzl+85VQmNk7sq2Ojck//BYI/hVKTFA9w3aPjfZ0TLtgx5if61gnWlUZKlvObV2YwJ
MpJ8q93gMeM+/RIdSg+k0IXtVOrq3q2YKXFXXciFrGJ8LkxuSDQ4geX/w5r7JgsVhJUVHEOq55e8
oBdD0nEa/nxxlVlQxVQZSSGxoEl37/tWXSFcCjSGSYldzD6ooo2JgyRvNJ+UdcIMf7X0wyEm33yU
DN96Z5dlnmq2fay2FNulQ1OIDcY1vcb1w1f1dixpTMHdaJjVRVIsOSE4CJpYcRlSNc1uaevDGcsb
L8I9FREH/xUctaXgX1tDk9AjSb3XVcjLP261L4yq6u3Zy6iLcxz66kaDaJAnVN+ugoVCr63Gko/a
mqlV/dI1GDULs8ccDh86hvfUsoTgG//02y6MAl9h8tPoYLw6M37wun+geP07sMV2esLaNVUJ4p9h
WbNtFPOR55mA2aRPQsLoT107IG+YlgL6noWDdjVBz/nZAh6fLt4iWlLoNtq1JDorJnrnc5/ZB7gB
CdbgktjAaRoRtb2Fugq32C/7Vz41Z0q6yHRytBjxlsdyfekOLVj6eWcD99ZQsQKHcmmoVURYir2O
ou+PUrNHxBsLg7+JxAKLqTf0vpxx0wMhbVU0KQGI8yxHJ/vtRcqFRrv/ijv2EN8ncToVWnnzGCH4
ud8wYY/EeCXO++SMicti6H2+4VbCgTGrzkOqfdlcxz/iPN7Tth7FBCAdPxC2U3HhMc3x4HwDyVTF
ZEjcX/5rFls/dQPyyMkVjQns29aQUrkJY8PSICVtrDacOqoAog5n4EfJr9lJaIIbiYYA4lnISNIx
QGX61x5YjqZs+uBi/nHx/ywe6e7k5Z6FKxIe7I7EJc98LXYBE93tf2mU1ol1rkpe2k8+i9NUFW0D
HCdYdHd+1p/1D/sAXWmT0T/Iepm6THGipumAljA3iMTk9N4wyukFFnkF2qDirE4aWZQZqaFeE8om
m09e4tERDje90ryGqFpl/KrKzbo97gYblmnfTQVU3Ay4U9wVbU20na3nBg8a3pFJiag8jj0CcO3/
Vv3m4IA0yPb6Q5o0AEADKpW+JGJtpWulIMMRI6NP3dwERSnrigEwneWLksU/pHeQuTmVnTtlIbdQ
ywhY6HRNagDWHjhFSzvJ+8AvyviGic3BM7VP7PsddT8BILbvUj3FCavih7MjRtG2+X2wBTE7qnmH
SXpOG2FkMi2BJceZjR9q2IOYwzpgxJiopqGAVy+SIc+WWagT3PSK59UVllGUiG8LlgurPsjeKsoN
sy9IS2pVGwtmrh27Q37QUggISESgc+3B/8sKELf/fBCHMplNCl1131IhI/i/tAFUQhakapVLa3EJ
YhYInewQxe91JesAkZUH+UgJdhgvEE/Hu+iWTUPv5p2Ye624YUJRXtV9/Juq/n9tRrvAubYcETHF
RBTPAueGdlziD9V9rs9wMcq3mSid24fOStidn7hD4WVqMDe+tbYRHTH/9iDq/53peLsbQ7EkTi+V
WJUGL6JoIb0jSHxSld2VMhpsA+Y2L5Eus+Fhjk/+YRjrumW6essqzaJjzhf7/TN2UNMoeeYcPNsC
1GILX++ysKxrgUcBmxV3gnwFX7hJPjXd0hE3zS1ZchsaswXLbn4iYYicpCiaw1YtMAnyTo8NorVB
p6ZQG2qN2Bn+n3uL/BcC3B/aIC47/6ZMs2TS10tWPFbQk+fAWhYTWMgu4BKRFIyRrmC9gZGRYfQi
2XrdKtpDBI61e3H+7HSiDezShtxmvoy+4PLCRcIaKqAS5qtIbadcVi86hN5JSxZc3OB6ki+8SGyS
6S5YOMDzUCZ0LbwGp/24Ldb1kzNkHCSe5Q2sRlhOEgborngrNYOoLZOqxQ/5wKFy8TJJa/Pgs/TU
+f9I0BQVtbs8QmppBV7jq/ZJ8KCDnccW2LyeIquNvxfHTmLzpfyv/tO+gVhnFBBP6KZdjHtbO5sy
cQtn1xDtEhNWVSp9fHwb1Aec2fs/69GXRO87xadGXcyuxHi8Gnw7DDmcxx8ojpeXUI9Fa2DASVXK
pKxZ29bRSqdxzX8Fx1e5wAeCYqo31IjG7oOjerm49YWnhQRYUaFzjwjuzRfhG+E7/U9E8iBMoMKa
pSm8qDXmm3fjAf0XuEiK6J0pTnA7SU9uZkxAkqCfyHG7PPlvMlzP5PSn+BhamE5HMmB7OdXCt03p
AO3IVEMBWKUEATFHWaYcsAvLZfO69bNfih287qZya17miqRWa4aukuraLtbgZjIQMmYHt2r8aFUW
VXG7aawa7+K6JAb/RcTHVYQD6D7QSdF/8VEhDHpRg5/I6m1AOQgcBqDPSURmWdHwexM9MsPgtyir
K8bfLbY5lQQNzF7ZrnRCGRiDUo/0j/tMxT2bEZ5DHBLUuKqvVdVuNbb6NsghoN2616Xnz9h35c71
aKK26ixEKjHnkhvlPKmFH/TnqwWShBTRxrH/3Uq6N0TMpok+nezu56tUCN079r+mssbyBTnkuwmg
sfVkIUbfDzYIlPNRsy/Ikr96IPO0M1ySpBU9MNxEVbyhFOXeHAGk16+A28gfZdyXSMyjuawJtQ7+
Tp8PkfNyJB2919GHjD/kdZmraZQx4Gq1vmaZ4/Mssff22JTwsAB3ms2jK2HSFutJm0w7Mrb0Fbiz
Ox/rKCTfj0kZfm96eSvAyaSwyO+8yq3vz8VwT0g4HYlm3iTGHodpfssoQHK0bYgAFQCAny3nk6sP
9o2Y3JE0Utiy6FUzA/UZTBuN/uT+ecgjOvSONjMAyprNCRx4HTX+MhtIBsXXk/TWlKPfRvWjkily
CujcmormHAQijwJqNgV3BjSm/ugBJVnDycv9k4eQiWCrzSKQ4bc6xd6sNcxrQncRuXsDZCybp6Ac
ZkbLr1KaYeoE8M4rsYdqOW2Ux8X4y9UFGefN5EoJDoImqufwnxbQ1iTbHKxIoMz9Yqsrj3Ynze1b
PM0s54dzIHHKpC4nQ5Mxo9/ZkV7fFms16sKIJX+FlUzFdjMYiA2DLyIMDjw1E+S9v0RjbS3VOEPe
Oi5zS3EMSq267DE72yBOoe4drVbZj+n+SqKSTgUa8fcB77nfYy3UAWhZt7+bx9/2PH/HWA4msYoH
lM8zVtVo5gjYES17xwyH6mRebb8O6rBEU8dgnrWb0KWocgOuqc4qSdhHoQMiqC+Fm6O+JauqmNu5
3QPei7xwG9vqFc39M86Eqs6UrJncdC0yhgmcMIZTWLBd7v4MShCS4AZHed7IzblwT4Sy38J0csUU
w1TTnVPZkMShU6MZIlP2SkeQRnrtb2+/eux8Jm01EWEyCVyE7erMejkQ93gcTGQgLgeIo3Ay+US+
83i9ph0JLdNjDt6Epv/mBRbXlhODzGxNAoT6AJ4HLxlnaZVgHkEryuQmIH5KhaIrZV6sPXrQqt4k
mX3KD2ToXY6jHOWjpOh9yb6P8JWfPmvWqk/+0BOYDrIJ6f6bEVY0CEfh5svg2t2fwtQh3U2mLV03
vol5evgOWCGfP+ZPCXboBec/DJx61C8ILpCPsr/UJHtHi3yQ8VucoBJ2u3Ckee+clt09JK3tGMAq
LNjULQOboFNxXhJaQKAy5yZYcww7qOXS46zL03/jfK9AYe75FAbJA5p3O10IuDpfUv4kG5KtdLYj
nCX1CnY0HHeKdkkIbcwsOgPCm9Zcu3eFrE7X8TPnp0kXDvCKrhEwoBl5BbAL8XW/5pl1cnje8M/M
qbbGp1rLTUAYMnoKMAccfEnHPTWlNrcULQaLaPCLABx4Fn0IaIXIu/NO3Ql+emcstAxt4WSKIxuf
1ZbhtDPQufZOrmxP9bdvGnhY+ioKsAS17DD/BZxR9RkfxksDA4lkJ/No4Z6eTZSYZe3bprF7y8rk
9/lbIpW2cyUjvA6rLS/PzZaiOtnUyTiRrRcInvAqfveDpSHbL0h78PFG2Czju2E0yJwmWCjsUQJH
lg4yMRSwAbF62PZ7ckBPoX9rmaexSIGWJaSBsfWMlXwJe9Cq7ZHfDPnI8Cz0AMMg5KH6nj+BXqky
bBPan/OcfBoZU0sg7n12LNygzw6tAVaTzp6YtyjKvq4Nzevr4R10VIY9lfwEwzpXNzTxIrlEu5jP
FTMdDoUCguiNIy4xt0vkFkHwr/88NbkFs0HY0STbBd2O5/wt+BoktX3finL7ZWfsHINvM9HeoHCY
90T/OjrlqYu90L+QP5RGbWkfzb+ON/VUM9iXDx78b7R0FF1RJzCgv9cgGDROCXkW6H/8y+84ITty
bpPx3ZCJ8a7kWwQxXM1IXGF4Xj7koc19lVYhf1aVmwKKTAALWht7wgRbIGYJmpxQxv4avqi14s/m
TI9k1jMSywigruTl1SU1+nvvPqhkHWznMG3g9oNIc99gbHbeaLhWc+nyyEnFK45o4A4+61AAqEyE
gM8xkt8w/lKX2ikyFh007mfeKqzAKPjJe5vHXxbI1cL+tNrt4cgaWR5QPQMlDx4NsEniL418ylge
VxtxXWA5MQm+eZoAfNMbjk4EsbPmD1GnCVy3Ie3DUvIVSXQ/s9aLAERJZ0S9dLIPTCm2afBYIKow
73F0nyqL9ucSErDQPq0cyAdYeQZ8e7IhW48Be9KK/40SLZIkDhb0ViETswf6ZWoIBhcmhODG3bH1
yX7tojCw7/GdtZ7mz0Hk3JNpYnZVi3MJgwBIWuRhHXPDndTbesRqGyu9cGnULHn72sfFMDTNR5k4
7pze/B1tzzTFLW9u+Xrubs4C32S9dhIeNleKh6PgEQ5kRUnpeEn3spnIr2w2f5ipY5iIvUPQIoGE
BJwL1krAv4BfjRA789ciX3GGxPNsZIVVPZcw5rzwi9S3cdu1bie6aU+cDQ8Mj4qgbJHOp67YF1cq
N7xOUyszwf1RYrohio/Q1pP1fDpgv87DW5hN8jjOs2ZgXKzU5KD9h5ALF07hcjjomRncla6w67s2
WEzsaZO4FCPkWSRIkLuX/NX8kMyV3H6RHelxFqWrLVv6WPjdb+hPDQDhmk6TVok912opdAxDiUTY
DpAjQm1Yw2e78Enyto8aS5jOjRN4a5jbie8fCSet7VCcVfj9/QnB9mFhuCnpr8obaSbPDtqE6t8+
/vMSK9CAFoEeoSZyBTvCrxkIifPpzSSwhfInGv7dTAsrpSgr+GRBUAFmjKoNEntSLU7T0thqzYHw
th+e5uX15T0nK1KIJH3/TExpOl2yyR9RD0MRwCuRDf60BCjaxc1i2ZXR+uL6bZTEdZGpq5XXfFso
/KmjAlZGsY6FelmXRD/LAmlFDcoj3ClrkjbXJ1oY44Vp7soXegZd5jSzzsE1Vv8Olw/21KpWWSS9
CWXMfm2Y26oLy2CBjYC5iBKbOCs8qB/eHDzsuj7koaOduZd4aB3XUbDwgGB04vyFslTLoaVVEqkR
v0EXjIILy7eFWj/nliL8CAV5gP+b5uKSRO6qoXb2MhoxbsPnfaOAwUZRT9QxQgArk8/UlrjVQaRp
OmhUpqHMBilFDtyfukcNgO2fxblhntHATTNpqxUjJfSDpeRgxC6AkNTsXg15TAyfYtYXww5qN2wF
xrRjVgk8hQEuorZWy5NPfo9wPlSX/n09Nqm0yE9bdvuY4G3dvQiRWR1GLU20X2u/+N33kxNckESx
2g3iiCHdOuh5rHvhE8ODo2oHvtdZSWm4rKrgCuOayhxzglU4RN446v9QK8mLnZ4L05viLQPPgVwc
lweQmYF37yXRsfe5InBFKdpsWaaWoP2y1qqfJUyR8Xcv6xnwBBysCCE5ipkQB2dbfHg88TJEQr/n
H/Eu7cZPg3HMrHh99mD9wu+gVTH9wGi/YxNJoRlWIUHRdmzchNoChJPSQSvAsP02QAfKYAbiMUbs
5UHLkPBGCuIHG9/6a9r9+N6iw+ET85HdkIEYqDzOLk+/1fSR2NNS5c3WhI2FL0HBOdjq+GQWFCr5
dfeSS2vEKtnNWuth0IGFtD24OTgNurI7n5XPUi6RH8owk+xWR5e1vOodRV7Eg9jN1QKs9yjS/XsE
Wbh1/OSQ6zD3sEoOVgpzgK0QHqpoDDDOo+2/kSxpCTj1ppUPDQ3ll69saO409FkH3YM7Cq0fIYyD
NlTRRo3EqqrOOOWT2iSdYD/T6F3ZEAf+8/+c6EEo4tM06XeHz/lVRjzoWQt+i/nF+OZQ27SqLNp6
PeGGnXPulydzDuV5QpB+O2qGmKTevfconBFypuETBkXjFyNDPYhmA7WQLg8WxFi7YZdCjcqzSzVF
h7W42KpiFH24rEoT/CKJ+LgZzIxYAUgUBbeB6F/I3cTVTWXbqhjJ42hoRVT3+4MunRLyYhg4m0Up
SaNH7No4BIKfGQFCeuFstjANMMqyAQ4kXNFP4L5tizeEaVP6+SC/BofK2POwSHthzJ1O2miKoBv/
dM/B6qMmav7oT94lHyGCT9mMTJ8PjbfnHSECPJJ2V3RPMjeX8BAaeDw9rgCqI51cgzJ9BfOMkQOj
IRpRSz+sCmQtwj05HAsEWvw0KTxKDGWfdn8Gxm1L/ZMkbT+BdCvhEThSL6h7NFjpTnWhiOLWmgET
ACsGAEMXysCu4E+JCoRPahHUQzfG/32+1al+l718CoCsPoYPmfSeMKeCMbgxSUfutfuHbBoDpqka
JOgkKwXUZ3YomNc6dkkDbVcfZ/6O4m1LQj9cAa/beBNVmWajdYFjE2ucxwEVBHCmkfrIFJcSuxs+
jvMNcUu9TbWKCZeFjC7XpGu3tj7wBEFZS2Fz/p3vP1V6YPjytWpJd/vdHHLnwjH9h3yPzCwOPoev
0Ak3V+o7g4H0RtsZH/jZq+BHWrSk7l9ga21TMbnvCmgJhrrNYG4B7KM2rS36iX+OKGomucEzK8kp
+HlcxpuKdORt/7yYMuPZ82iiXloEqA0MOZFdeh4ONH9muTk8m2l7W7kjWzc66ELthmdBTW8HU66u
YYgZAZmoBDZWfIfw6xnqu2GpGS0evLe13swn98OACtWWpwA26p9abnd4qUz1ZH/DSobvRVXa+INr
Jo5kn22fW0+De8SZ+K6tjDRZqFuy93FlE/BtBSFQNHGmI4iG0U7yBhoT1oRBptW1Q31ahZWslgt+
N34CG4gqAQxp3EK1IrNpHHT0szv0FF/S8zqFGf8g/vi99UjnKohPCaZEHzXA0EPMB26YhXk4PK/Q
ZZTh+RZJB+fQXVDHHpub/NqR4yRrdP2UpdcD9hM58icWCSJdlrze4HVcvwvOZXn3nYL9Ug8yhZHh
ClbJyHZFJDf62lsqKoiIs4Z4q1YKBkkSdBgvTHg7Ja1X9tbUg519Y8HNrqDnrbkrghgl+IteX6xX
o+CjtyalJqqdpYHLcPEeC2IaxbzKfY+hkE7QlAgHN/gm7QcuktN+/2+uSXS3AsaeJcVNyMZKJkE6
rrf9rSf9QtaOjden5x88J1bBXF3ZLkak2ktpC5i9w1xOkmOB8uI1GcCn0CMXqg5lyj/fPbnl2cz/
dkWh5+uxIWeyNslti876cSucLo3+AvpYzqwWb89KG7qgHZPfEV++F+Nz3vT85R5jmxxBF4tps3OT
CQ9f9se16eSGQNllqoLZMXAJTjGq5sBE6oXOmwZ+oNYvhWgW2b1p3NUrNMYanX8uvya3WBC/YzRz
+/Nz/eANstESLe18uOOBtmxZoGpMwM823jZbYukKzDpxBF47DgxF4tc6zj/O7M2JWdWuPxznMgvJ
4jN7VS3nXXZlEqUas9OXA4kOta4Aoqpdy1YS8aPyWiu9JTsr6E6VuWni7V7yPnzO/dU+vxlLYN2e
mGAXn4I/xSSy1sClnH6m8z4TJLl+PJWy4qzsq2lF5UAIAwV+ENfZ/G2lvchqVQAiWvvnpEEkwdZr
RCDfex/Bu4DDbxEDepIawrEjsYCbMRMi+6NDqCJsuoH8Ojh8krgC/+7A+MBEhQnZY6xi5FiXeMFW
e8zKtlqIS30xLsGqGN7N5F2GcHNZFGVbkAI48vcbvfZbTvjQZ62HmhVkcrcu7NgFlNEsc6VNQE43
dsqMXQt+5K1taEkfjQiHi3uZnQ5U8PzWocEyDGwfQ+Sjzzo+sLJZrJh7aikDpAZKhaB5Xn8iEXwS
rzk/Nnv3DI03mbOOEtFaI2/kHz84MuYcwqsTR7T9lYvk5DlZ3B0iyA+n+ydhUDBFJLrZVENJ8bum
wYfjz0yfBYRUBh+9OTUTG9CGlV0ghIw92V9zG7QREQCBvNm+VHlnTIotJofAvNI7bcnm/N8TSipn
+GW/hlSP/2YzTkGMFqeJBpFFpRbKPlZ1/VhTxbEzTCiFYdunQ6XKuM+Bf1Jzq5lvIujcGCbORlJC
lJrqtguM0WR5VugDMGfjwjgDybOts4+SPWUgQZ4NRoENVWpQmtDONNUNBP6zVogm/2QQTkabR5Rl
7uQVfzHurcWihTWdc6szKcgxI0kR9CQS07TwUQIJhup3Om3hnZtfBJ3u8MAgFvX5/6rqE8wEUd2h
DQhqf8jqiueBhcB2pmVIQlGT8FT1uBCv6flRdzGiIur++4t0veVfNG8zkJS9K+V1nnGtWIpd3vJl
I80hEK0t1QrSaqMYybX/xYe777J7Qa6ybU1zo+mosX/sWUCj6E72YJu20EA1m0mepxJEw7xSnSfn
A6K+dCrIhJloMhQfqvI2jDm+BXkKxixlYMZqyw760OUMfjLefeUCICO360GpJZZ7SaeMGFYchoNC
A9IP4+CwHl/QFopTFHK/LAHwFyYNac8OZgqAvCRU92j4q20uH7TFRVlDMRUvdGIrA99LaM2Qy7ZH
mTUuP7msM+NKIA89u92SWegudDY+NiuP66sMYR62MDUbiZT6qrkoyweotd9mmiqvDN3DLvAQTSEv
3JPwz2iJ+bu+bNyyszbx1vj46FnuL76SR0xt8w+e8dmUiQGT/CDa1Wtx6TNkyepwD4iY9pdXWwzk
CRVhbUehCpDnke7HMSLK82/KFtMsP2sLsouWoYzLl0cwHqabqS3LnjG+BXrKVwGI+4AXgvqwj4cP
byZaUy0zWiqdV3+h3HO25vVphFKuaszzR3y6zzxvLJt0xAa7lw/849p23DMrcYnCT6EnMxrwKfKi
Jxg83ILU4LoDRV5cd+OMHkY3RBkQ9+dYdzGNIV3FvuewDCIpItYg72G6umaof5ECyDHqrtByS89D
pq22QEfc24DvH8Ii+XEBzxnRUaDv6kBh1qlGm44+plGOUZ3t18raoaF5XkWg8FscZLu3RoXP3YLd
3W2ycA29TKhhVfqCLQZHkeA4d0gTdO68vfeXuuRZ+7q9hfH/p5MfmsdUTezkwDmP9DT42sWno9g/
iKz7N2kUdMwBBzKsp7z3Diz7nLfG2BuSpPfDqNqDQQ1HV/TIwPCNkrksBMCT9AotuneQbxcMbmFp
9FERifqB9CdiRSnDStEHyP9yCIs/UKv0UgXYqrqXTEnAd7lD9hxsaEcMhXkaslQQqCQnAnVjMiCI
ob3x9RqU4uaVEfgBbaKdima6OTN/Jopw7aUMeVKkUhWHhJfQEnLdINtcSJQfVolsu9+/5i8Cv0Jj
3K+FASjTqvW9Tgmu2qeFe5l0dA2eMitNWEF6XRE6n9DfyxveLGJxkPwy1nBGvgVoWyPMGYHBx52Z
2ml2ZybZd53FmBBTjF7BglwL4delBe/TIjbdfkPfrEfHPksidyz12koHi+4Ci5UWNxWl4UT5zypD
tLIqDu57l4TZL1aUEikZgxLGJ/p8FOL3X3Yv6JRBdCxkI8l22xMCAYAFiOHx4Hu73HdzJ3hrjZJU
/5/HRziDC4X/c0bfgnI1WX+YEhAC/5dVhg+bSVyAzqjk8B/Jt+YLdsoh+lzFEJWeKtydRzldIVUC
650WYEfTHpY7LbuW2OUrSMjaNm+AyFVhHixqeoUeZmeU1c6ngM1j3Cr4OOgoVeVETm2DZX2yGFe0
MtEnKvHZ3gcMmYrwQj1yX5HO6IdsZWdls7XVFLF9MjbazVx45tcuozKQ0ovHYhxg1ezEx+x+Q6lR
ohqKPVlyBn3JMLjtvKs8USr6ugu5ZnFtIEayFEZ37O1ar8+tym4isyyeXDJaiXcXeJ7ESrlypkI2
iN2eA5YKhUNdT97Cv4T8g0fDAXoXU9B5RhoVA1jeuWRsDVfgyRFQFpkkngqhzlQDmnfRQSvevUrZ
ZzMy7Qbgpm3n0cn8OlG7LfnGoNwmZSdsiYrkmOz2lRpm1hz7nI9Lgo4eEMPDFi99zZnB5mDS36/Q
O+WOq1cF2qJDMVO6HwqonK9IPcyMThq/y1x5iZMda2pYIeDdgZ12Ry8pCLbgSnMsSaNEQBgGhvHv
Hlv9lU+FeXdaH+kJ2b1Jee5tRclkfPK/WjE8xmGQtG6nhd7bC3HriK+rAN+WqSV5GEx/malhaMdy
3szLe80LM329EiKJ/qoUek+BVs0eD6rvRqjCBho5X1xmPb4PSoTLMZXPHuQqhANSL2Ly3beKDZBf
kah1wWUsYjgvWBd4VOCZ5kjcCm8QnH+eBDPPJt0DnP94AhiIUgxtSadM2pktMgDxUzC+yko/sGu1
A+IuJwvk5EV3FEmUlcPaEPChHtyZp8wVXjsIAyUTQoKuy3sldlDjMb7dQCLlexIfnT47FlrinMHF
bRlVQOZ2C7sndQNmPnLI0wuJsuC3X0nGXPJUvQ75ehzutlDHekF/wbmoBzNzQUplWdtBGniCQvTD
wX4p9u8ayc2lVImVRV//2MIAmbUOvOwWee0ED0wxhe9tVbAg6Q8xJNIufgzNX6XklD6ddn3L2CKW
zZwRYTBzp4gBASNdgkjgCCXBk0xf/iHMHK+JpfvBDSLOWgmRc9BdfQEy3WYGfvnmmDfLlMoMIxDt
2JvHZ0WivqyjUjzqgSjc35eijyzHYgiAFxBc08VREhUhRUZH9QnLq7QFIb5qCLEDghgNy4JfpPZD
eVz2jQlQ6f+0GRZcZZJPEKLHv3WiYCEyPm1/ntzlA72tL1eoPZ1IeXO666EJ0H7+ScyadJ1y6W30
03qEPXvUYsj7K0Wml98Nw56YzVip3SUNkpVOH/vLNhmoDzf6k8YNlALFSZtM8Nr+DHFzoohytv5B
QdMkVNUkaLeSbbUcTaNrvd/zuwSxVbJr242JlTWLmk4zo4SDQOffFzrX8ZpwWDl18vIAku3nBp0+
uzQvsAlJkRoPhQpikHDexJp/lDjyQXh41ESqQGTM8nB2PdRmKmJR4R4I8qOHRIdxa7rRdlop0ejc
gBX6s3x6RHsYISg+ZAX8i0yPsaqr0e0+gLB0y0z72Akx1oITW5p161xUlNT6gYllRE/hbX7763OA
V4mdHm3ssl/SfN9/o42UXsq2ZFnrxtPxzA3UadwuIBX0GRJYSHBuxQKei5iUswiGM+ClTgz7FqRN
fANVhYYsWN4+FVSTJKZoDF8nuDLKO9smBb6VCHHrdLm/AIIlXudAgJWJxFSkUuWK/tWk6O/PgZNI
tbCr2ZLdyscbc3+1SNjpy6syYU+eFAyPmhz2v26PUOb8HobFG4zeLBjJPcEa7iVYFK6uZpg5Fl8F
slHMomkx8mEs4Q9Bckl9Km4l5EKrLjsZSR+tYZHAgJbC47TCTvj2N5BSn3OemSJmZMQMmGLRU93A
RSzsJ34gGDM/tmOKIM6h17hmSX4cg9mfCm3n3rL/PpQX0mUxXERGC3MHUlwE6tSDxXHJO9kxiR3M
gYBVn3SdfzsJV6L3lcE+pHkI/qKPfLKSu6r0pDam6Qk8bMyz7RfsRBibfOx6o24B+TkxQYnlE5HQ
PQ+w8OZ+UMiZ2zxPBkeLASZ2oLBluF6zhyI4NPvKEOZHsweWhssqn/sDqOHye2zJW9dBcGk8hTZ8
oj7Bv1CjqsHcPue4wwHSWr0Gk9AYvx7RKSWix35UB9ZcVZWhKLBm3UqanwCQHBaOC91g72sQJoVg
O7EFA1aIUGUoHkRCRBXx64RitKl7oy6PvpPNPnOWCUVqd6ONTtau1CYClndgDdgDgNC37O93+SoX
SdxDrNJm3eFbkuVccdFDeqwTtkTJse3VvyWUAPNDapaJZ53MH03DTqB+io1eOx5VFd9g+7gQNbuN
DH0HdkKpA3jthXRS9I91VHn4lwicvWhtNF3lk7ez58lVDNh93mK7ce0dA9stjyTFrBC3tKcjkTFJ
vDH6mVmXuiVvQaY1vwAxARCoxLMiktaSfdq78NZE0HYCwd8bcu/paSlOwqp72pB+I3mHU2+TEkR4
+0QgxvGhMqtsQySnBn0MhWyHxPZx3QLDw6K6OgX7mW1Xt7iRah7PiQeoPOKH+Tem6tboVz3d1X4r
gADq1KryjEbfVbFSHBKBQsEC8iF2zLePRWyjH/7PAdzkRhrIv95M1i2ETVl9Sq46RwsrQWGcJXzt
Gaf45Z+XD0jjEbF6ltc2X0gIh/jeymA8os6KUSsOU/v6jSIy3qI9pXNNDRv1AIKxQMkkqzOTPggn
Mp/93iZ2s/7Pjtd+PCLeWBkGAK+EAZex+PXkvH5eH3mZdh2P03SHDW5lJvHDy8qS08pMrI4hkJ9H
DbukcGh9cK+oE+c/W4bPSn63O2rOoiyxBW6JZGXHoi9L9BfGbUtBsodVX9iOGFWCz1l1IxxHz3lw
8Di0w3RaviAMqmHcVi3KZUY6B6GIrZSG2pPOMKmKhNXSyYbZL5B42vcSMM4gXSsR3/P7DALs0sb4
YZpiuRrUcI/YjKQSj/UnNOZHYMwvU8ZGRlwNoaqFaUv79caZzm5oemtoSWwJAZQpZmdcBOCULW2a
D7/FDrNBIAljMVo0nqbvtmn+D6qGaMUJY4QnADFOcqGpMAtF/1SJKcRUcMg4uJpScPLv+GReDX2d
6LSe8nccorBYdhwBliHRgw2EYY5EvLxwFPFb0jWacvl6TMOEkud7woGFyIKvkulNSpSgyKZTa3vH
6K/eqcx/0y4z/Fr+xEx6scs/XJHamrGeLcvQTjbaEooSn/q05TIwWqjiF376Uw0NMwCZi0HRVZIF
8UcdW3fUGZMEPgl+QeS3Ozg1AuQBdPPsp4SZwEomGtrGcJpB0uXyFwjvELtHoj4Cz+Zesn0uTP34
hzuCbtv0kKYSSOGekx2fzpkKDg/PSZ3R+C+QsP7uKoaDF5V7cDi8VEtK7mYqQK+nQ1gbfBSGxJb/
UMp+UsLJHg/kn1sg394Y8sOdUko/flq5Sc9KT2MoDLZIcQPl/HuY4TTUhuBWMQhcUp0JBTuABweN
grukkDUTuMRHMeMNfd+WPKiNdL1rt75SXzTOS2Dn06hiQ2M9FW4umpN3LuutBlCBdtfkdmrFThiV
m2ibS7DD30SvaHbJcZ1ayyHrfiHSdf7YiqM5AN37W78gUsH7gEo98+XmpZ4CYGUnz5gty3ty7KAd
srWOdTfwL3vcdai+uRibrEXF7XgYt+0RS3VLyupXF+ORPC0OPlGt5Fd9qeYAlRNwLQ7ronAPRtyy
JP4OWcb+M30ubpKpoER5J9V2IrdZTveJbe45oQMGrORmr6EtjBpgDgBgzuJjYuOYEYUvBE/JmkNi
8iH6j3dffYZTVB/8HP0yfLPxM95TlIPIuHZ8pFmumCCDh9tU6F1NTlyId5QiAJdE5wk6M7slXtu4
gO3zhssA4ZFBzORM07xSexmMRq7+rBnZBP14qreujo5wBZzce6UqisaR2xFkkaOADT6E+OxN9B1f
6kpHho3HgoR1+Jxa0/1tmTEFbNyoI4M3eq0VDLBU/hFjPAxWkEEIm2w4tNkMTMzyWYoyAQFlwAsm
ODxWPAr0M4wCZpdteMgA/dnOMirwRyoP8ZN4twRvKz/iKPNyCnYZqvXB6xt7ixXcZ+tP2MDe7Hf8
Gg7H3J6tYYN+Itb4JF8osA3TXQvQDt85MI0oLm1VaNg3yuwtVqr9okTCRvKI4LwsqdJkgVzbM4am
X4LsZ80lE1HfEmM2fl0EZ2Pwh0AwsrmnDAgFsscXf/R8iUo6/yX+DNW0wmQsX0HzL8gGpH8I8uj+
O+rufTSBIe1b47Cl9r8Rgs5eugov073Q/hYoIB5sxIQRs/Kzvr5kBlKncv8mjwBEgUFgSaHzJPXr
yoyhRcjh+G/oS4YnfAlsx3U7hyCc1OjaYLUjmg2sSMik5NY+CUQ6YdZErxDS9BiQ5YN4zAOKU2qc
2v/5B4dSX3Wq9ZgIpYxW5u0yojX6iK+N+royF9xX9lYoy4xzCCZXnWgZgZLGGFQ4g7ACMxa0Esyb
q66+jwFqRCM8+QMJTgS137OfBgXGir3I2qpvG88pOx25FoYtiac7vYAXAjZRMarwFliJTq7L2rIG
UrPLlgHaHLFIIcHxUhqmbfmEV48DBKN7eklwImiGt1zy6b0cBJqhiGILNu5eaZwdnuGAizKgJ4SE
peG/vwFScvmLsUA2sbvz1Z2fy0l6OZ8Uqy7H8HARctLYH/gy7hks0riAfe7Zk6AUGgBX2utnCZq/
wxiH7a+HtZ6ULdCP9CCQE2cGD2p9G/z2KPtdsr1+CCiYLpK/a4t3UDSabkHKakmhyR4/rM7EpGGw
nQrK1tu68R/24Hj7N9hup6mrbDlT7ofc96Rq/CnfhUhQWxgeSCx88hSLQ/ja46WjEdJ/t0a+qSVx
sBlB+DEhPAoW+lhiCzZtOilfXvjOUgurrmpJ1zvqKW++jCx7LNUkXitUG2C5mGJ60336sy5+Xpp0
ZSJ7lav6ScPywCQ2hKzQtKZtgucmtT+oX0xjg+o1KHKgeelI8gAiLariaUgYqFPeBvC/EQ0xND25
f5q+tFPvmNNQnfHGVDNxTqPEt0BpUSUJk6f8LAnLev46EAd7df0VlOe4SneRblbygbOwfozz0Jee
sZdIZ/MCCQnCgkDa6tZiDWngL+MXunBph748YFNvg4JVixEa0LFWdfhtcnxaNNcT3VtFkiX6sIV+
EYPh1wQh2knoE8bZhu96bkysO3z6a3vJZEkjEjhxxaFb83DzgRE45jyuF0aVOqBh0Ix+QH+8lglR
eC9o2VI7ge0OZK3PUeaENQmFufH5tul+vw21M4qtqd5WCHdD7eeX+uoM8dEhM0wpasXliRucvcAX
j6d/kKvSGYkKYbqJfhBbxWJrxKXDMob4r+kiL3UIBamjxjd3LqfRhaVDY99BYLhHqwLe7PKGAkbg
9KThjbQWQJrlU83P1JIdQLWT8D7Xa++KBP+xbyFiAeXHbZDl32xBy23Hx/MH4i2CwXOrdGGt8Jrv
mKFjxW7QFxGA0G3F+Un1ufpOovRh3FGBU2+UnllfQ4SJwubCQ+Y5jDgEU5gQhFcDC9/FVh7ptFZr
J+fDfm6SwS8Xe9WEG1WYfs3pMSefBq9MhoGAORAU8w26Y316MfBQCNLx+N2wvxu92H3Wvu13wWSi
KxQXE+cwEKgdtrOu0BhzkL3q+DB7dAuUXBDr9+oWIUQPnRfKfOWLUcY0GfUL0UGWyr1R/KT3YlDN
hNkV5Vg8z0FQP0E8C7yjMC0D58/R3Xv8qCLpTvmp7e3W3w0YuWVswErK9gnRzjzXH+XG9A3gcdAl
HkIf44woa8i48oVyfHp8hMRxpBHpX3ysCrl0uNU+HRB7nTqfpeUq1y8AWIeg3nm5ow9oQlzAmS5Q
aIdV/Cz2rfbL4SzvNwV6tNtaohr4x8KnnYIm6cf91BiMDMtUHiu7Acg/5LGCOLEIIHQUCxukV6Lo
pao71FywuWguEarIOrvt5ZNPWnP8J7mFx8bbPhtxKCPtB/14XVBRG/+rFwYDjD1ctJvh/Wvt/6J4
jKyh7zoR6sofPyjkdXq8AQH4hVMaJo/FvrZQO4D+hyN6ccUvqJs9/LHwot7CstlwB/NIM8F7/kT1
uJvf9RY380OIgFPbaedvqvQGxvTobXVZA5MlrHAAmJMVeb1gaNrbWR8DE1guBEPXE+mRpJhalhFw
IQP0vQKKsthcfndZf8bhK3a0G2FkbSffOHMA9PEe89WsM7Rb5Gc7DxY8VmVCTuGUhplrS/b8sNHo
arW4riTY4R7r7/24JNuXr46d26nQF+WGn97W4cWqlqxrEYoWZzP5RUdJZU0TdhZnqXn4sz2gtURJ
RwrpR1DySfpd7UkgRycAg5FjCGe0pzKa9FOcME/foDQLG2X5bV9Upd1RVCr75jsU5fCKA98YJLON
otHo30OvlFZ3OLlLFfKPCSowH7mbvS7pftEH0o8nZfL2KsbnMHUDlohdRuHTVIgAwb98egkZa9LD
zmIEV7qkCKuSLrQ7qrquWTBi05/Oc7VK/QsP2O7JcXWuPiaCPmzlmZHPic9JiiGbtlvwIxkxEFRp
2O/FC1f62C1gzmvIRoBTSSt0W/tlRqdMTySn0zChgU6pCSfY2tmHCPCai6Iq8svO9oKC2Q+bG6bz
4YAAjg+8bM1z2rYOrj20xPjjinawFk3DFK2wJI96W6GUUmZUz2cNcjqlK7xckYVO1RO/5q/nvA5Y
ieK0ekbt6egcxuuTQRT/zLnRxP+5Ukgv4Q9vJXM8LQfpZANB6C0xKfgx9KyVRA0nsRWTDBtkBx64
RML6Ro/Kv92/Zqg/BlDIlv9wjZ2a+OoX4ow4q8QjAkD8O00S0T+NhM9M0TXVZVavAeEM532jVqm+
amZHt0l4Kz5ytGQ6rb+QvNWWVwopKmm8NiRM8C+hIuYJHhnHSwMzwlT7MKIXvne8RjKxKrWGBdMa
c5FeG6VJkNi03gHy7icAt+S+IE+8kQAKZByKUN1Q9jVA1a3SlrV1ijfh8HGntkXtNHjTzC4+X4ds
GHt4P78mmbQvwagX4fQ/HLdNewSbKx+vgZm+HoAEbGbQXAiRtQFejTIWoijByyXOdCDWv55Ziu7C
Ql6W+WtbG2+ruV2SSoYPow7iMsiARW0n/3Gg8p4mcFzy6VTYyGftjjMIL8Jb/J/ylj2MfbzEFUen
TPk9Jjyv9910gTVVlxQszNYW+kKYOD4X8fkfIgV+diTsUzVqSHdZ+yAIxrhmqp/0XEMUZxv+svV+
Sh64rTwGFM09RI9ijH4pVW91sAo1gLpxQOOFK+GVT3ril1+8cmcgPKgTULolYOUFAprEl8zCRj1n
5vNL8Xu4bd/ChRY+7EMvoZzjkhiC31cAdne7QD/MnntG5/KQ58F/EXbe0gEcyvlzWQUCbq8snU6p
PzcmFy8QVvO3EHd2wKu7dE6uhqBOeOsrZ9EDhqLQXs3LUl8wz+gvGNoQz5xtl0+hG4hmVMWwB5eC
cxsY5nsgqKkCZiqVqGEt/l+i5pYX7HULCIb/KWKiApUhkOnCmDD3B8O6VHR3VoNluQUj4hcWL4rj
aIvzfZclhl4j3GvuE5+9LFbuAmh5IFnIQRhYCvFy5QFoEvsK5/3fTZoIF0jy2IOC7nfkRUwaHO82
R35azcdH3KW36PRYKC59TSiRVVmv7VVHwtBdhr2+DvZZIjWrnW3cIEPEeaiTMavZ9zqqRcfPO85t
DDjUue+Ac2BtJuaEK1MDha9jEqYbTPqQYYS8zDbXiY96zhw6Ivl4jhS6TWgI/PbkD7vXLqLynTTg
lJGE85MR9Dt5/L9FWQlsHgzpu3bMzUNhCrwo3Wy2lJbcthiYMDt0VvyrDxvOGxunKBO+7PrBp1GP
DKo6v0V2C/TALWsJA3VOZVeh4yGwqmSYUUh445B93fEiI6YRQJu3v6S6SaIy9RHnDxSsCzsi5BHK
/rffxJbWkaC7HCpsl53zzzEkt62StFuIsvfHuTJQO4CCJvALqBUvz/UL+gzgN1X3UxACiPwwP6Zc
kx+tPSgPdm/AvlbYBsRqB06RxwBLlMwIaEvXzVkC1gYnJi+cDFQvLCUILBsS/x33MgFGm99mTmb5
A7NLnX8pZ19T44/rNJd7zY2rtWTaRnDdReHTpI9xT2gJCzv2eZUPPARqf57TzCVF/eXqiqqfF6Ue
uB0w9M2bEg/TaIVwqAv6YEmLJ1YTDoVIgQ1T+wlEhs14aBWO6hoMidXOgkceINCNRLgClScxrGQD
zo8BBzM3aovxW56PrHtqrwuV4hA66ludP5yOP5Z78ZlxUfNmNdbnL9RjMsYKSFKL8jJAjH6aQjKT
34dJZ1QyCkIiCcPQiSXhZBof4vq8wufLJwMx15nJYWcyntCj04VRBQ2yGX9JsldovyyRiRvKYhae
IyiKT3MF3KS4L2Ku7jhcmJi9Vc69LzD0LYxNUsxd/fiVFkAYjOXHI4rmsdCHcyZ2L1d+TuDC3S3s
BNjH2fOL1ODdG2C5S2V4GCAS831lov1OMwMsHAm5nYqNc/uwItO1HF4syeg+WaQ6fnucsGRyQyaX
2IaJLsEuOgxlc1C7h6W0scCDTJylu9n3gVwNEMQndgaZNVuIEwCCcIRebX64uQ/MNwVEGJCHdYnv
RYcd8A6hgIP/UPdc+aBHkC+e6rHFcinMdlIBC3iB+GMXDjoParKO/xmfGwXOzi+BEmCo/mv16NTi
f377YKTUt6Tyz6nxno1h9kM6Nh61V+dGmWvzJOeZGh4GEWpE3ymy/otVu3UR9LlT+sSi8NnjtYjH
5X6HrjvLsyJXvU1CrDaja8kHGvqcKVEsHVddJYLLsa4Js0y2nJAKpVrBB86rTMsZXzQMItQwUQPy
7jAMP4wJND4Pw4J/s8gj2b/QusdlypctfGUNpmT3F8ubozm40uaQ7X7qu8bGTnYjsL088DyyikOu
XJFR6M/V11cEpQY65vG9xldFvzbcfwyaBm9sWrVuEEZb6FwpYMIO6s5qaMhaqbMF4Ahntd30N1Ot
132xqWqhxoiYpKCGgMasvKWULAnYVABW0oEvqZPiOa3yIWhumrEcVi7mETXhyX6aw99TCxHPjaT8
broRBrA0vdGYhnuX1zPKHqOS49PjYl5l3p5F+0MEeUrMVSwbQKE7rJeiCHCBJfbXkYuAcJjvUBer
Wj99Rxjm64iRVqn/TEC5eHi7mrIcVY8JQq5NZGQArHcSVEeqp8ULNge5k6qIzaG0FbH88qhmA6pe
WyEQtQOqlhV99U7Pm2S34eMEIo2bGMd4K39MfmH4UHh55W/VDU0rVexwuYYw2PC8A0o0gKY2ZlrX
LbTQfmWqwjnlZObG7diR7cjPSjAOOXGrLUayubdM04gU15VSZZzjBTzJixr1r4a8w9DZmtRLnUzJ
ccz6ERAA6ylaV/yXhH4634MXdUZSJSted+y/iqrDadfUmFT57D2BBBLrg5jrl8G0/F2IzzR4onOi
9TxNn8pZ08bgzaMO4ve+rKIXMucCwSVaOlrpwEjglb6iDVrp4sspmWC9i0Ytn+wSW60RsnVdg/cq
8m773g+CigggWIdWe/uJHof9R6r5p/+2BPGXcJRTpEJX5WEd+Iq1DMn6mRaOhCvewxcLbKMjh2Kz
sC/0aGjeTgg2WXdfbcJKNm+bGt2h3oJpiDCPIQBJGgOujYCRTK5Ak+a/2Bqu5GpRtf0wemLzTYxu
IGh5ecFCppW7b0lB3uOF7T1/wVZTFyrWE68JfVo3H18D8C8HeyFtoVz83slIGm4W71taRDyGofUE
T7RBLgQJt8SzdUvwmWaLnosDMp5PPYU/WJZgh1qRqzPuxU8FlKI22JCerxckIEnMkeKWhfVc7BA6
YgkAA+j6IYBP72qJTRMqjdv1vWR3GT2uofHQ7a8F61Sn8lGF0vw0JkwHo6wa9v4+7SKRQrBMjx9/
GAr0AWefvmtOdPzxLgvfe1E/sCPwIsFtb+eeb5lrm4U2ECaTrUtA/0Ot3ZTWO8VKvimL2LLDfXP0
sHb02loM8oNqWE1eMFyj1vCb6u7aw6NJHZOaXCxuE1rLqLMyQzdwChQ8QIIk9ICMYuoUVtMuo+cO
qp9Owf5KPyjSfXwoZrdvb2AlNVgNtcDaKlMatPkhSWzHCZOaz/TYELGAzaWt8UKWCc/y0chgCYXC
5hGT+Cv+/oudcNCwxtYobJNPWXnPHzmO7sRgkrm8RIE44SXjAYyG2+wF6+cKuuTvv64vwKKbFRtO
wEShrnVoT1ENSBWnfRPZOBGA/6EMa9Fv9mDioDSm7Rjv3CDNND3NYhWeXoefHooinLeJCL01Q3CJ
ZELT10q/pcbtqXYUDdgO8VcMrSmkc1v0Wqk87YbqDfWKtyCAGqWBtzig8Ch0dBdAJUvDTp1vnuBi
D8ms34u91KOeb+2Fj4sJZine/NdJZCFw49mbpNXbYHFj8OW33q2C2uefXNN5gHMqN7jrxQJKuWn6
ZC33J88N4ZKiBTb6vIlEfRF6C/Evqv+eeKUW2LBKGV/AbYNbsvBSNHLJLzIBVDDH5UF5IX54VR2J
MEMVr4Y4hxumJ5RJ6vFx87X8mO2OJq7hk+IKBYXVcgJtXIEkDlg815KTeNhgIZdqdjPZL6cM9zJp
iYBQa1XQd+Pkb3gmoQ3GrjT+Y1NjLi/VNAppCyJHjvTJP56X1EwDd4j9apkDdRPG/EE60pi7q1LT
5xRbHwIkNKEAUdqBcEh7el4NvjZg1lKbioDr6/A5hO5rvZzHDwYZertyozdKCcf4rEf4jFjgosko
od/cbu3CvzxI2taw+ZJKbpsZddcMCCvZuuPWq1CYriwECpAiFX2b4WbG/5f9hHuFWll21cA7yJc6
8sVPNATIppPkgrLbWqwy6oLT++THp/DMlpIxL2Xv/l1HPbi4+ih+a4nTzcvo2RHQNHOtB3sV1izW
FWqX8t7UaeZdT7KTe0TcAvtgBHxipJJrZfUJCMOtt6UINCBBlVEjqPLMXO0FQ7m+TgYHwF7cJaL3
rJGy7ZI7r6LB2Qg7G2gpGbIcX1vpd7kpdB0gRyDENgjhtUBKqNWiDELlWbpmNpIvEFXgJrqX/mBb
ZS06rLUkapk50EHPYATEAypCzgGg0RfWBY3Ya2NEjM2LsNmksmlSVboVzyFxeeGlhmeoJlPmmvsH
dLdnWKosM0gVNaSuAyEYzI3ktaV1KNRKRUhO1uOLhZRTqX4FER2J9W9Yg0mRmO4YNItHJT0Fy5ng
FjbOuAw8n5EAzpthNeXIZJxMvIjw5FWG0FhUuKhOki/QyuWUATSLiurH0FADuWlU0btLQ7acvdyq
H1OpFqkPdGWoXJgIszMoCeWHKEXyaKB6d8CcMC9QG8uuwBZGh2vWrumV5aGpky1yguOkuiyKVCH6
T0BKpJMaP8jCsu0nttM9akD9J1QEWgHQFa8nqBX+pOKhW+e2/SCqYc8BDhqO/lQb5WpRkKNQLjqs
+xuUh9VfQNFYV0juSlJJPyP4HNupvMPDsp7itYoQc+1Z1ZZOwAiyvuFEMoQDD1WMuJs5GCMRVnOa
d6NBgNEGLYqioDaPGiKAzssk8R2Fvh12L5Agk5rVI6iJs3+mf/0KOuuiOX/52kRO7G6q3PR3Hlco
1x8IikeqYMM1uuGRLs6BZdxRpBMwHWY1Flv2cfzlpPHITcctFNm6BthRCKc52KqFrhP5jnH5vpVO
3yztLuUKEaq3gjwAD6PloNX83rq6md+zd7kaUug3nv/LhHlV4qtvl59Id3XkRw9HgmE+qbiGBVaH
nrxUxnVz8rm5CR8TK8dX3OSuv0UM3LHK7WVVFWg4HdNCsKB56y9qsWzIDAjCKz6Dqn8Z7RECV3hT
fa7MT2lw5XJNHKwLo1O0EcxmY815u7wkzoDXrM1JMv4Wr6a+LA8M2sGhlKLS5HRGX40PiARfY8sl
8KgVs/0XBzDiz4mA1iOZg3oPArPldzSdqcYs8RMrIPiWUwkV7MdUYeOqDbUcwgQTR+vvjKn2QM11
DQd4ePcqdtKIvfMM+UyIvxNcPEfKX+Jd54ezLkZUmC0qeaXcWaRTIAGS9Zi/TXxH4a1NIkaxgQ+8
N7MwnrfDgvo0i/buGlNRFXV+0bINEzl7HEEGu7UCWA0RMmKg8aiKOU81EiGBi3aLMP8bFTMXxQ+q
rKIg77CrQPI+ZR0McivL1vkFDnqS/UIjSt/7Wg5ImvLFnH8ZaZPujMMROV6QQoTZgZZTNZlICH4J
sQCMxhziJonwu4tMSKKb13eDVlkMVr4MLTAWD2U9xgsUVKW0uOvpiw+BUh/9Bn0yGkDi3R+s9Kjk
egjGIqsQIJYtwDrEfXG4ylMeaQ7tST7gy1UzqjMaciNN+ld5CWGBLOWridHRHdl79w4RLwQ6cUE8
kxcoqNKWVdGBP3mR+mEm0IYuSp0YlfBXZD1RJw//aglVNROfJVv5Q7R7ISqgnzu/FNZ/+OxKIT0U
7dASMRc9gC39LvFO9hf1dPUQKhCCAAx23QIe99m5KAXHlmNuAKZbNH4KwARJrkbOuVThH2lFnsQ0
T9tCh/UtTrn6qx9Jx9gH73bOR1LoDYNN4N8vYfLZe9/F+Aq3MpiBrmifL1PmxpqbT9xrE//jkm3h
Jb8RA4RkOSCAlMDqRZk9GF1nzmNpzWdHHZQsqVyro1meid4dD+cPCrDx+Lga5A1O6r3RwtBAt2Oe
YH+qzwQhUMTzogHyPrA225FI66B8t9fwI3mZKe59PoU+06trF7uIz8MCLwgTX1rYn4rwOQATBgXJ
XDBtdK+Gm+2krPwH5AcuhNyothXZ9pDnV0Q4Lrl7+no6Y/G6WC3+vRzuOrm/SLXSTI2vWM8p5FsE
cWbrXUZFtDeaitVFG9dwZJ9livcggLWC8jDPzWSAbsjEZIPSkqxNsXpeZkZ7vrvYA8w2swupG9Qn
AQEGQjeCORvqCF1t+b0IkQn6D5YIjNdh+fjeHhIQbUxbiyd6Ild9KBcZ/Mc7eCU/sU8QgaV+Tqqd
1yoNl8anob2KFeU8ystrFQPAG7AvX4vO9vHiG+RKmQqBXOlFvryRVxjtCaPCMC8QGgnMv/yP3a0Y
lgsJiBVgpOKcXSUSuyorVdCSEB2aD1ax4biHwcPt9AsxuThzwsRDRe5usl1C2WbeqsydvsgUaNm8
z6yVefV49Qf3OUZymb2SKIxP0bo6APJ+sTwgcRS64vadYuDjKFBc53na4CwIOvQ3B4zQTiNteuL5
w682kUON22bN/EkMqYyJabnRH4Nbnpm6r9QL/Rdao5fDC0R/RXmRHUat5YUlakCA7TTLEWw+1LZh
CP/452XgUVdUVzAkLbxB8KFTd+neC00cQHH2xvuzlI8itNeFGqxdPmkWlaac4Sy4TJ2D3V6WjnLs
QSvIeHcPQfWzG/zC/2gHt9avFLf52y/4Ul9Iujk9lwcs3qhz9DYpeqThWg63OuXJuFixzDLC6gP/
QsXHEgzxVhfVfq2IQlBob0QYpnMh14xb+IxvIGKAPXGK3eYyhItyUvbKuDmtWcgYWmRp75MBt3kP
Wd+jnzp7oHi382BNrB3Os7GXNFqoiVeUQsW5o9aasTIAZAubvwEA85sfv1QNEK7YpRNjmtyW6PnZ
GsbbyeVdVZWEs7+Ym/JV7cO2j+bBoJp5bBgvmZPuPKKChjHWEJMZ8+HyOuukchILHteByLCOfaUS
UUedEtcmLeW0eR//KWJkRUt+mBosDhFVZyCsCZuIl4Jfd8BN9rITndwBaTqPkMjjn9+wYL3xAhP9
oA72/C305ZZ1aQfDEnoXIqJozevIO0gjrAYKm1+c+k0LhEJ3KkDbJ3YheDPM4uN4hIjeWqAE2RvY
fnDIxVVZhD033dr5AipsFu/9Td/tv+J07U/Hqx32xYTGaorYA37NcUAaC05jUIiaVFL5hdgsykcs
NarAde0D71msfqaVIVcmyCRb9EMYm6uft7OA+9S3VxdCZ1wPTdN23CnaXLcxkwEwshe86huj0DUT
xbhnjOSu2kB6+C5JNooztcMHQBZSeV1T4LBoZ8ZJjWNCdNFH++CZy3okwN6AsUsyk++A5LRAaOvt
yy2fZdlUGOUD94fQh58Nj1heQorsemSdGvWRWPssf83cVWaRj4IORMnBJpeGoFTYPQ3mdZjNkbO9
6Lvn3mpJdV6ZtxEUg7V18/pZXb7GVI2CcvsnFJarlfUtjhDMF5q4+CS30THQSkcSCgxJsSx0rn8u
nmM3959WLSlDx/p99MbLMxmY/Dk8gpP0YDA+8VKIxnbWzZhGRA+Tqv8NkchXygJOgq5aS0y6IDbY
IEO48V95eibQ6SSZdVmRx6fGo9xrYIZ5eQIorq91CRXNVK90LKrjyagHknrKHDA+dAk2SsGA0XOA
dDREamFb7NPaQsGGqgL9q5sjWw+3ZtTlrLKBcif2U4QmBReeZdoJKVE+4Gcw25wGLU/0N+YQSeJj
ywtzYdBzg6697/h85ycUOclWIGHyku/ABI/+CrDu9P2PwY2/KFNH/7RIUQSQD/3bxSVo00m+KbV9
zkORYG+wqvzhQKC0hWa0rkYBjsNIA51WEW9PzT/eEXX/X9r0td7LF9tRO/I46AeRHf9FR3VN9bwH
wJYNbrghk5lcxJuIoFPMVhZCAOntbqLWDWOtQ9mMs0PIe/eUCXali7tAJdvTdVWhqSA7skeadulw
cUeSKgw8Pp7aKdBvnyGvBlXaJCWgEQeJtr9qxiNmkhvkqXopJ6OKC0jmkzRLcvLMlrnxlKZ8LLDw
lAIiT6+4PGswG8CaQ0v+A+PPvWbC01yh0ssD9Svr/l3TnrvTJEPO0ZREjEji9yZfmBSZ3+H1WSDQ
nHIgc3oXqTfJjS57wj587dvMNw/WHsfgXyMy5RyesKopjuHHm1dxx6TRhGDrDWmHAjOVdnyAFifD
My/2htZWPMBH1kKbZC7keXrdt/QEX0q/1nZ3hVJ/zsPa8MqFEIIusbMO+WgUElDaW1s6M2qbSoyP
p7eELHaJTeAyIJZjEzXMp4ftKR4V3Do9d0QY1Z2SlWXmPpR7uVHwYH9xaKSKQH6YUv2V2kkmTrh8
7VFWmkP5y0YbElgQvrXmZENl1jt16YVImRJcbLshV2DpLbK8oisaBMyWjTFunQR7U6u8YzxqVU02
TGy7hvHmC7+MpTbHPCt9dOd0/pSwffICZetNzvJtqAuiNGoPeaaOeDk+r+pS3KyAIKWw1vXvPAET
DF4QW6HlxGzgoHRzuAgSxq/zz+WvFcFrWs3FutW5SBqTPy+JWmJj6fXH0JjhRPWyE5GNwOHkjSjl
XfzYhEy12cDYB47nXJ4zgOSXzCheKzGvxTku3sbXeDt1k3OqjgLYBhOmhlOis1HRZUs5tkxGvxbe
a/1D+KOR4yE+AvfNug7+89deMxloaOnn44NMuTy66VsQF9Sx6MeEwhOQTPy0oSe0N48bUs9OLgBK
lWCHOIwZhIxNMHccnSXq5U9rvPStyhBwmFFvCYVYcU1FQrFuwUgHVH7vpuIPqiSH62e4ZStgtPZ1
Y3H0pFtCWg7716C/8LZJg/dFiIQtgyMDZjkDrgZlnl4Tf7IOzYVsxISgJLWMfy3m8m8kUH4YMb79
JVOHpbTSd/RxY1TdAfMnEA5uZVmNcSqYQ8lm5YUsYkblpZnKuWMjrUkgU6P1CPYCMT75SASpJGz2
agSp+555mKVbyDHv44Fqwkow8ft1lgY5LDQ2mGAXmcess9mUr4tK7nnNn4l6lGBeqIJQq9HKwt/j
34XnscqdBK54mE9ogPyKMyFWn8Py8e49UeuCNprHKMDZa9wVilubZeBMSPdOjNuUoY48Oz0iQlXI
tpHdS9RdQN2TSSRVR4gwBFx6yQph1QW/sw8TyCIz18aAleFaiHqgv52Y42KkMp3eELmmfnl4UaCN
jl1boSudvgcx/j5FPf+h6PCYD6684SzXG1aPJhudq0ujJsfDrE9VA3InGpbvBd2H3IM7TVEzcv4o
NW3/CFTEFoFNH65HFLq1fCCnYUFAU2gipNGLT41NoR/xDBoohrbMsGvdgQke2nZ/5QLGOn5cjTlj
tZnY8OoZ6zabnIhqRGR/DDwELp/qpQctxkfEdznq1DwpnZNT8LOdHtluMcE1po21XHoDxcDvoDaR
GU/e6jtP9+2oVLIvBybXSNCoLpDP8lMX95iAdOpH+x4sm74nAcWjf5bP7rhmEyhdE3Ad8wYCCTRI
KBhKdqpzHtriUWsOwtocU9EfXLeLykHDK4pxlRUq4t5NqFXXXllpU6dmlkWmLLYu5NAjaLzcb+Tz
eIJtC85EbATHZ+e2dJqbaOZhLXLwLhgHhImkg/NtfWAEoxt6pRoVUwLZlIXVS8P+VOZsi4Aw0/yw
7CCvPi71MvrW/WtUKp1DHzy4YtGx+4cQNnQIj9QJdd5QxpUZO+33iq9/4E7pyECRcvbQVLERhMDs
4NaRdR/da+mbiHC3htzAfx25adOaT++M6ZCgHnDme6hNVfmu6F9nixVwOB/S4eWdmYwBcBG0VKo/
o/kAjqZA3Oqb1SrRmlJp6vubAdZOMwlnvtVcGYkhwMXovHpjnVs5c9k1a0QsYkyiKOifOEUOShcu
Eb4LvsWOd3jbAR60xDCxE2XxcHsVRf1EbC+pz/Mh+t4WFUZK127jQs4LV+WvqYc6Ilt7GQVBev5O
TFB6ofhWBrOLzAk0VJi/Vyaw2RbmNPM3X0GBcDd+yq6s5+H9R7k3i7LbahPEUqm6USIR7p6NtWTo
jBMCHRzi45lx9d4zwZwzIZg3mV7+bipSCwUKiGMAyHvq/XDSQDt1KZd9Mc73T0+Vpv3bQCc6xHhl
kadyJrlT6IH/z1wepVUzprKLJEBTmzXR7X/+WGPKIi0GkacUYHW3QkogZ8M1aC8STJQi/KRKXLk+
ogvzNV63oBWIkj+SbA1PqkUHU4R//16iHyoURTrGV312PE/glFXUxpSJimNXJsPLXvTlR3sbSW/Q
ExCTKCzmp7Lx8s4299iq1/WV7zL8qYwNtyCGKasp8A3FVLmdryzk103DCCrkU2uqd8QbG9jI599y
D37niGHOwqJKlkis1w3eFgx6FTHFUhcPL2SznxrnNcG//INmbKj7yHStOBZSOtEj+SKfpA4ugxi5
9L82U6aQECbz35m+u5IcPP9uvOPSorfMQslZ+08Eiblq6Hov443gcTV5H2nejAA7K+KEIf3t8eAa
wyO6J5DT8e0DMfeyhZTNYxYu2X4edZ88HDqs/ViGBb65ixZwgh3iDThaDeOEdLqyXR/wqiZ+s/KX
0aTFrQYxmV1pece8xa68X+vIyR/LvVUcVR0L89i04WC75t5hdm7dIjSUu2XZqE4yx9CDgv9ASz/1
1oMOL0lhx8O0K9e3K7RN77pNB5cbvCHNcopnGOiQEUMjlXYUwIPyvo2/ex4ezgwyZpaHBOJtVtl6
VJKRvwQ3J0oxLowZ/vtVHpNHKezLO7ESc3FIzRBh2h7/dhng/kzQsXoMcuU6k0pUq3RO/wJtmTNC
Zwv77Zz2zcmjEApNv9IhsxKowO4Ldt3sfFrNZFrM/Y/YWDTDxlhxrgIPy9rOCYnW6kZI4Dm7tE6u
xjU12eM0Bi9cmQfiIUhjF1GMs6YVCeDVBANKZ9jhBPX4uw5s+FIZAVpS3Xu8WOgmRlAqsjcyZwVH
iydKRMX5zzciduRGGq8MlJq2dTge4BY/Znoh42qjrzNizCIVVlKQW0FdDxeh48x81XJE9lr7ogRE
Fuhxf5V0Yi7GobfzYfC2l+/cZKN9N9xjjkF5Yj2DKpWsxZQsIQeO0DAxjMbGfZkRpmFFsi6BKKlK
L2UM7fC7S91zj5rojLuri+0Pg66ynIncJQFpuS0BLMXckIldUeAF0BFWvpW33y4WX9dkMQNO1/ME
dpLi6rsuUabPsd7e+cxRH1T4qLfwEC7DtCHSuR3glvq8Vz7qeDKFJ4CkOo09ugkIHHezB51ld8iZ
bzqPsWRRMLtCaayg8Qr3g4fkmSzkQ9ovc0mOrDrBpa2/aRgiM3ArjO4pLdfwIhhFRIDmEPC0U0Ks
K6tAdwszgjiOvT8xcS6um+C6mo4Pqn6/r3VIM3BKJK4GsvjZayl6HrAuNtslt+nkpwqC1XuRc7YZ
Z8qZ7OCl03zxnF2J6tcFl5sg8w7haSlKIOnVqvX0k8U/e/lE7eTESRfr6uvjRJktt0Cyzm6z6gE0
zrOw+rroZyc99BlbqCdLVkzkRejwAgz3eouCnsYRZUfB4IR9gizGHrt/uv6Xc4TBg4woRk+YcVSq
rboCELR77oC2BEDs/zOf2s+eRlOi7a8LmCxId9pRBz3xaVxho5Kxl+/FKndvxWFa0kyqFXe9sXGF
sZZPk45EgxtYAVxxyQ1nSY15XCWReuPfhVvvUACSYaJqUbunm/Q3QSyccO0MUDlklVmFAgufsyPb
YdU6LFnx8qfNGwnktFlY5pRX+okn0s8bzjoVW8LrOncaZxKp9WC0YTqUBe7Gz0Ikh6gLXf7A+VZz
wXRDkLCBu4J/bdZjoIApdpb/peLNO/FkJoXk4o9HXDYh7OIFY3LmlMiK2JkdKF7xf6rsGmvE/ayi
uijpiHana0HBZdhN9ZAktenMAZMZep+BvmhxVooDox7+kUpsUhjI98aZiCK6fcEEN2wZxt+heSeM
LVcILpLYZP9U9/k7HWvm6iQP5wUna0jNto3nAWhcrGg6858TblX/MFntIA7z7e08va/SnRPR7vXN
fcPEUOhFTlYoDWFMC8qqpV2YumNb9Y/0gEHRcDTmZicVvqn+j9I1hEGZ9gOA8v46WLBfdAl674IV
YcIxsM9tjkx5O9TCN3C1+KZa9tEP7c3CkegNb68dO2hGHamCEZm2uTihGdbJZ5QqlG5ors1RqVTx
qG2TRP/lpOs3C5ZhE7X7z3ymo5ZjxchTMLwZfhDBWES2pG9iNvVvIoeAgROPPkjnEZ5GorkJNwGQ
bK0BAnZl7U42War5XTQO7Kyhiq87z33ABYpL9fHZAR8r2BSDZSlEaz/1ustaTXjdKDwX8UDJQTNW
XyFLYR55tUBzK+6vpIGdD+4sONjTIAFFwoek3wXtAQ9uMfVBMbQDRSyx0UoGGkXB1QmcxB35dAt8
G/z0U4MyBEML88ggateVwzIg/+pYXap26bFhkf2k4vjzhgt3z3NrBcgPMPqLnojkqtfsQKCQNOKh
iyeCGEtR9B1Pgi+EalPBnai+CEbPKCrWhNahrikk8fRKj8GSqxEMXEqIoD+RZyJ+K3nA967mAiI6
V5rhfoDzZBw9GY8aNp4HW+/gTpBRJR4yj2v5QnOVPhK5XWMP+15qbZQWuMHatBJRvxbzUbn2vsbv
9L8ZgUMab3X7CUuIF+8YvAsIQAPxnoEJLYonn/TAOUpFrBBgmJpqzuFryHHY6l5ZhYBFsfJnEBvw
86caKJd8KdXzMAdbmGCiCmRaUgtz1EIvEz087CEKt3fl/jNZOMQtLU3htjHOvNJEja4tCYYVZoBK
obZnNsc3DJrAyKKF0SxLX+Vau5lCc4xCRIEpljA+lbBbzjSO6+DhHUGHYpLv+mBLGPrk4ibAuQpA
DNaR8hoZmIrrxPHrReFxSb39bcDAa4apZi7TjSNhPnyjTkI8jFE/nfSl0gbscQyJQzSnVuu8WWkk
LcGbZE9eaNlBPd2/y4IDL886LcyjGRqBaQ+uQrCOaFPf7zAgmXRQ9UCw7PglSlNEoiRzNl6OyvYx
MaUcwSLaLsqqFY/cC8VW1cii0oSNvjTB1XlRhKMy4fIvWbYJ9P2V5VIAcnVUCTDkzIbKRr33ZQs4
3/NHR6cbPf8k+AbQpdALrdNfgxFhjCCHxrnspnC45iC4xC4SIPHQFuntjeHdLBuaMHI9kTC4etob
sbnzF4nXzPUlmNRtm9hXPJmRJlkKm5HaDEkExORoj5Ht1I1URnhdpjl2SV7uDWZruI4lgj3aITAR
dVt+QSblOCbL/hA1Gz8Hwx1a1vGIZwozQcHWs2uMq9QAk5roDzoDz/CYJUs6ZT07iKvZiWIXOmou
Bbm2VZtlPqU8jhYVKwPmxurmLMJ+Kb8n19qmReKYxhnwTNJmcevYCn1nTAtXbyL9B2DWzR1pvkKc
UqBksXsU4YMijjg1nbwAT0p6VcFheoGpLA2xgIzg0j2OdKfAplfLywdzlK15Zo3ClKG6uCbDhCsN
yDMSgp3ArcvS/v1TkgwqfH5Pv7kfSpwNONCEvu7xN0t/wM4hK8hEh4bgady252phOVRi/8oGdaxB
8TxICEDbmQCs/X6nvHC/8zmIx59kmFQSjHkvrUD+ve/GDoRnEG70NfLbA47iSEXwx1K3kdRtIBMB
J55+wJXfJoqGJrjQGwnwjKM5GBMrpz8opnUOeuBmG/S29bgpjDQb7BzNGshi3PqPQ1SAEshNSacE
nz7SHK8E2oO1c787GzrP0RSqjfUqfKUbYQQiAl5oL2D4c5RQq9CxIVOxNYMzSykkkGKgjTHJQk2o
TtK7a7ucA4uy+nT7Y/L4KinGsDMuKo4eCbllFcZsLINe1pPk1OC3Kyg0aPac4t/mp0aX8/jf/1NQ
93uCF53EOSNdVDMM1WW1RbyjVsi0W4+/EXKmF62HBRJamGxnksbQhKetzeUOqtl5BaTuAizCSdDM
mcQF/QvDHSmznuSz7rKmHV8GvEGk8Cxfnhh3z9F01ATstifVYDYPT/HWgFVF+lNLVEbNuAzLUBbk
K1zH+jMk3m4fTidwZl72cHnXuxxhFr26BpKWeljLuDq8ekXHg0aBLyHlUVf2tmtuzXks3Y4uB4fk
UIiYCO2nET/zrXNMfCuHCbRjnEnAcXWb2s7HkXCbr4jFIbbOrMKN/e6k+RqgtDbp9nG9Z1Ax2/42
pQQlTY9NWoEWonAr2CvqMZ4fzvWj6Fochmpin9qNSehV+1AACC+mtZ5VnWadsbL6i96A03hL72+i
aBD2XfqfQdn6/CYlP4aLC9rXjPM51yshwC1d3aDH90lRJYcP3CJjZe69gkY6wivoVgZgdY5OF+43
XIFhImQCg4Ucbcq7lxcL/6uzKxUNaGbec9od5Bah97wooKG2NfZWnW0nFR01GjWxuuj3ytTfXFkn
F5EygszAxPa4XRn7W6TaY8DMYrDn2yyVk2sGQbAtEqzMFq950IRJHR2IrCnC18csId9el+h1RX5o
nCRamM9GoI/nA1ixIW5fJ1tOcIvbXSl4/6YVB7QUsD5UXSn7gftkHKcInDZ3NyWkP2S2nE56bEpa
ixbPEgl24b/TrxvwkmtoxBkbcJ0Kt0mnHWUZhoKUQ5HbTawODSkp3mvcaJp3V3Gj+ExIGMbCYgqN
cZQLdyIB1wzdPdriqSQQdYzJh9aqWtxoub1sRI4Mi32Dem9PCjQ1cd1+ohQyHdrHEj2pWEVFo6O/
IPCjh5F30VV+mMiCMYS5FOSlCWQtu3ywNelP03gXpkR06eA7UmYkXFZe0USPH7nm2XnWz2YIDrQd
+t+ylq8qbk2Cip8UUEWGotqZCb8cP+R9T7MrHthOvNlsyVXCGSr+icZewjV36zSyp13GloO0ASbB
96XcO0JcBrjfD9bpFpYLxiphZwaZXKeF84ExX8M3aqQJqUmt1/JBWmk4eQLjyBCLtqz60KOiZc0t
xyvO7aW41HYrTXurSUbJa99gT25PsGD5Cjn4NVQ1sAmGRblS6wGA8U3NQh+zwlVP/OFvWkXFXCso
u/qAm49t6tPuowxAUDHvEj4U3Dom04MJlx52KQU2DdhZX2n329PY7Qj/ryW2HwAV3Nd8NqKvD8RB
piw28EScMDV2lSmS/u4qBP59MAYFWYCsqdPXekBg675f3MpV2UR+sOzbOS1F+aIp4EMvkr1quRTx
wprC2QYlDKuoNkcLeagBBbXqqzjeiXdorxjS2fR9dZU4AMSRYO/SZFAPcIhHfYwULzEK0O8/KbGb
V12snQsZSIDRnALmRAssqnfMH+G3Tqr2AtOP1REi7m/cbMSAnbGJOtbtqJWaIIT9EwD0GsPmnJrv
xX58Q18EmLy9dK2l1cSpCGA3Rh9g38Zy8jUzL3hnML+cYyrAybyvbmxKdWJOpc5D7gb1QA/m54oV
lizPLKVWUzbJJaPbzF4z0ykz5qBMRoaHoc8lC+gHDHNWv8o8wDSC4B0iqh0u0hndBdm1rNFIuWc4
07RHABBIRLgrdkqGGyFOWEjOu0PTv83SqaqJJUTVj6xKceS9CB2jklb2NsqrftuuOE7++jYq77sP
MmRpZ1JW2JSos0TAYsg6Pq1aF7RK0j32xwunbkwoaq6NsClnsXpLkkNs7ufa5ChastGzc3ZrupRU
LDtbarUgcV04SpIDI0eiHwFYl6m5cVusB/AXU0yAt+P15fBoSnEK0CtV4IwMEdmF5bP6gsyLPYhZ
5hQ4vC5cpQRIMYjwzhGWfPrDeUb+I59WV9wi3Tr8THGxKtknC9mdBRpayOSUC25r4rUkVcZ2Pelm
gEfTzezeFQfbHkXTUjGrUb/9+az+KD2HqtXZEv4JThuUwOvbI5/O97uxgEpi7WM7xLMD+0ReL8qG
pNwYbhnfHu68HXzmiR35YEdKarQUogGQLLI08JbQE6OdhtlNxiRsaTtwzUvcgIgE1dtqKtc/8Mwz
EC/oZG+o8SXgvAVIxLMwxrGJaKgFO8mLTq45mbTwKx1WXkfeCDjzj42Cj5dANM08eG6NJJbtWc/W
CkL9z9IaBqGODjAqLIFL8lvtgCyB+xuJ2XeT0XwCJLPnh+JqbH8aTbR6SECOqgrsUCOndYPqNRTY
HD3Ou8ujtMm9lf3G/iYA4ezHovNCaz3wupNihmubwd1XZrYB5lSQLVy2pgDAvJkZ0nRAK0HZyhzz
zxL32rQRCXiiqg15cOr22Md2uCQgshyvxkFY/yqoPs7crbkQ+CzLHm2akwIka8D2FhvGgFZLk44+
dEwuu4D989PyZ3gZB/urNnsF8qqnExHIBxKMnz972PgC3KI8LFmIaSg6U5uNrs1T+EaGo8H4dRs/
iG01r8IdK7FI2lcdFpOpskU97Grpha2I5niHv68welcn0J4qA2UpVJF95+rJ1PMqd6JcdipNU6ey
K4iK7kPo2h7TKnQfxLkwf8Ma32dwN3TBIfnN1EtBuypGq7OH1GO8NtYkFjeP01m5n7SUaYk3r7ev
ezdw94txHba3Ta9mCQPViTk/y3Fv12fVgNLGlyDSuP6g9A/rIrD/1U0Yo95Tkaf+5ZN27gLWxCye
n9MIum/xfA0vfpiJLR8pB19neT73nQ5EZAk/4MGfGvkF1O/4tStiUDM0WDXg3lCeTLN+Fqdj/C4V
/qaUGe0lCGpWIILDQ4z7AGpMBCitu14WC9R6A9nYLSthJY8+nsM6sqD7OySVmRCrQA/q2yOiD4RK
tG90LR7zbBu946XR5LeaU3DUWfU4C3aTTvZRPs+f0KO40L8JfEZhX9kRqxypkcN2wi4KwDtuNg4s
ItEw6XzXLrVk6TJk2Gbk5/7q7kXfRoUPamAmLwJjf3qFnu2mB01laNbVmcUBa/MmSUOUNU/WLurz
/7i702HQgfQRIYWVI4t05QCWRcDcftRGD3XoycMqu8srOXW7ITJOUjBPpbqzw2rr27xxO7Q7Som4
+CGh+SayEEsEE+jAHcoAiVk6Q5LpM1mVcxjD5UMiQ7dADixdVH4rSvQb4qjQYQDeuw7l8NrjlR6g
HAidFU/EtFBU58NVVzDJEXitFhkS/UWweBWM5IQeH/nBKwvEgxow6Zz6APkmJSQ8+IjSrKDrlEj4
NipDSHwG9e1zlZNVrkylBzKG/ctvMSRHoRPS95ietZUrUeAqPxFFtaTatSjdrVkBQptQ4wTmDmBP
8hqK6VML0OyjO00o6AL9mK3tbThnAU0r0TG46HvJss5uqvAcGcCtQjfiGencA8qh224zFTozxExO
hpjmCRddYa1k5X/vKF04p74Hq3lyyzVOtN+CMd4tDqlrmq5+iGEAlg0hxoO1pRMRRkDvA+Wi1dMm
HysWB40bcN+turwdoPxte6Z6bOR7Hnf0MH5xmFdYWIDuKvf7H47xXugPznpEoJ19ohOkpK7T63vj
c6VgrB33xp7ysqizpls126h8oo5CCR27L1Y5z8g5+lrfxVDcYcDkmOiadfTMDQQGk7Cgk6BnjDxj
SK1I5voT/sn27uT7B9uMxZCff5k0GVJJrBKTSOKOhb9uY8ix5Nk4UHEUFDl72rHIbxAYthqP8HsX
KUj4e5aVErLJKC08ceWXdhDFOcqtKshxEgX4TO1LFKISm0O76p7QTetktchWTGZE/yszRxT2s58z
esEN+4yIRlkpTTivNN9NdtYec6KJxMLLZdvHzEDuVE4AoNuNfhyHIjoW9Fg4qYNyjd+V9CKi5IBg
r8yl7zKO4aJos0PTp7bcDNbhr7vfLITRWG96lGBhqMagPk+fnIlZ9SnIEdJQqQ1siHutmVQCzTAp
Mmp0FWMarpnBGSMxmdM7xte+TsP3I36WW5pMHjNztKyVygLngP1GcsuB6sizi2roZO95awmeyu4J
4lPg4YoDDsrbCihVzAljWlXCZ4Kyhd6caOXQ5SAYYz7d1yXVUXudmt42nuJoEie6A+d07owwP6Kr
5OJ47BzRXaQxhQBeI/zQ//gw+aIN88qxh9ulDfO1JprdHvm9axYRv/n4GpQZwHLEFTT4nZG8IYXc
+dRv5g4QYAMRsOKi/kVCQry+tgd8eTrGaHRuIv4/U41zlroynqO+Sy6o2YRlkC0okz53F2B1wqeG
Ex/37BNY+oFnI5vIMdbzP6Pu+YrxoaBwBBYV49OO35i2sLvyZUpLKHJmgxIz2M1Qv/hden4VDwCW
gr3z4GJ9R9eWXFyN6BvBt5vVAAXlMA2Z7F2x9oFh0SOXtv/73VvfaWdVjX+s/UDSsjlTQPiOEh28
bPoR0KQ0wg0B6iv+OUZrQqDW36sa7sZgVj7NqYrzAwclWl6UzhSoWnC3y+Vh1mSq3bXVtgJGa6gW
OVFjOSegOShTOMaohOIGTSyvhb2IIQD3w8Sua1fWiuWqJ1bDyj3ZiZG+RcYmzwoXhf23lLqQCJbz
4cVbmM/AlZ05JhcEjtPa5TCsVXJgVWsB7Ev6mQ8xuTF/8wKCdK3IDKaGZrlsU7NXFGQaYskGwLdG
nwPDrPdsbj1P/2j/AnUnGKKGd6DF0M6aWzwhTdBJJ6TdW6JXZFW0FH3PdPSIkEntAqG6eN2JdJEI
TE9GAfz9aITNfkFuzcFwbooCNhrQxXlG1OdF+0prIuK3IbyDpdpYhrUfgwxJeaLudiDzM0WhkyBJ
iKPF+OjRGOCnj+TjbE5/fplXCPG3UIKkyrcpz2lSPsLqkeoCZkteiLdKQVgVOYdiz9zNCKxhi80Z
aPUnDEYdjjO6qq7H7HqzC+ra69hxHhQMePPT9g20u29MqXCZz3NB2DJyQfslZDseKO6+E1EaLif/
8Br+HLUMX1phdc0DqjyqpxeJeEF0FIjsm38hJpiuIafFuBnfawgY9VwZXNsC8buabyDNVl/G+4T5
CEIhUQ27d58WSPEwwkADiDh1cPhHojeJZDVdFJJHGADh2RX9vfUJk392H8Cdc6CYA29VKSTPIFSw
NtEOEKw4SBcwEX+Io1AYQw4TBouBHuPhMNK+irjaH3uw5IGSa2oo4CdqD8ee6ihyQiExoyFT9Fa3
hNRwW/XQNnmTdHO6ZnFvWNBLIHsMAnZRdq0w7I9dSgXTW0mF4L08QDZl1zwo8lL01yJrF50mT2HH
AK9ZW2FCLQIm/h9no5Ks5sRKgxL/U/NoZ448IpkedfQpoELscYW7695CvEEVpQOkI7imVOHnNIN8
u7uQccYau2gjUPe47Rljh6pKgGtUzHVZ2PmxX//lmmiRIGnE4ya+35NvXAFnsP6FB9p2VrYHZTFk
UQ3Dog+UnKdacOQJJPWLIEtx2CznLK07Uy6hdeA4CvkgMbQsDfAAd53+YZjCHci4VL5joy/B6ne9
dmFRBRUbUrju7nIo03BygYcLawYjjsgR/CIauG8bB/BfpwGK5M1Nksw70XlsCLUFNwecm6WYQr7h
qKt/c89Te2qWzxko+cWZ0P/ta1XmBBgy4c5DR4Lyip+tnAn7GOkbPRxWyh8+7P/fQO+L0S9KSere
iPTw2G740tlM107SM4BRGL7bJyXFKTq626Siwb0mzE0bc0QRhnFnndCg9dTIdDLbNvrdZYtgCLDN
Z+yBH+3xL3mV/crlaCXRm7BOBIISVyIt1v0yYny84RHNSXZxuRHV1UEDXel0sqNWc8+5UtlHh2Tn
iJ1Nz8o8oQAM6WejAzcSNKKdq6gYp0hNEHploK8hUTTy28ZXd++Sax1fIt/exWdMclVbTcIIpWpZ
SYyhPaTqTIZE9CaL9INgJv25cqgP412vIGvxvWRA01Xlg/3mu7MsdKTnFrJON9E9cnS2JctxVs8a
iYRaPHPcUGlfUxXkp7GZAxcrWZAaOOktuAyK6SRSjkEDeraSck2nMI6UJN/S60SliWI1viw+c8cm
rE077IuP+4Lpx1BwhFJLM43nSVrRGXFcEC7OTelDfzAFdtt6dEOctcD/W1ljAncqRIvqaPR/Apd4
x3hJ1Q9kq45uribJB2KqCS2YQfGvktU3gmxKxsvdK8G4n/KHGQo57E1X5WMYj0BXWkxcJB24pAl0
9giQEGrvoMGZkN7TyNYP+J6WrtdFp6c1naOWg12asH1msxS1nGOr0/AsGXu4jR9FibtTaTVBmmz2
4brFbcg9lj/FTx9j63uRcy4Cf37NQXCdAEWOvQURzXzfPJjMMFp86fBYpf27GRi2vNmNifvZLTs2
U1wBkRx3E10XMZnKyTrWxErJ+HHnuPISBD66kdF3JHv0W8J1QCp5tumuGUgx9A1joOfl6WHSmZAo
6cY/ToQrPxwJy/M0Ev7nAoHd7dHTA3JvA90AkDiUcawKS4RNWRl8oBv0Pgddqw0eIz05HWBd8CCu
ybM103frICJXcCA+bTp4O8NV5QZ0xap9BUvK9hTdqgJfhRrYrnpMz0Iv1stLXWT4kbMYZhPtW1jr
3VzxFXhR5pOqASsxalvZwaobJgEkj2LyP4b/ONO8HX3+b9aeLnhA4nnr5jyKUJmJveAbkRNzSO1y
zMFL+IKW8wUuYYPOKkUYJbXWvk7z1rLWGxZIbbAm55kuRwqHSdTL8uw8GFsTkxuQlK1oJvbZh6Xy
JbGEjGgLDfG91gRJMe3WnG/30110phSfsP7lMK55HFm0LRyh6x6QdkXlR0jATgafR8RMcj9id4gk
il8ulY9yK/aULgY595B5B4H01mTQmjvvgzKWz02FVn9lQerUdl5h0NPmKGINNL4257sSAz2DWCbW
5wmu7enLY6t+YNdbG6rHMpMpPNyFN5mMc6aHTi3JSFrkSIY2k+oW0TMKFC23PC2MJ5vkZqGuHyrx
LpgbYzFtNQGnS5etRBivQTHsYWcBp4q9GbLTyhY4qHBIdyRG9p0GjfSywd/v8L9ZUgFXoINam8e5
ait82rTUj6e6coUrAMzA5Uhj/bUCIdQ4nNM9Zwb11Aa/5KaoVo5QAo92XuvLeNPyVAyp+77sbg/T
4hTxtU30kQerSC4LAvYKLg8JTHfJBTj/kZhLL8+lP3jNHdGa31MAatwrITn/ghFXVk127+J/X/W9
naB6/AjtAnJq6wuE+CwYKreGqeQoIe+jBciROUi0psLMr/QYK41HD0cxN6dFSst8k+/MwyH+7zrE
y8B4PczZxNSLBuRz+FvnMZXCg8GCgq4h+YlvoTkmz2aKYvJh2thrXNKbfZqh7iEqxLEoZ6Lsj3wt
xlr2gW1A73wjXM5Wu1sL5wdkI58VSDAh8xwYTX80dj6wDtYpZ8mZWzP4Qy6htk9aiGZhAWGYcaqn
QUErBrwC6IWjTIS93GB7rgl+GBVcLdadyZO5jlR7fAep6CTBiuJwYsiBUCxVc5t3rY+0F/qojg1x
t/9/34uR/GepZ7vrYzHHcCDtUOcphez+6GFzP/CAML29A6q9pjHU2M6iu+fFZRcwt9qG78B/t5d0
V8LhxJ30BfIEAPY0jJjAwgA6XtVX+3LOkzlFX0Drvyl4bzM8hwcvea5d7NX32ouxPUjgAf1hiSCH
pZ5djiJBuf3VA2x/16pxnx7G1OEbkbxB/VM78lw+74g+0zp1iofAq6yO7sEMalUD+3ofzIpLonw7
HNdZ2g71QvJ0toiPPaDLwukNRGFAfrHSDDVf5EaVgSmOrlBdDee7b2oeMdlAG0jVhB8wTjuCSWEt
WqRecWmdWInN3NZSsyN61l3VmNADTkJw2kmZslyJnC1TGxoMDdWQIZezprPeBFPmTNG3KOLJ4kK2
MrzrNAi5pewCWF0rw1qG7aTRHJoT9gFUa++dcO3yPfcauvofl4nIg1AVge594BUE2JkQo4HBzOm3
Trc5iiznwRrcIlxi6gIus/v+nyrVrERqf1ASXMLBbkp7lpTQsQ1qq2Soeh2br6LuqQw3tDilKqcj
ph/YDC2BgrdmgXPdyt/yoW/9jHEsVWKKV3roqZH+qUdDLtXKC4lB4+BVtuN5RhntmWfzzjCwghxD
9z3LlfAf4mLMDLWz4v5pjksQ+aRecFnwB8QDltpucIN0Sl7SG5x/CPhhd53Rf5aIjBqh4TB7aDbE
J4k76wnmIPKrJhf1L6hoMMSB2oYA+o/HW/XpENog82gqM5njP43NCFzKiDXTyHQgBiTGaE29MUiT
BGQOTAYBPES5L2BTbNFBMZNLQ5E9FCANmaXQOKqgr6hRNj3U9HEZsDygCfubg9M7I1KQYQUPOsYg
51erhzJwJCNsLy/7qToQRqyWrHIi2T4WU5Z2uIgzYX7qwuH/EZm4dVOdOnB7M2zCsyHkJn3tOzOm
7bILkMpThzbS2i9QlHKBDwKekKD/mOtdGh9q7YExoNQooebu2FNyOiGlWR58ZvP8l17s2tuN0rge
StTqJI2yQ//6qog3WzijxwO+NXsgt3hc5o5xqa02Mvr2E+69UhcZmtUL0SoLdsg8Bx8ntWXX2k4Y
b2hbrFWLe2u8VocKRilIOIh1nBEwE9wgVEhLqvQ8X/8ki9iI1QpEyvz8mvfLh37bS0jR4YL4Bqzx
TM6RJjhzrHGFyTDxj/GpR/sTmmBAqm/aRfHkUXePq9wK+sfGWf4WRfjP1WEbkZCj/UjCeSDmI2pG
nzGg18SlRLz9PiS/Zpv5N+OQr0SH1nXUc6fQEpSQ4VJwBr4Bw/3+DJ52sRbzKcZOkYQzQ2KZP4Ab
0hN6wBYkHAPr51UNcEDRy537QhpKrlbJDAj9tsa6uz0V7xDfOAl+dlv2sNvD4Inn+Vtckn701OO7
dU9cCUnJQe9exVVes0qxDq+FxgzkZlXSRAf05vOKBIYa1RrIrCYpoYIUXvi8IxfMsNICp50FBa0k
tEDvThZpIKJl4jz3Mte2qy9t2Rxblqgm2jcxnSz7ktLgHJ0C4sNLoj5UvKLJBBaMebe2Nl5Wt+6A
YpEm3jMzXYPZE9HBEyBlY1XvVJSWaWLLq8EKgRyKEIE1zPCmioCkK4cJqY6Q5zJoe/Lb2cUSiQJy
VIutNEZR8jyXiP3Tr8yXAEx9RdJIgepJOXK3SnGnTk/FSSgmy9pacKaw9AXBTTLWSy89D7BoUORS
VL+HaM0Y/C8juuMiwgdcoB4aLdrgtLKPa00xC0Msz1VB2QYdbEBJRJ0TP9syRkixrURPUvq0bRTj
htfEryTWOh74Eyj3j9j6ONsS03b+bObw3eZlUp3pvS7NOIC6u6vnt4xrgizk7HqT0r2QAg3MQq16
DhZe3H0vj7ONTGQOboNhwBPWhWGab2Ww8wesbsv7sbhRPQe2b4YY3muAvSy/xhjaEW6UgNXr9iVE
pKM8z45TgejlPdGJkPCoocmTISRv/1xmrZmobUzoU11TVhxXiWvXGmulfmbQ+rVdFSCM9lNGJOAO
FE/KektMh5PCiaxwoVVyXPXsGIXIvBJqTdyjuvl1R+3Ju10q5gzUS5asfH72a0ToqanTlJhgdj6T
3nXR/0c4a/xk1n89poIh2ysx9zuvm4/dCHYAS9gWAXboImjClPk4xNnIVzzR5YhZlHxMczSITyM5
gjNqZGoyBPSOqgvAmGENHLfQdTD0uZjusWRJXwD9WRqZhFw8tbtp4badDKOUplYfK019qlkyG5n8
C3rk3kxk9CP898bqV69fL/01S6Iz8bkaD1KBuh2b65NOimflM4L7HFZS3orX+6Wrl79bOMlLvL0p
iZLZCXLh77vSE85oJ5a9adPQeeeYheahwwzph834az0Qy0uMAsekL4ZREpwQORie0apLv4+4tFIO
UkElPB9RI/VlmPkRxb8rtRe0Hj0zaYCCElO4inDdSt/tfEy9ibjwFZ22UPE8MerJm5pDn+Ngcaed
phVamKnk3tPU+ZDZJfOfkTFgS0SDMWn3STcTktduMHPU7kHQgzDJa3XjRIkkTxWwMG+CNzGZBbiK
x4UC4Bc0B9vWHL9l7YYlwSXm+DVytUcwIhZG6JWZalL5Q93JHupkgoZFwjbL2T3mE84kEuKEC46G
xMLFlvUMjjJzoJunwZkR1vJqCDBkO6N9x1TYAxEshI0b/q2UNSWzJ5qBSIkW9+YJXYtH2qgP2wlC
hUdWR+gwvBdVZw8moOphPRZD4wVvFQh9I7xdjOThLrUJG1BwvbNYX5doiH2UuYaDYl3a90r6wAvJ
VWe30SMD+FAra8n89afl4igaFFfqlhACx6ynJAylCEC3O1TdCbjkIIfo3kBRftGvzcASQQPGBceb
N1aYnnN/AjcqGIvCul1rnVA7aIm0LsW6K3ukygxc61H+ihJVU4FB2ejVwApC012MqdUGFmFJN3wo
yzTL6cGwYXdJqlclIdEU3I6qSYTrfs2H0BqD3wiFr/9APDL1nt4XdgA5bYf4I2lNLS/ex9l0eXRS
Bd6KSUWiONq8b8sLuU2yVPlKWJ/SV0a3+wqOIjsP6NfONH4mySITEPbOwO7Tzipr9pNezFFFQUMm
TLVwK5OOgq3aF52qwkOLpEgBBnT4DQRjk0Cj4vyevV2REVX8QwoCoP3k1tDFzzt2c6o4uOM8v9mL
vMIUCPorJTrCFU+UHDWVxZDOowcFO7XXeRZdHSdCL4RGMGInirEnjnyi6flOupnXHrqKY2i2pFjR
zLlRunxMqMQRuXcMyFRZ8MCvQUpmQ/BMeE8PbgkrRIXQD/BlpFQtkDGkuNqCBNU7dQzRWgd1HIAR
4SXfzVnF0C/R52tIiWwacL8Jlz3JK2zFZngi+5YVHPMwwE7awmBw2FtJ8el5lMtA0HhA9hyOmD+q
5fzVvkvJ/E5YaH+A8Rh8HGhxrBnYiGIsr7hdSW6E1dKYVq+t45PXjnYXZf8bwG4yqmp84epF2KKT
SmJi7JZkU4i9/FFNNdZ+1R5U6QpYsDfNJYDo3Q6MVsV4kcfbM5res7R/5LQA6VEALSRh5JvqM0r3
/fUblaCm15T/T/syIP/zvdEo22r9tVxVK3kVPM43VZZ5yNDGvVQw/6fPJHXiE3HEaaHU+VovYUZB
kVofe7W7Py7fHZVnKtRlmJuZeDefKOYwui1EnXcqcjlahmkyoGMN8mJ2XuvJCSM2TDJ8XhY7t48n
BFK1uUq0qSgpZi8g5bx+7P+w5yyflqfXV3AZhyG8trwkHo56NhRp2sPCR8JdUO+S1undqTgwZeZz
XdYNgW9NuNhHij+WA3ZITdLRO0zZPekeUtfs0Juutj5TklaJqZK++uEpgxHgpnMR/tYuEHf6h7a2
GfpEmqngbbtz9j62IZmIGraUqgRBo3Pm148E+x5USx9635GRqRReqNdK8IaXOB9myNPlpitLgwrY
9OStraLdl03M+wpAbktQej2+fmiWgSFwXKHSPjmEXptChua7SOaKnNcqemiEr3qYov4AkKmHOBPP
mVTkXVSA+sIvx3OH+ybp+im4tFGePN8dxACqT6D11/INcVhpqM9nqgC/jpymhHNI7nhToZLGmpfH
fzPX7/z+ScFcGidLAnvsT42e0jzNq6LBMnkHgehQvEWB6+fMPY99wDa7FjhWFq54hoMAmwr9SV5f
VafoGK9xTzZjavLyS57np3szS9VvTRgwnsgJF0cuivGT24kHk15G/tc5gtgIFlibn1xZKumVa3af
D2eXjjg+p1nwEQFVMWXj/0gYqRYzyxZPmtdEr9hAyD9M685gYhDH9+QQhgeVxlhbfLVh+C7WJcL4
yFFgtOg4DQMVfa5HHdwclMnrinbGQLluFrkaY7R8t8aaJvX6Z8SBWO/BJZbdnvTEN3NmQM2GkEsN
OFEbLCMBK0pDXYZAhTYi23H+V2gLeU2RMFPFOfQvmirnuqJ8BS4JIm7VdrWE+FgJ1MYRSk1DAwFZ
dnwiGIkB3U4uWdEieX5Y4mmO8gACrfJTt6QEECWNc+WtnRkD9BuyP/Zy/aFJPjdTt69ucMQaDwJX
pnoAFvjWsIoWCBiczzhS0adHSHzsyGWSgOHm36y1dXkGkjWYE8eRnKQvh/4CH1OuT4wDbpLDsD0p
fZUvJQjFa9DAEEYT+6EdxSTv0feqiZbyNCBiRVVudgw+dCNTp50SCjkBj2iJ1xgIwHs7t6KjTOVo
N2b4Qb4R4l6oRvVNcXEMMfS+94mR07Paegbcnp1uswFpvtM2iEN10AnEIDjb32snI/Vb0Nn56lLU
jtMEj0Q2v3q7ZSOLlqNxdcsuuLiXfTMcWwaxn6k/NtN8R1tGzMrFsd/3lZv0bSuxrZBCGKtUQQ0g
jfhBkzlQJ9U4MsXonFILwIRyju0gE/aYEqA3H3GljL0QDzqV1aSIf6MWvt002qEkqMxI07ftI+7h
zfRLncPiKzQcWXQqsNjmD+rhrLZgk8CNqQu+bZlDLkykTy7/wk1Fav44y5PVrLdRA1Dm97YWiik9
R325VBkBopKhg9abWzsZiworDq2VHZ0Vd+eGxyBU3vpwPBf1yfIXaT8ZKRIrcChjtsFMG8gGlGMw
IrFSByAHFtGnujm2CY1W0XLal6Z8TPouomtCoDdIurP+bRq1q+VDDcttPRl3z0dAeItc73c1nGqN
JgZ7jkEzY4Nr+Mh+GZL7hUHFm4jxD5Esqwohwdo2Bp22ul7+j9i232Cgk7VdF29pzIeALFaioCeX
crJkHCza6enh9Y28sE6shS0Zdcp9anL2x//XAu38R2WdeJFSBoOrqTi8NwVdgIgcXq+eDPWQ2+QN
9k3Z2s1NVlh7a2B0f3//HOiV2/++g6CucuIoWg6yJhLDk52RNUAqgGcW6n6rQKAC1ziRPzJjbx07
O9iGHaOQQVAP9snut9hZyMQNwugiDvlU8PPM2CGcVlGNw4gc3oFRLjXX+t4S/r/KFm/KVZ1My9bw
A6lM58USJuVnFzA/7MelwZlsZURl0LcCca9D1rIdzYvv0NUfe8OrTPrS0Xjkr7KG926gkElPBpct
prI7sRg9SSlXBuHTn1tN1l5FoDwGRwM/B4vGz04m/UiuJOId7J47qMDDO7kf4tZ8Jf4EDA9k261B
Mq2eMOB+NXOdo8Bvs3Qnk3Roj0LA0/kxo//SQTByFbQvxUhYLYrVeK1rzxPyxsV++pJTUgY0bHh4
YasSLB4ovatQYR52bgmLggN9037v+uowyEg6mBZHdj7kdEovcjWqKczq35173vE2D3SLpnVPcNYq
2X0UBZtu5SvlPVpR5qvNK79HR/jRN7lokNgY+pPUsXZQAk+cmqdmoHtUdY2IA7i18mBMMFjIHt0y
KIpWGtAgh2TjbyvsMudarR2akYgcvSben8GuRfe13QXwcN1Fvu8A/4JA19X4NpFfR5Gzlj5l6sJJ
XSmyTptBpLAZ20+FbZaBwZ2h3nvBo7/6PFtdi2NKLqKIGHO301m7ENsAsYKFbhEJTz0Zk0B8qzdG
pMatmMm+5sNyoW5F2BszmLRMHTzWEmCkOiqCIilrw60QMKZdLdRWzhIFYCcCxj9F5CtAeFT8FgJH
gv4vNGegmK2U5ZNY+uj04qiJQLwHV5xBzmERGTbM8d9DIJPkL5hmz66/Z0/iD771z1jhDokYfPOb
deDDl5n6U91gyg2aYHU9WdKydoKYXOXrvahSNPlNuXafIqzkdYmTB3Zxq07bSoyXYrwHTd8NjmUU
ORqzVPwEPx0fHnuDAUZXxe0IvNBtQKNMrPrAvM05Kvr1iotykGbSe0P8sey4/HnTZiQeHVeMyxeU
L/vO6Ph5VCj2Jf/r1HQQ27KxWIcchNyav8ERs6IjXwTMLGxxxX0DaZMAHU8DMV3gLn31aoxZcRVv
VzwwTfCATifbmwI1zXSODerwZES1wVaICVojWrF3RKlOnrPQbtlTSXOrBqV57LXARlNEycc2SFIV
C11cp38CAb0NdpYY3/OoVHGL5c7JJduUyibj52RpLbeTE36/biCw2ld1ISFij+5u9wVwAYo7bNX1
z5oDzmBj9AhgecjIPBtX9xREIOSV/D5E4+b1W4/KcMoKDlopSBHbrmVvJSePZw3QVlzyp3gKN7r2
9jP6Su3jGnIxMwFF/JzH6PqTAU1SsdGst6gHbe/RIr2M+nhdN6r2i3batd9ZfWouc48jlu22CWug
TGR/YG7wwdsPoK1pyG/Zz4jHcT2vyYzMHuPwup4pVMXWryUCTXAos/mExjPAutDdT3187m8gYH5y
UxYGf4+wHkC4pRvkyBK6S/disl1Tr5JUrnnbdKq3gW4S897dMTJaC8/V6yXa9LSERty4+iIdJ9/D
sb0uPod0ZKC6FQGsUHHCiLduNREQleeGqmGr55NJMBWmgvapE99OUw3h/M0Qil8d8GNjOTK0VMWA
fRF+EGwes6ZFQwnDoJ4LAYoamcc1rccIwfVB5U0BXEaaIFIHFjBrjewRxm1vcrpeVf6+V0CBZMrv
P0RBEYPJK2/TsRnkq2ZXiQGZ5KBV0ZPoiRbBgRWcWsk7z92DDillIRZtiyxCSb3bnzjE4JflIc4q
3vtlZUt4tiqpH7HjiVV84z4CxGIzQgGIyH+C5Z6Nk5mj4+tb1fbes4CwilEWj141Ok+tAfgT1OLg
xUTHko5G7A9LXUduat32GxGBi5xQ78xfEHvCYs+WU/nxb7oL0BYyFbY80CRsWtFgZq6Nlm0hxlxW
5ErzPODRHpyc1JDhXRcCg7CwFLT2mCVoe/0Ksm3gOlJfle5Fr4DmlTk62Edd+dOEULRDI81MQe4U
oS+7TrdFUZzEvMifur/286HDyirUnl6Xd9qWrWJWOFlvSqzQmNcAMtJ0264TCGC3X+B+C93E7iAw
KBC8agjpbifwuhVOI2EgB7kh0TSe+lBLGIQpD5CYqFxPaWFahYDFgqPNL/XxY/YM/DHrgFkE0M9e
taMU/Dp/d5nkH/IgrFS5Ejaon1GIx8uXq+Tr/sWhPoyKVQcxxthn0A0xjPGPDAbwIB4lHc6WFZ9i
+s7GODb4+WYobWGnm0gqrg2tf6wGjVNt/AoHBBpDUpeOKx8i+Dxib/dTYlNWQ0y16XzeFkYU3X/z
ADGe38mBIMqMAV7AEFD3qnyB5yVS0piInHu2YLfgvnJd/4M/TVNMCQ6nVFaUFTLoFUyKVgxmTcqW
3IaAjhyGS3tj77OFOhxeib/2HRpsksFQHv6AoAlL8XyTchq1GxuYMFftmwQNyVEL9XXAuNi+OQg0
yMbdEA0W9i3VLEzeSP99674MJ6AyjGNw+kaIOfUtO9+Hv27KbV+eXt/xzQLfXLxvzpMukPwOvOSM
Ds59guHmvFZfVYM57//y92bn3fLl6quCv0LXC9PiHnYOlr8N1ZaEUxCbbuyCcp9Xbxl7M8xgV2Gv
rSuJwL1J2Mx17Oh6JwWhKhMbM2WQfDZQOovOwXBmzbAJQQRehdVsYcn76OIkrk0eshvBp6cpI9Bc
cz8kLz9BAIB52ZNhy99k+PWkK2Fscq1UwiWxrzOGHB0K2T524gKY03xMbqN88C0vd61bzJiFMsef
vS+k4ejCOBHrADGv0hkxlphXxeaDcZB0+kC4CTX9v2K0syGtx0+gymrdeIHx47wgX3KaWBk5BmXK
bTNAuy6AuQ/ouRGtbiARCBE8ARjy7IPc5BWLY1kSCmI75pUJ2XwDfRaH5q1ZSVapQIQkxZb1/i+L
LPddhJ205wNxde/Wa8B+Qyrxny8iNi/ASbVE5BUTjVqElYYBL+DPT39cfSkUZ6N3WSuKV8/bB/Xc
y6Cv1i6hcYde5hQk6X7685GeXctHgEKjAbQEpbzhOULaIksNXJn1gDa2OcMxLLqN7/5V+FIDJJkp
X4/UjUDoVuRopCUw9M1lTBtl1D6UWSQ4PkiOCn8uZWZpwcCelYKMH4wJbitT+X3bSGa9rZ4LvFLV
ShPZCgvbb7WIrTGzMIPfqIHQJLEVvBGfXo2VWF43Jq+8jzSej05QrUHk7okUdC7CDGAeJrRG3rYy
t0F5WsIntVZGckB70w+d01sfMEMydow97ARy564oR2MWDxS5o2jvNd6H8lR0sd05omGDmcZ4eDXX
3N45FtV+Z7pAavNaAl45AFrmybSPpZdcU81Xy9EgyznrUIv/zgD3OpooPwd8Pd/fFO5V1kDyaZiX
HXPZgF8HsjtGMECn26k2Lwgzc/Bq1FVkR46kuWozt4ROOKAjNw+tqvnsULShZoETHKQD8z/sOVur
/huvJTsn0Od0CWko01wbHewvuvFbI3lx/vjyBxn7IriFQKwX+rMy8FCEk5DLt55mUBqJxgaCZDQ/
Rk/tKSKfHoRSwzEi1EL8mXYZFQHGJ5vlCLxo0S2dkyPGY4t29shqH54yzOtccvYdpro3Z4KQ3K8j
o2uFmgk5Jo9IBuTPpi1eb4zI+0PFHGRyrcFClWxLPprK9YdhwXZ8MYrPyBXhHFC84MoE7xuixRxh
Mu8ivv7sbDYHs3ahr0GMHhXg+cpDRcCfe9y5Zq/HpTZlkNxfyGEV3hH5RVFo5pBehnJ9+VrU2Chg
wDkvoueebL+9VhsF+rIFKPr+PbKbgaDpp6tVFCqjHdci1UALtMlIr9MbLOx84Kd3V5GuzGcNJI7L
gCDHdXGMtuXj3lE2VAZPQsS86Ft8P6TbayNepIF7Vn9Tgzfd9XqQEhAZPn0KTZyUplgM5p4gP12R
r+vlqqg4bCBRjsZpaPpZ0fD9gkg1poVgeYw37E2bxUFE0xPKwhhE0wCAXneXemPesNxfzYSdxrkj
zT6JbK8UMuFY4BfbcBJSIUqP077TIxy6pnfXLG7Xajd3i9Dxaey+ELN0ocUCSYDwYBmeJRpLH68e
yNXHqIzKbq8wwoMg65lfy206gKSd1ZNywTjcK8UNwcBnnnUS3n7NI1O8Ifh52qdls0jNokSXjqrn
gi/mkfyAj6aTwkeZj1Pav63ZFz50sr+f1R7DRr1pM1Y7Y3hGT1xfbfnctJT8A9twJJ07dK6dcmvc
KlImfZbtjJU6+Djjd5wn8KmuY6kaLThHzASPHJc0seARui9bN6yJwHo5d2EClvMKadyFIthyGjnV
hAOvzyPvn/J/DrAFyKfROX9voiVC5T+hnhNN4S8SJlAP+HCdCDEVCb2d9xWZfOp20gpH1n59Hg4c
OdSZwj7oYszyfQfplIiEa3z7d9OzYs2FD9Oy248SUcsYQmeV2KCrL35gS9906rGKZjAy1f8Gal05
f2E+J/56L+uwG4ShtAORInu9jlPUtGJ4KZNGvkFRyO6LAB9ACeGjMtVf6Gkjkn8/T9CTQgBEJxPH
RrKytJSBji7eGVA2BJGQBlGXWTYd9nDovwMeHiBVhswMDSbyNv6UH3nFNmjeSidVXC9ANUuXNOTG
RkiOnQ6VMNd6e7n+XqhRS9MoFUe4e0U2NVQhDgwQwy3TTG5aWhfWD7QjttD5jVZ4EU2NaxuLteES
/IWoJ2DzmxJZDw+VWpXKHZ5N2DVaVhlNjrhIBp3DVtCiQxKqaijTbCBFNxLZPSWZTokg26Re/h+n
CSb4jKaTxBmeH3G2X0kytpqqUlkiovTi/KKLfU3dmhn9VM5NscjK5BqlnWYQiM6rvZ7CU89clEQZ
udL9QAPm6W8oTuIofjeeX24zzlCwsk7/6NoAASCh51oJ3LRLWJYewTAql+PCCgXI7Qq3BuBqB5BN
fnEHkmeLmViVexWgcUoUyIq6LVF5FG+IYBIIKQfx3CvmPimYhjwCPDUrvwBWtVBOGPKdT5Nw6Lp3
YVc1oCSI2Rx/kP3K1ss3ikJNncAs6I5V8yuz5PK+xb66UjlGG1Ehe0eb3ensvmaAs+OTMDscBDHf
jIbg6jjT7OPYKU+ddgPge60JBZzEQrJIGmXt1imAcS+1XUyBTzjiXuE2aTT6pCDEwQUHelel4lTh
05hL3DHEJWDbICi2/MFA1D7PG5jmxZAgak7Ot4Y5hpLFktKlGWPLGksDJSfIllS4th2tbOakZeUF
EUXMwMNILXXZ52+ZASAwOkGtlExOfmMLJnZDEgyboTRgRrDnPDBUS1jhzhKiW3HlLdq6MIzSA5/4
LBAcqC5RL2z0N6Z3cyeBPJSHBIGctNhQaAgt1zsb9rMhgAKgJuIQJil3hZ5o5S+eA6Iye78HEI9j
yMHSLMq+f/dUIfpVatGHK/IY3vFP87dP7bV+rPloK5VcJ8lIugkkciCcphBNo9U7ICbPSVGrSa81
GCEcvArugyRCtPIpFCnvuOphCq33Why+UD1rzDYjAop4zrNT/DErFryWXjMnIaFA1Z80WiTATBQm
8VDEiFAPFiZm6zuUyQAMj8t+biE49+NXi9krDdCjdsYvfqzhVmnXbKC7aqZcGps3tBcb6pZwpx9n
4FpsCJPrFXxzgXGZPCjHH8U4aK0nRqLNVMiDNtRmPT3HAoS8KWY2msqmhiPzxN8VOfxVF+V/VONn
AIAmHDxdm5EP+nol4J9jR3ooK22h2647W4U6m//P5qS2vYC+0GR+r/AjoKQevE3KwMirGahSeyF8
L+nlh+XUR+QQcGHL0ZO2kON+j/xl81LjUzx2+Bblq96DycNciv6cI9ckttI58qrzLCXlEPbNRoIn
Ltn2GqgldCr885xb/JVYmHMQtKdFVlZooAB8ywrGPNbmDO1YfHOK5z67pgyx6VBvbYK2lnN9XYII
eLWCeiAbkwWOqF7BrrQQP1XG//8o4RXpB1c0nWG0IwLCVf/ba6/VqTNUl7vjDmXnfDo0DV+PFsT4
72leuAX6+QPfA+wVQFAGe0rUIWVCn+CY0HZu8X8h6RG+kxW0iThpQKYy8q+FMjOWrwnLqwgGmkiH
pCyRi+gNKKOsawuxRN4GY/VysSsx6StgDrA8fS8KRmIdPicvINhLJtDX4q6gfBC0fLzbnrvdJ2CC
xyjgeyqdGRPUYtv9HLm3NpdTNSF0LIzoJfgRfcocQ49OKEnVU2pG/Xio7ZeDdhuPEd5an75gT0U6
Md0nAILlo2MipFLr621N1jPZqaqeFHQBFtPf+So3WAVC6CT6LKLNI2x35rzmIXF32OI0179NPTIB
+YY+dKAWqpBYT1vQgY2r4/jOG04k5WGGr+Ba8V+kMkCsKDjHTLNX+Np5j3W68HGqHl1QgugK5g7P
yu9fAYX5jKS9FvL62NGHP35FWEFcz/ZdzOeGwU/J9nX9xY9SlHIn8M7NgrIrd4RWj4vx/yImRZll
qmILqFhmxLNyELn0YTujLxGCiuJGu1AcbFPhr9mD6s7lMZS3z4X79AWTPvyd+B4IOvjnt+eVbSs4
uKkLbmaHVEv/4lBlyEnzEeb8hqF5Qk1l6NsCboe/UeO/MF9/d/yiA/PhV/Sm052SON6xNakjEY1a
cOfCf5/ItsjiZiTucYJ6RkPk/QRzfGzvrZ+3lC+fPqqsJz+QCx+O00Sb9NOoyZ+Kth35t+4R5yaC
eVFYJXWFbHdQj/HNFFy9yOR8cRSuVKjPziYMwKdeFRyJ6jHKNWsdCJx6inoHRGBSmxMC3zSM9ylZ
gii2wyfJpYr4BftNmG99kPe7ayRsUHoqSXBjomXe6oXSY9MTVs96BRAUMvspD4MOtmfJQ/OSfDOW
/Dm+JbGMkQnuosn6vd8tShavsjIgdTKQwQO0a7vdBUvp7KoowUkmXhRfQbyLeAQ40BcU7EbyMdGl
CKNVxxMf+IKaVxB1YkBCRWAQplpcOmvaASX8fhgkRQOl7KVyGvPeizIco3MDcu2bDKmwW50XKB3w
8t6rwfzUBntN/kfMNpQWGWTWvQpQnK9avYKY/SfjNhV9CF8MuFOz+ZGljG7MULptLrJKvK6F0hl6
AWp1hcOXQ/kF3/HpNzkcpCAq67pj9Qn/HzpRmk2Mqo8Hp8hEL51RLjlo5rGMoyv08G2oJDoChSW7
8ccmcXsEHIPHQwq/lGpB9EVi92hPp1evrX/5UhDH7DwPOwmDPRrFxcNp3S/Hd5YkNri4llbJUdkn
x+c63fbzs+1H0jZ1pluhlot0SmjZaRBB3dlUUnTtt+uNeh1fuugI3/KFzgmSIcYJv1T/4Bo+da+1
OEOfzyCsWXpz4KxUHyCT/cfjv4ZQoykxgxQ2ERfgp64t0P8Pmz9DcVQqsfrol/54C5GPa6ToboHO
/Ju3TdiV/ryhohGQ7T8CZ/DHpC2K7gGQtJVj0T7L4JYiBIQQRcMo7/pCi18MWcKk8lCn7kAF7DVe
BiKxAPqlF4DRP9dtjhas9pnrnfCybVHBw8lt0NgvBEXu53SyHbI6J7JVA86RkRF2lVWWrGotqfQV
MBxDaKAuh+yoe0ff/R28EQfCoBhEXz/wELAJmdukBrXWJXcgrBlgWwxDBpH8FhwbbTYYwvyhCVL8
xuCJTQGt4Z8sbKsaHNCapgqHIH58UOzVoNpGkeGwIpLs226/Qb9QUIp08DGXaqkAyUl7JZk5d11s
tM5DJtZl55sZieNs+5w+4pd6vRpGY44/n2pL1qQ9Tf5WWO3grggyrqqgIzFBguvRwONCxvOiKj4z
pt201Rs6eYV10msPF/ob6C+lS8QbrYqZ1fSxFta9RYtlUhYH2Bp9P+qol4MbSBhBJUatcKk95Pwg
3tFUO8Kzi5bN+r+YoDbzQhmKBrefpxRu5+XzcoaiAg+iD1XWBGjQqY1UAsHYUc0YSY7mrE5AYyyd
XXLuH28XUE391Q2svAew+wGeygkW6hvY0QnF0SoXocjcp4KAsLzwqh+fxImXhTjmKatJJRtjUidQ
gApUPp6De9hhdcxYrzvOpZvDN4IpWiP/0X0eYq5TnH9zQUVIXBbXpdzYzaxE2RU1i+MSPTIHdYej
ca59nM9t568RD8XzK32o3KfflBYMfi/Somctgp7txIGk2Kysakj78MwThPIXFz13doFFhoOqVqtY
+FeHLsYi54vtfgJ8i927kXpHPZMoFOG/agSocG68el8nLIv+5E6v7iNIAHPxnY1NFdzffuxCUE6B
d4VhgYfh4jECDQg+qmXYXegWdZjfvvZ8N19qVYZhWatUCWDkvFx7qlr525aobobW8PYRsYnkOyef
V2wuPckZCoNnW1lEY8vGqD6yLv1I1lah6ehZ+fx7hhmfkbqGhBnYJK0pAk5G514lvRS/+7pf/CI6
J/+51CVKKnV/GRsAEh/vxocjESjifY99GCKeAxZ2JqL0yXZNmaLpmQGRW8zBVlFrrzJKxEHGKTwO
fa5clhnhSeu5luqV9jr9EkZqyeF1zAMv4IcJSTeBnn0EMPqmdqzLkSGv9ofaenxsV51IE3Ykpk0Z
KVGAYMiPXEMJmXsIxoD9yVIRT9sOyF7bpI1ukTxkL8s9DZ5H6zk3O7vCsEbGpD2nO8mPA3pH8a79
2Up2w0oznotPKsz2LKOMaUynwFl6JRLNXFao+LWS1/UZlWE1PrMVCqUcUo8VxDdYVhQtUTHEJzOn
QKsbNsLddGWVVq5azlJLsFyMsskHq4DjXJGSlithDU+JHRQrTg0fINGDjo2vV5lWZXoMAt6kuOG1
pf/8RRGOUzSrN5a5HYCnlbVJOJIl49R7zoN3Sw5fvqekNfTdIkQ7+W1hWS5lKotc7Tz+eUR5uYdo
p1wrSngiYaAQQlbpBN/BbE0l7NfRK9c9XD467wWuK63M8jq0YcSGhvCw486rZYornsBCLdD17BTf
wYCDwMv2QzeIxybc1xtK2Z9N5pIeBg4aVI7D/TZRFWVd+eUwgSeXmofdxc/CZeWMm5/iEtvnNSjz
JpgybZ6OFyz7F2EzkDW382vQbXumA5L8l+7fKcPTX2u19zLRAYEGt8VCnok9Ldl7VUH4tiUxbFL3
QZjMOZ90/7vAGhuW0FajdlTe1sIiIqzrKlnl+uTEgSg43ReLMYyJhVwp8Vtfplzb4HZKmrZ2ksxR
GZU0Bnocg6tROkRcbshmrzAyfojo0fWvxjDSAWvYUVDNM+Zk6vaiOnfPvxu6H3WO8HlhKqGYHTAO
6vPDiRjxf4ofba9gRJavT+BAqOUudl7KjwFjckr88vn4em8kI1iAfFP4SRyISz6WRx8wR1cFq36g
1ouEaQK/DJ+gbVKnOhR5RACwAfLGtTtt9dkSJ0eqknENIR7JpaCTGz7S3gdT7xqXxZPQFQUZdqNI
kG0WJPKHvAlyoiRorqqNRZL3Oq5ZKkZ6ADG5s7xyBI6dyLgwzmZtsD+TeEmvwKDZqKOqWWHlwv38
RRcdJT+DX8a0Gv+9fRtRgaKl1LW71UjmpbmCZ1va7ahwOznphAaP2FG/uJza0CZ0/HGcMh9jYgv8
4IzbJYBoUrsROd/iJsrU+X4JsuZIvVEYC7szi+k1MwckRXY5tSbzl71jPEbLXyJV9iWWeQPv8f3d
YFXGxTOvch8FwBc/d9x6U0jbaTZu4lbIlpyt9oKKQh/TKZ9eEnXRph4SNIbWHXzz0tqBO7IiKDlh
DIgYPJw5pYYqeBckqmMmtXVa3A+/KDacUXa0PjuT5tUj7fFooj5uca+7cJkpweU+Tv0MyUBk9nt6
CYOZgBz29k7RlZsh4QCiVfap6IDQfRLfEvFCea228HKLgF1H5wJcqICxdzba/+LemlR2losjyfin
Or2Ssi/j6CxtADe5UAPyDVZvpqBM6oJlYLgnuUeqiUCCP5vOkAJhCn1YVZrFdsFzukqBAi2V4kfW
YBYzPNeFGlsm13h6sSm2b5+2FKnI2c8okAl+2IiQokp49D6PSbgnr1bLJ2Cqn4udLG9IAM4BCuNr
5hdaeQLJJOvo4KJh9h6bvXy/ET4GCPgJt28b9eBUp4otHBPUjj0QL6EA1bpkKPXNU+rQRKdxEiOj
S8RZts8jn0+KtL3FDUoCkpJYpd1NIxIkNwjozPvEHt7ilLUmcrf2OEkEbeFzGn1yupW+CfuDdT0f
juZkByovuzkpm9EPYx26HptIprag9DF43j3XrPr/ExRJ7Xsx5WDTlkBBhi2/Onea1i0dllnbIvl+
6Iy+S1PEqbCgtzTPe/saOm3udvrV9f2AOivpKic4K0LlrFwscENI9rV5ElWIjeV1Z1NCSBVVj/Ge
yfKtYqlEik8NadomAXx5E+8IQlTvpBUaVxElAH1epbmTetwfEp02MmM0wZXjNdQE0n4thLYyYl3D
iPYVXRW8wNyaepCgq7jXdwKWLMzqx7QngyRjyMWswzV3vzlSvC0w6NEKjY2cM7cMo117FBbpPl6M
qI3bauD5IAPIjMeH1uTKYLQ2xNaBWKC2ESChVpNznwp21uzJeJ4Lty3ProDMe+wuUfnv+gfS3xlA
Zmjw9UnUcahyc6huHtJ2DyFZsejldSjrIX+ltfoEKXTZHrvrV3O2X2fxjnwO8m2V9pYaaZwCs1IK
yoJ2sGYpgH2wExzekMTQvqQkg+GhqfNwZJzaSuv42LNg3K7d7OTwwn5IrhJ2+ejaGuZLYu4HKQow
EV49I5ybauY7Lw4HFPiNl4OTzxynr+3sccXv/iJ1DvgdUNQxH7b8GVxHj4OG9n1u4cdBcdILtXoz
0Lr2mtRCy8e2FqhsBtSqcSoeuHiCPvyajnAX6SRWB3PaUMGMo0vm3a2eWCSvLJuRKqAL4ZTNK3Dc
YCEwzZmrD3kJolOaseiOIbUDvca7OXLzcTIUIiYsh8xx0WUiBth5bems5L94nFIALV+/4KGeoxN2
GX2XCm8/1Gi8HN8kL3ud6gDcNrCnB0ZiMTWM7/UTAvOj7j3/IuqNoG6CUBPNcRYkecoVqdA1WdC1
jikzfjH53ofZPrGjpSAcv74Gc0fwlSNUExJVC8x0Ny5VGwxumTbH3UYxcIcS+0pjHwm4nDkAisSc
QQYg/OQOS/Hfxh6CCrGmViYXzcHFTmVxGqPnJNudAaPRvATVUfu4vcqIpXQ+GSETf2vDNJ1rteuj
X9uMtIfCa67tiM1MsbCFA7yYu2wqS4nqkgPQ5fyDkt1D5mBKCHVZYUJ4GWAClnkv4xQiXPou8NGj
dTsBowbloWfxkLkN1OCePVvw++OVTQmqLDME7wFZQAtU7IE36kMQI5chgzgv6IKeKfABEyX21Q7+
UDJ4/L4KOnlxx41dQHHREsjmBjAPcBq3UGbSgLnC1X+5xDum6UXLDOKl8vwHnWBrEqzOn7b7f7e9
ELAlUzbyVhHutd64zEtVonw2P12Vu2XGLcmW1XNMh41JCI1Ay8h+OSa1FE48L+kYhQV924+KnFkO
uW0ww85GKZMx8De9XNdrsTiNRWV75ojDyXOoLy+g6ZwQjTca++vm9gRPzZbfcpKL3drXK36QfxCj
P0QidiE2XIaR5gn/TKKy4Bch+sxPLmoya0qBOVlOAl5ZS0IUzrLJFGyak2Vm6JgSmMpPjZz8GB4J
/ikQRpnsO2MzWHUQA5niND4yoGxxi9DhnUJxRLczWGxt+j5R3JbXuxdP1wsj38Nt9JgEAPfl1MIw
NQt1gRi7Av+zaDg8XgdgDYynaJhqMTP1V/roj5iRna73xcNDFj0LdjEURB+nXwX+h97GF3X92Dc9
BywKYrAJ5dd99SdUbrtpBkaL7np0tZpy1Ygpe8Ozhl+JNUJhUlA2hXEQ1/nbtPsP7Pzdn+XHwXd3
ZNzkwx+6CAO9pTM4xrR0K+b0i0PFVcLDhyJjOk1EE9mHZYcX1GEl73r3GRDjnFLJac8O2IJuudHI
7J5s7aKwpSn1pvZHe+zLosagIwF7dpbb3vK9yw1IHvmDX0eMZR5gDoYix02z36rE1FqSd0suO6CI
xsyuGxexfCW4xnNJPl75D6xgxbyhcAs0OXcuOoqzsptHZGjfLF3MLPBWgYzyTA/8lvraivzCBPIP
CTywBuCUkqOw4IGoGixD8zAFitLE2gHKSk6/25x5mhktPOic4xDQTfCTTS9BLQSsOf4jk9LOfkU+
S+VphQ/Tr0JtAoblwYImV1WE6ZCHXBAXVzQSaSJw+Io+KeoZZyr8zfKAuiLOdXKYnmtIrh2pENtG
f8EHAF3eE0MjFZ+HOYOgu/q1GWitK64MCv72w6M6ZpfQAheui2ovTw/8J47hQSF1WyiOqxUmJgOW
Ym5B5yY26OUWu2j/aphvy0+eMQy3DqboJi7mroAnnriFglCQAPnrEiBS5pfw5egHKAtmFVR+VoFc
ZbN6XWkcUavIGTL2xuf0itUFeD+JHblgYWce6bD+nuQqcbO4BHRB0wbbq2wDvbts21E2840joyR1
QGDuAApkWGjZn/vedIN9TwJj+X0w00TlXz0Dia7DGH27psEiGCuY2WI7Gtt6
`protect end_protected
