`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CrZvMcRTbJzopeUzE3WHs8tg4BNq+nGqKVEgw+1mzTP4lUhlSY2Ml4y3RYecjxvxrhvVNAf2LD3W
21QqBm29nw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qh9j2FnmiDcGikf85N1LNuAPtWZt0ZyjxOdeDOjPiw7vy2U0Jt6g2rO3SZ0NONTncF3iI5rUSQfb
RG+Nf0I3cuLQZaJ15NX2Z4E6J/xNOJ4p56V/jYkliiBzwHBc1LhD8notAPU79WSfkKqPLsmNm1Lg
L6X7Gh/y53k3l/4WLkg=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zAVHAQ2uoHVEPlzwvTfzeTtSdaaD4hO73vuH7IdyX5/CYxbhjGg3Tn74s/jpE2p/rQD9ql7/B3aL
7rtbEaffgTq7ZCcJ0KQdTGRjo26X43w9ROYS2VQLaJhylEXo1V52L3ZQKEPKkcWD/XfmH32wO6k9
Yf0Fg70SAFqRIVyI618=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o8waKvjSvUZO4WFJkdTFo5kxX4lE7JEF6KZiZMNrZ/xkYd7RfJL9hoh9Cr7f1cMyh9Q3nV+EiTxq
ZocVFY4ocZb/5y+Cu8mOZ2I0Qo05n1Av1xltfhUlBCcGQhOrUSr+f/dgJiIi2bKe9/nH8MnSGqxz
NQW8ZtExrMqis5LnJKLpF4/lA01EhfLr/GSxZLXJzVGL6Qtp56Iq0L08ujpjE1y9hpbuYszA/ndo
+0Oc3yYExS1k6L2HfslZgjNLV6elFhsiQFYJ09BHN3cn7oKnI/5ZLhw79zxM3KDg/KBLmCar6Zut
DkC0Py/KQ5erIamb+oHzogeqZHCIHHaLUhLFzQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y4E8tJYFBYgPuvbDhfHOsy5OJa7kQfC0S7yhoVks96NUr7dm62HYVq7efZxDQUEGs4fk3fLRS903
jk8ba9RVIcj7KreaI3fLTl8R2JGJE8sZcdWHcdsK/6LRwL5eQSrMr+wTzaJUONYGJ1a5EBpKuaG5
zj3gk0wFeD10Lu50YUMVwek53worQfbj5o8AIiwNiwAcbLIU5vXCAD2kTpauw8nyS35K3MP2MjDu
DU+q145Fb9915x0mg65y/ov2ra77ZWVvCLQtnKZ+jZ9fmMjLfC+g11QJ0m5yum7Q7hswaou44VYI
IBxIeIqJ3nfB3s74i3Lzp016Yz2AIS3fi8k71g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hI9SQF0K6RI0kLdSmHIzoNiZMcgcDVxDdkwelw2NQT9EtCHZ7SH8TDU/R7UOtaEL5lVQdgTfa+y2
0ONsLdQ02iWylryr9MKv2/+rSlzfTQrFETuzGNKh0CNs+YgYdOYEbqWBxm+hnSKyLJJSVEG745fY
Y32Qt9TssWLU4zqFciXf4T8O/BAj6TbxIYeWNuyuXPcoe5I8yAb236ayfN2FO2v8s6otpx/a7pie
yXBxuuOUXx08q+AzSSZlIkVvBIxRNgwTe3qhHeekm1YxRKl37TirZlKdCUev7JBWU3TaExPOUoDa
wAMU8Ysmqv/zIZ+01v0rrXZ7+8iUBV1EMCatVw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
QnidroiFtHGNE6OOr0EuMkyZzrnGZ0/50LYOwegQT/CfKnuIRc9X/wbqp22GpqqM+kAeaZDb39l3
QRuBFQYcCZe/YbM6Vwfls0Y2smzRlxDzCOUKe6jq/IE+nGPv5Ac6z2sojb5gChNUzEtGB/LQQFn8
i+reripZh5UQlKPdZlr3viaatI9mhHZoKpJFd3hfg+/eUI/Shc+DRDM/ggrSfPjpjY31pR04Pcp6
UiJ+QpCzKpqSoe47YNrrKO9oyUxPuBEukL5fVN6ebQp2tl/5uDbj/fvrq0RiwFifgpkS5VVvURst
99OSPddjqTYIll0hr2Gsg79/H1/D3K/yXAllCnSTYCa0LvU4uOCVKzQoZoaHxwvL4zyL6UmnXss3
MoEe00REQk2uU5nE2rQeX3bthPSFfGIj6311IER10mRJi6Oym/5E4EFGYBiza4lPkG/ZUd9F/IBJ
T1yJhicbcpUDx3vplj/FHHKE7MKL5OOf1el14pMddscVyYSo2bKntB6hfHJsdUATVXjd8sfFHt88
v1QkF+WG7N/1f3UtRwKVcGeRjukyV89GDb7Ho1UHrQ8+e3UxlGM90XWUQuxR64SaAbCLeTTAyztp
JGVOFFujLCSq33c1R+p7LxtWOki8F0l4NY44xqboXhdj5Toc9l7+x/laQofV+eIr9tEVAQbKWJIa
k/2P9qtXn2ddv/EXXdkwhPyfzK9oF8t4mILoaIoAwxNJhvCjXA8JJKID8gVcKZ2OqPnONFuAFabf
FCIHYWoXceRBe/l7MoTN2vAYJTrptsvSvnK3qrMyc+FSOH2ZEKo5pXHoe3XY4gZbfH0vVN+6GPCQ
QMRIhOle5+Or3jyLPCLs4/1WXNvOUM+n9m778gs10OioK2r/gEycRitWWjMsrdkxWUmi/QGSPKmo
WAdIjGmtwSU1yPjHzIKBqedDU6IsveTyvBa4IIQ2LTbxmkA5F79vbap7BJZVQzfFGyewZUa+cvne
dLqm1kEDw0NnhkV6uAgH7iLP1w7fuR0UfczWiHocjWwQOJo6txe3KPJrzsKNLMW2fIPkF9CfwStR
fgGaIfc0sz7NHcVXil0z7uE8n/QV9TrAh2D68W2Hyzi+wCG8xwPZqb9pdBkUdY7n6+c7l1hhIdgE
Vxnn3D78XTeLy8uhe61L1/5NLdHp9vAK2RQrgjjRt/DUw69DwNR2Cem653P32mvbpUi0LrVSyDvJ
rtS6DiHTBwRkE5vV0J90XE2R+bWoa/ppWkq6yrfFBLsaQ3nSCt197o/YjBFl03k9lYUj0jzH+QDk
Pdvy/knbilgCprr/ku3uN94CC8vLRogsbhJsmCPaikTa7X25vz/KgAMyV2E0BKrQHcmyY9mONMjG
OctgR23grwLPItAOa5mmbMGGuqvwf62293vnjC1TeuMppM395GuQduWwfC+6p/W00o5WX+u/BhsW
CJ8+cCaRg2hGL4/wXDFhzHTIjvyp75qYNA+m1vuZ8/fXFNE52/jdATfZErkOtw03WmYDHyj26YU5
yfdLndwTtnmQLUlGOM64EopolkNuSwbWSRKdQ1mmBwvgqTGnvZ6UTtZJqSYfH6k5kMt427S4ehJY
Zqlyd+AzHH/5K0jElVU4mqJNvAGfV+tL2g6J+AZiTL5ECxHaPcsT+z3r7lofGQFVKxXoUe3YXvfw
y8B+5BlBA6QtTeNMoxYPwuFsygk7yHCuSRO0cEG2q3sJzY9falItI+ZXCUrukSoZAN09d6K3DTtY
xamDOmt4oz/NDH5tkZAVTtvbhAXTrvPunBNlF1xhyInLBj9jzupE1RHVl3rW7ArOEo/kxmtE2qRg
KjtGoZ28YbFuUZUrivF/1OP5HZTlwWGYhJki9tVsHh6foJ9tPmaDpIFAJhklj0c9zqmalDOif4gm
Tm4fMSAPUoEspxQ7uGAHgK5rMjvZpVArvQinRC/8fHHkgwK7RRkJlIsiXCB0pRnAXJyeELUKkfvt
kLEo5rily5aq1oV+SZpjNa+Ly5qau5viNuSjL6bouFPD3jCzoU6Ays6XIkra6vPQL7COgd7H6j4X
f1Ej2+WfLkpRc9y7AjRqEobZ4XRzYX2F957+cxvBeokZi2MTiNuvE3DiqIRA2IYEGRRkvE3rf+B4
piTe4XvOgcdbdtu3zr+C9zMkPsXbbGFGGVTm8qO4CgRuAzpafLO331gSXGWnqSNdkRraHe7HtgEy
ebaACgh3bKRgj6hOdnHDSg4GY5GW1eEIqSVCrXQCJ8CGDJo0dqEO8tdMueODZT+lrHkkMr59hdYn
9d8MjkHver7Yr2m/tXlloNoz8mUQlXBix8Lf/DteGdCo9KgfcxEwUloPfhRZQG8tYqUNCc5Fmhm9
nkKlSaYLhPEfdd7stKtDo4QVRliWTFLK+emCmQBG6JXs92GC9WM56nu/8/MHfuLdXy8ze5V7uHhd
vsplUfSk+YkgLOdQpWRybegYmJoWlAaIJxdh8mkRZWdkkevOQ+slE/bMmvMxZ0jE2a0YtCNdetZP
kj4EunZdDrCqYJOCl+Av+4swxvReWwXu/58AMuNjDUurbJeEPTN9rLt2vqwRfWRB3Fi2CcESQL+T
Aj4x54JgyBDojUwjFki2p9lWjWvJvb5fBZq4k0SVYz7hQRfdaxQKWwxtPryKt1GdAok2pmMK+OHM
XFcIEz0OMYtDvr1M94822t7Hf1vgCGhgLkgbuKxnR51MiXE0M3AynHoEoVm08cp6jiICgXTxJ9/O
9pZSVGqka2FrnXPTbj7/l0oZX70h/tx6BA8XiQ2K2ZsIK0MB+iw4uqxo7LhSz0MM1OzrM24nFFt3
57IuCSkFlJlrasxcPWeZUmQM8qKtiXQbzglZy3YWczRFeYXveCRTafZYhWTO4EvQjsT1Krkn2NvQ
PGIDyqPXDpKXRO4jvEQGT/RkEXsnl10sC9kap0ff0DeLgRF4iXwqfUneIL5XOKT8VKloYqUSl+0T
wtF4xD39zPCOQffBpkS5ArElvtdDn73AvUOeMSg+mWzslapEJS57jicz0D/ocHtE4WHUEPDkdx/M
z1XgHeNO00hoXtWX468eeIeixx9DtHewwL96O781yBizynFydqV3jM4DN4y/T/OG5FJ803kBWYPJ
naOZjd6TyVbxPI0pfoVV51h2Sd7sbfVO7hmUyg5zzLRvifpn+WP01d/vdk20kDDx5ro3vLN4i0KU
2UZ9h9pLDXhPMPu49TLspN3SDmtk6/XpbsyWBhYs1k3zfJL4BBR6G3YuIr4zQ4lWzBZnq3Awpvtw
J5Skou8MKKg8V9wTmf4nQ+3tWgLnrrIyLECA8bYfSUGLpCB6P+Atx5aYy0PmvGofCjozAbQjzSlM
CtVKBzeU4SxpJwZPOBhJS6TXi4o0boXjQZswhSYTlILBlpeafEegG02LklZdhaJcc1wrfL8zMv7Z
y61RONiIIKvAwkftQS6YTvjghiyk1BcpXTUctQ95dfJo/6byaTScZclb7nM31pcWPhirX99thfEN
t3pAmAQx7lUGyfTo7DMyu/lxg3qbtccyBoDlzhKckCJFHwo3mxQDTQ/Z90snvNbBdYWkB3XsZMoe
SFcepp4kr3HCDF5jh4r0UAJ5OCDnrZAlXTYW92PjPf1SKsSoPrtQcwZ5QO9z/rCze0WKtEV6NY5h
4KZ8XZ5LKPDf3MQEKsV8OXKQFMZP7x4obkp4hQs04woGvYrCFMw7poQYI3ajnrF1munSe6JDUMzx
WSu7Y2tzcbSVzWgIwE66PsvpmvejEKfK3sq7NYsNePI4YXstPAx1xOtHzsxFycRQ8GXiyUadZPUm
oaVDAhX+D0Y58aBRUtDfpa177T/TbQVKazRwZlH5OfwPbo/ZbqkQqc2uqv9w83uJE9GuXVXU6fkm
eZY2i/Omh+D47aRHkh+SBohmXm9hpL7SQV4Bgxlqt22TwGqzp52PChjNQ5ujYBekivS0HG2f9ST6
x8PF+YiAdeoNzaNrhkTszKQ+TGK6jBwfO0UbjxDKTwvascmGckbw8N5SCjswQ9NYUrPPp+5Twa+I
IbhFGspiK7pBsTiPxMM6FP7KheAq9nQUJ+r1QmNTgsv+rzGSVlgNVMOcvOUp/xbd4SGF/v1jCZuD
ow5tXZYpbA7jAdvI8V8bZNgR4T5QYadrCZhJxEnfFzQWa/Yo+ZjqzScYiWsOGhZcci0UvjvjmmRf
1j6CbVpSn2LZ31BZfm8gDG4/xmAd/DsJirVccbQeJzuDYrpSD+ZKHDLE+N5ZF6YvpHkk/4PV/D35
JUOlOtMO6PtqN8p0w0kovdVER78Qm4EhrtJSCh6y+QnGoelJrjkSpLsrIhkCXGLb5JbwdLJ5M/p7
XrlzKHR41laUGwBT8WVjQ42wNpMTfZ90Pdocy8sG5Q9h2Tm//24rqG/8Mn5KcgXO04dt1zg/TMCp
838eiOLkjQe+eivjDm37RmCEa1M35tDip0DchK5s7tmqpLvj8mAdrmoDstQo/+EgMsY+EoWnr92q
udmKIqLRhdZO/I44TVLBsSKZuWvNMrOm40C0hvKmrIyf0gBinLZXtC0YVnUGc/o+LamOwGdBqKeW
Y3WtkgwcleQmcOBmJQMZgf/g3PIGbUs+5+d1G0EbWC5zr5P1+q+O2XWmfKn5zsheyLLHOd0JA1fw
z4cBDbdb8JZXlc7aafp/jVWA1KztM2eAhz/8s2VtT88HjIPttaQtL7b8x1QS/1B07/poPJxT13Ll
cNukkrXu+jkN36gbiVTgNKcm9pR2CB1Tzm5UL0wPNX4CNdLs+vRjDYaGPq8sqjNhX0cMP3r8Qmeo
a3JANTCK1SVjIJ62GhwxIflBjZpyyBt3LUBu/tKzO8O0qyALUsj42BT5YXYhrkxzzadkylf0TUFW
GdirCVUYQuHHr4lb/nHQrOz7AbuTyHMGyhgUX2vsr0UN8liivN1JgrlEcIocE4ZPbAYO/9PQ8ae1
D3Z8JYTU37EO6yX/ShJBcoY1De0f0nI0nLilULMz3zDL3Lg9m88fVwFgf80Oe4wXBNaeO/87mjax
cy2G4rNi59xBxSOs9sMVg7n9cF4GZ+SXdV76PG4E9OBd+lYytvTjO/O3e+PG5npKpX/3Z676DZiZ
Rj2KXIIYiampgaRgFBrmWylGbfJTfVVcbSf7S1Et9Y+NZGuOvX11vxFifkQC4/V7IgPjipQzhbSH
FP92v0pSoUr18qND+mAw8EUBcwHpouRRFF1Xk8VzzNU2A4PByGQyWYnTm8bvLb/FX+wyBII3MJ1p
w9/7j0rys8OaWJ9a2ffETrOxydoP2FP0gY0Nj+pMZZo8SCTEQbsSRT32OPPE+O5GT+79wphVdpI8
/KB+hAcG5Dit0zq6qsKvWXoeX8gI6q/7DD7nXUp/aWFY+Yk472psA1luGTTrq8HuReFAfa0rOM+k
ZeCdG88lrvpBBPM3BEPydKl20piA/Pm8OtP/Y3Hig2HvsQ6zQ75ak7QrXnDjSWW2yJdAXcx9WTqm
DWBQ1lGmiWuBvuZKJmy/QmJG3IxT1UpZrtwnMCrffGXe+vPhBuLJB1U82h6S8vZ9drFMznQ1DZ/j
FHHnedeaX+9RpddGuHGo86o57qxjchw+xy9QW3DUgceBUMinnO3DkIsXTr/TawexVSKYXR0Kg6/G
uPKjQDi/82SYcPx7xhXs2GYiAU2RiFFDIzu1/iI268rNTnsiWbZ/IOS5TuewF0z8tGC1m94P+N5A
KIySWjP6idwGK7N43IhhK1KeD2ikxcpGhRtBI4EXB5+RxaFLTuNLbxz2TxHGFKrVRDn2v3oN/nni
FNYkP5hBmLWDSghAwAER4m4UyxnzmVtdXhB41c/PpZYhcNodWPGUGWbjMIMVYr9M+kHL7nHxt3lV
9VkxhfH4gqRucOsCYl4YROHN1fg6Dg0YfWjYV6jSveHEggAYh1ETxV1+XaPr928QIq4n/RkWq4y+
x5H5ecIMEG57SqIu8g/MipP+0G8i/pqNZSmKfpHPtN7j+869gZKWjsjIVOeDl+f8yQ26MYmqY0ki
9h9MWg8cvYAKNRFTJ1QPsehmLqQNyYq2Y3aNJcghgPSBlQwlUz1Cajt9dE0HcYXdW3SrjjxMo0eO
PUjtxxog1vOUBCr0PnjLEcKoF3GvUHOPcmfGSgaZ5lTPEEdH7A27lLetSCMRlhcGLB/vHXc/uz3x
NxzgNoeZW8jjeTFCHSxQqhDq+jNQUKPIDtjIyOdsDQM6sQd0EaIcaSt8Ncx/iUumgEe04bR5XRoG
xGgQrZTnMl3e5mCHaLvvJxzJ3myA3m7lX3UmlSblyHlqEzHKNal1b85u1JNIVGu+U3LLrRkYEPhk
dDYu/AepzPJhny7AnvSnJLFpYnV0Cs4yJMBPL8WDhUNwVgZDstF0PILOCN7+aw4p1g9D+P/BHwJa
N6T4yeYt3Napfh1YffOsiQ3zC9P4nUBWP5Xlygh1ww7e/WFb3qyoHO3N1vIEDdSFydATDYtvl6H9
2M9C22/VDxKjKPucAPpLCB6hV5DZL9jBPk5gz0JLDidSk2M8dfBKpeazsmXII3phMfjOK0HYl+gt
2/K5tP7tHeQRi1YILJrByaZ+EAQaoTvqso4SVIBvbJ9deD4/RXw/WbOs0qL1RstaO6hBONoBFbJm
1KBw6vMsDbQlMHCx7d0mawVZRECovxozKuhD1unST1IG3jLuUD8hysVhDrUCNWSl4Dpq7GahDqc7
Bf/7MqSv2G2uXQPvDEIF44WTNcAq6tsqI5szhvJRjjgPAl0q4330GUAD1b0xOqnfpDHd//uFDlQg
fzlA4w+6eAHhT0+p+ocDaSxkoahrdpJEPoVN24shXuUKIwCkEd+n1tqHm9mL6ZWjpzzARPe9aBLV
XusSnZ9Z78rU7Uuf0bWQaQuDnLNEJ9cD7NNXjc40iIm50SZXosCq33N7uihGuEQ+AgalWl+iIzAo
vGpbLTPZdqWZTmCBfni1uG+bHfRt7adkE83EzwxkfblQzBeNVEXLg8Plzbuv9pULW9YSRHwg1W3w
t72hONT2ff1G7X5tJKbGXKavIOjuPZHYtHftt68HnYxDXSiMAULAzkqTzDWZVntW0EL5D7kXmEx8
2YKMngjVQb1sTZ1my1afYdPlGF9aQz7atuhqs8SpEtYi5jnY5WGIyTngVJmR7f3m8wpY7qUwB+Ht
aE88O80Mbey43hCe4+Ii9UDEhalX5jO2n6RzANxfuCzcTiSowN+pb3YfCVW2391YAMXgr1rnGPty
Bz4mpHIeu6bPLCKrTLNpd4jdSQfnwQN+IOFKgHxgtEeEg9ur7fntLPcf98aytQZO/X8ah9MtrQ1o
pEsRT2Hzga7NZLUmYXtbGAQtaX2Ptnj4AJV2laFMhJmYm15gr+qrnfOdC5lPw4bq+x9UUARxau89
NFH2lo6LIvDD/61aGDQEGQeSFa19ZMKqUU0YyjtHu+uLSFIr59uC84bVMTZkd8BZo8fWeDSM/5tB
dJWLC0gaYLndXldY0VL8jy1MeuxxZ0OYXdaRlHd3Tcdj+/2SqUMELaclpBByZnJZHrBZ+yBZ7Wuo
uaMOzMmyAbkvq+BcBZMWQ4pjWg41IUVOSQVYp5Z3mLW7Jn5vFgPekJP/8AIqxX3PcJYYBwQPffAu
Y10f0rGe2Kp98FfdN4iw/1Pl5BCyasTQ4t0PCOfdOgNqTcbLAdc+Fse+XBc5rGBVp0Yb+xBkrbeN
OAjpgIfsHsWQir15JQrx00Wk0OXEU8mn4UEZKrgOBJYAWmsu6p7nzbUSj0TmOAM4kFDTbCCstMl8
uqHCfQYDr4XoUZim0UjckyQf+KgGrT9QsQoKfpuUkTRv9nhWLAT3CpZxzoItGzJPApu66EleJ+Hy
DflGvnDLU33DQPqzJuYW+kilbPVSZU1vZ9TvX1oNUtMIf99P5QeikysQpqMXdtcAtPu/PbNs52LS
ZwndCTAGheSEHH6DMEBrs3H3eoHlon5fTpiSOFsxNgn9t1oJNP9H7Ff/jpsQCcAwF862Ml0Emre5
+HxEBTtDwCAJlL5XOx8uz4BFAdsyt9oTTytUQJNlNpvc7rE4kIORAAC4gflH4vD6D85S+IxkKCq9
Lhj4WAjAibP2DR2cPosP3oeKQqb/fYcVCTKKRue8XAKkzLVTOQXLkrJOKlrm7XUgRUhCIj8DU6jI
OkBWy6qm4LXx1AYm0xK/pOaKkWFFymak89g2IKuG5rQETXYOyEqhdSDvDXKiXzyNwp0tAdOO9kSU
jgWW8ELI0K03KFiRWZVVTqpyd5FlpWgdKwQcjz9B4vdiCD8sAJ1Cmo22ADGDoPlalQn4XKoPwHla
cZDAA81gZo5vggZJetdwYLS8z/s6cKan8IwNmMnO3D74z9Pv70XeehJIfXcyzFD5hl7r7b7qXORL
x6LhcZdH3FrvW+xHmkSvAfOyXtWo+esZv+nek0qaW7BvEuMGBKcDHyZTkhoaKiDoILHIll89i6CZ
/rVyMgh3qQQUnCpWhTgNjd9oA4nRzQ/xuReV2N2Br8H++AqQqE/8tdbg8oggFgyWB+PKLHHeHrJi
MMcW/DwLyC16vPt42Cj/855wJWK9SvgUPR3ovd9jzUR7y+0fyXxReRDaGO8HU7lNbkYhVat8on57
lnjvXk5wuwQorg+0blu4p5lsBWDIzU1a2/A6OyojA6wZ0xdbOlSz5B4GWeEiK3R99BsHLtb1iXuB
UnM79Yvw9qgvsiwj0hAWVPYhIkAIod9MvnP9TT62Z7XVcXyjrrp8Wc7XjMne90rvaV+aT3Tt/yKN
EZUPSLYXu9AGGHB/z6NrqkiPDCqPNrNgPRrHiql2ZnDbLef1h633Euk1HrrG4/orFAMD9cm04g8Z
VA5Gs4rRe1TvgEQyebv2jQ2amX6J+jxFUAMrQ/2hJpO3qe4Txh17RgZqFhr3o8YNyQ2MRWH9rMkW
QRsXiVAfBmP4aWgbM7Zxjt810tpgtxo+cBDGHukILr2lCAOXdqkSWKHVH6B6FHfIaVJKs5/LJ9uj
tfbJpEOcQ786s+1eFYmzfgX/38P0GARiuAmPyObrKzaVno+HqP4338nT2DfZ6DoLkvq41UTKodDc
KPsCExlccFRQECIA4RE0adG66tXk+QQGHjU5mnu3yXXRdpwso/yLdtz2kiRH+H2M7vokmui9gElK
NDdHjNOY56bSVIkGDC/Wg64LJDojANAMn7Yz3WMogZNt22LdGY0DTAuswKsqAYQBv+BukbMRH4qf
YhWt0FfUD96xDwC/3Un5PTAeahd8mo/9Z+ZaTNk+JsCCBogHfAnS6Z+MxADBhgtsId+akKWxG9oR
ZpzdWgvyygklKr/VZmB1KXQu1iedKXTet3QFIbJtoWMcY/Ljw/J8bzMYZn+2Xbk7QtqyC+sGytfM
O2n9x7Wcfk00GAFsMgPaWcln4gZOiDCK6DyAHMSJW0Cl+6oTPs5iIWB+YetKNfiXXQTN/NYxS6/0
e8rgQrt7QMmIUZz9Gm50Tb1vKNGAMg8IQBEdowg7PiBUc1O5LQGGiRvCzivgcnDNjqCp0O7rZlC7
b0v89Th+1bFeiZ2Ip9NkvT1LeOxKbHzaBFPg8sudS8H87gJQStci9LkIgfrLm8XZn9MTDi+MU4KI
Gs9z8nHeDdSVVRa1CwVyTm3dqrFnWbxn4VNOXll7C0r8KTPiB9u4Lx9ashCOo2c5+4Cc3ipvT8LL
gCk9pUrgWkWK+e3GFC9Hwc3Z3uu6EwFkQnKxal0rfLq3Z1Rs5LYspE8WZWvgEy4vUb2sD54ZI0qX
sxTtQfdn2Xym5hDcsMyG5Bvh9qniumi1jty9c+8xWMoazq5PUvQ4UPRdt9NcuR47Vjw4BExQGpe+
EjIx582IkMiUl/c/qNQrx4WGnMPrSIhXYmFtlos3fyTMMBsbk7Hs36rknAx5GIMgpLj/DAvyj6Ii
s9v0liznDW55LVQ6z9BdAidZBXZAZNSbwAoHkVBit0Qnw6c00MH8dBnY2IkyKsirQzgW7QGqeoLB
rLVxGjpyKbi0stjS2R86nG++aMet03aEvrure6BaNOBvG8xImwwZB3J/BIQWyEOSo4EnZh7UwmZf
H6UpnTaPEcb0MSQDIphuhOPS2lc+GG7qMklJ1eWlu5+R1u3Wt965dkFHq3EHpeJhlguGbTN++DRz
71NDcnsJy+VkeVLXsp57CQhxB6P2wcX8dqHjSXagCfjLAvCaQUAYb6jiTHUv0w80LF5ioi5O9msI
U/Njk62Ynxl+tv2wXNC9wAxfoc96rM8xYEEwIX/xRno1dZUKr4w/ZI1J6TowTNmR/iiRCBtTSLOi
aPFhy12/htq65uS30kl5z0K+0sm6Wy+0/8avx/bjq+TsN4HmzmTVrYqRkdM7Y0uVRPLO7YoIu3kR
9By8kmmu6u4S7rMsgp8zGvDrXvoL/cmYZuXO2PVHR6vnrG5/Idz3tlJ37SDrvo8Uq0P15kMBRZiN
WgLX1f/vhjX80nO/gnBhANRtUpk1eGpI4aebOggiswhIoiLSvF5Vq3DpnymPK282wLcqZhTZy8cP
Do3M0U7VZsfSReT/FNOdWxxh/Q+lFsHHhcSKHSjNeycKsPUjCZvgTbPF8FbD5usobBHZ5S4N2VFN
3kCdUjR1C67vVPSCrCqqvl35H6+Nl6jU5TSQRS48nj0Ky+YcEnOYmI0SdDo2pNVqySoN/FghI2HZ
FBa/qtuXBziMqqiYYgYSp4kkewpg5omeTCbFXwiwul3wJ4ICaARbtk6zVIAqW/TqB3VLHd16NZgu
Rxif4t9KKuOlEKlusovDiBmEyvstDHCt+HCYBWFxfLsJ9wznf8mRnnBH7ba0pVnNHlpBr4OcySep
MKx+n8aGAqyx8UqgbtM+xYaV6IOIKh1QV3ETEozr8tE56A4BA77DMTptdfz0mc5a6LQm7b+2yh1c
qRMYrt822pHomvl7H/uoi9sBiC/qv6SXotpnZZltTKz7z3ROAMCfcCyfpTdmahMSAw4sdjVfBy7L
Z0GQCBtymqo9axNTMceEwK8WabhhrtwIQJdK6UhbSbCwBEJkm7MCNappKdzvxkSh4ESZZt30FLtk
aNsCDMHpP+Nf6OTutYM1X5a/xDnebNoAqc3g0/uzu9b/3RAuMsiRY9m+Vpi2NVdK36//8Uc47gTY
nE4/BO5OVrs3UatFrhgG+E/TKW/qTz2siED4SkB1LL15bCJutso70ecRPEEu19rLzAraHxgKVmHz
s2AvJTdNUfAvn5g1VMydgIZXg0FjuIk1eKfOxZsi2eVItdeQBU4uSOliou/wzhqwPCv+jwFdubV6
qcct/ARIiQu1dX/kr1+pwUZiKPWkydn/7/YNKP9GxVpPJU8NcuoJjDaNlEcucvkuNdxoPs7e8Rzc
5XknBeje4SqMuE6Wu2KE92MLwrzqdgi8aa7aJB4Ab9+fHcftnHhTwlMzGWMcjX9AaIY7hTRie7Gz
rG5HcuG58LwmyBe/bv7KSmOxk80KUbQl7fyenCPcrCTn2VaL9bRunl/18ywYiDGz4zETmFr1Hd6W
2fRspxIwUiNLizx5KWD5hLEBdmQqeYVw3emBVUBihdI51LA0m6QvymhM28Tkdc2KxyR9ldDYyWMB
jQSWXEvMkAtEkzR35rUeM7VB8WbkAdJl2rLh+MqHKIY1HbGou9d9IAeKqbN+e8WQuZYWbuWwpG1V
EZ1VhSjzHygQ1Wva48bTAhdbST020F1vJFfjRNTrVi+O3+PYaJOTXEhXi2gcXN5NDbc2NolQWos+
IubLI4p2QXgUGEPPq0AzJNgdb9JU0iftOdw3hL4WTt838T/XakAdPhVBb8zMZ6oH5k2lGR1OA726
LkvoJhKufPRL7I3LoA8/g3TkVEAFclBgQg6NN3naAjhamm9m4SUtWoX+aQR25hbXpJa7jeyejuLx
fWEZztQcLDYJWnzZIOlgkuGkbgHyTsCqHQf3sn9R8UnGcDnXMpRnUxlLB1h1k2tzKXu5CZoZ387b
Tm6/ujrlWXvcsouKN3yMLCSTZVGVivDxfrbncdjOVgxELqje1ej9l79yi1rAWfgsC/9gQ8Q+n18U
lroPJg/3xriP00E9vvEdSQ1lCnOhaF4ej+GVogYMdipQhU/BIotUmvu52nxoZ0GGoS7dl97jp3uL
aldqYSR33RAuTLdysi95YTWrOq7exUMVLbre46WKFzXZCI0kelthb9I2/Er+3bepDg9WYhq51Wfn
baGSSwywxoW5AF9//nlHGc7W7IOVujlmq7JcUVyhH9nuawDVH4zuqt3ktFGK4fnuXtOq9K2C1Q+O
uq9sPd3/GqQxj0pIhOViO50avGTt2yzYLET60YDFF4jtSbfeppbNn85oMTUUV27AoB3oklEWVGZ+
IYxPfo9ShyLFDUtFGi4jj4/qKVOLVuumAF7ffVIxX+33vG5YiZ+PRvw/iseECMzE5cDz0DGAw2fS
2ahiYxgmLer6at+TPTJuJ4voVcYkQXopyrb92iG6Qu8+AE3GhqS0DQ7nnguxDzVkA4pANDuKYDYe
r27A+XPTAU23yq836KY9rbfvNp98GMHvtfl10TPS3/QTO/zw8qrHkwve+u3eb3iL2LXJKHU2tzT8
g3ZzXPIG78hQamSMhBsRZr6oU7UpRh0qfbXzGvlH5Aod386onP0AdsfV8zxUaPfAbYsYHnGnNiCJ
+yAlegpZqVthk/YztKcXGKxv786K3YZU3oJmiDOxHIZrFlxrWQFitkM0uifyGXc8PAkKyBDOJD6D
/OK8qwzFLKQymUFFgwkhqfk6QDDZoPr6euhxi/El/KGwWsRJxLhRvXmPcMYI/s8dMcwkE2kybCir
oLFORn1goVwUMbMaW4W2dHQ5eemK/yK0xSJNJLdXP6x1jOZaKRZ+bjbSTxycEvpZai3wlSW3xw3h
cWLrYsMSaDTQtQ8HhEwxICZ+wpKgxI/iwddPrw6QAqLc7yUFI74d4DQL1CG7ZnvXNtMsUEK3UPMR
zmaxHYVpFKD7NTZOOcguH1luq1zYp9yLe5v/sz3+GtONXz8rVSeG75uqERg8lfDT578/RCvCQ2Cq
zrJwfJ41vaZKJEblJE3ql7PL90Rpop3deaOmvqTsCA563FsBr7J6+YF9aLJo2Esw10KsqOnra7pW
Ui8o3YOXb0S3/3SxSk2EtAONiamKFR/uXsglHdwfCba3EojTF+dbepoIxjFK6e8LdnJoghTD3l2C
p9lNnjNTLUpDuq0QZ17BI/+LHZO7/tsecRak30D5Dvy98m6W9alIWSH4XhoSrGTyVClB0Z5s9qhy
dg/rdky0WwtHAJtAkHWrxSxuTaee9VcxEJX7ShAKh/n6HQsILKRFJotTYSdmHVYzXFNlPg2OoXBf
lersG6aIIW386VSsJ4DEbWVsAO9ah7hdHe6GgGfwB5eN02HLvXNa4+o8MYTj7nc7SffZ1R70CGw1
y+R4TzFiwcJIDL34fwj+XExD5NPfkNXjCJ7muwu2hhf4cTOaQWS8Mg9yetKOvQ44G2AZhR7/+nzG
vtmjaUARpiZsUvcwPAQ4+dnfm+6AwrFectrO0efYrmyRpZ9kAwEbPenIYQfLEYsAyL2fFqofpEFO
fkAMh6CCJ3d4+FHqgF3WIWE2WacCWzIwghUCcAsRPppfXfp0ULeHUGdsO/f1x5c5i39+xoN5Wr2h
NNN462oYl8BLV016WdyDiT6tYPje5UZEOY7Ym5SzCgk4xFzFbjIR7J9MXpANwm3fqXGKAhqaohQp
SY6UahHT53J0DRGMFCdEDB+yA0D4+o7yprzF+Z/RkHjrTNY7xAs1J/uFaMbI+oSlBKj3Y+USTusB
TaWAVHqQJ3SOUtCSHJlpuOUS3XYxIYGMwcDhkPwzjk11m7H/4KkQlr4OrIW7NE5hYw4aBVnL0Wkw
lawgKOYriEMP4LxY0kVq6QGQibtc9YTXQOqP32dwaFtwrgnxcj+qETqGFVvAAqwDZHoWPqVQtM3F
4WJNJyb8Ai/I4lY82EVeD/vaPWouBgCgsHp9PYHwN19YGGSXcw+gxC5ghJLMdQXZwaXEAyJwisNJ
mxRkRKf8rvz7W+QNOZnrQsWpPho8r0CjUqSHUrgIUBSCd8QuWecr1i+0damHPZvaujS2OjoL4W2z
WyhvKPKuWc3dActgx0smLx1Qa9Wfsk4q2nqFmcP0qSwY8bMzMrTWhd4t4VZKS+2Dyu1jrh5fZ6GZ
vRZuvVB/PQVI/VX54820dK3X4wKJMrUfPBZX8vPxvQaiHyThj1mhvc7rQWxHWQUmp/Q/u64v6/ih
5a4CQlyEfd89ihTEOtCIVSQHfFSUvSnGdTcaG4FkbP69gR+Lk2xlnZcVRf7kBARYEQ+n9XzETpiv
DZiEUivkeFhW/8sfnWUMJrGOGFDrYwCjSKKbaLDqGxEEe22bQwrmTBZ0/NR+fXiQ5or3DBmkmRXF
bT0Vza3EH4ubFcoZNWAZIrMgr7L4R8hFVV8pOlT5VPEtl6Gsso1AtDmQJU5rMeFpz7Dq4vupWMWS
zBFw3TtrZP3kJ+I4qKzDk1D+b6HbIdkV2jnfW680oIO7ZcxLXnJzb0ZFM7Qh2BgNXaX9U4jsBeaw
QCbCOv62iTNYV/6v1OmOtHyIxXixEhCFa8ao+OcxBAiHMTc1+HI3A/R5M1dWR1tbtAdsBStMVaUB
JGOMPqr/ZKA9JlxW7a067Kt3EmOaMNtjFUEW8RViaUeME/7Od2MxJdgTlM+juUbjfV7xQb9U2IUN
82j3reduVoap4jNe1hGzYOS2VUJGdaUG4qqNuntSslC8FjxUcWnKjE3qXqe7ieSrsZrMCRasudp9
vRHalu8e/3Hqf6GxtSrd2mZJZ03ytYTKemYz+uXXKLRNSYxbUBdJH7TFHqiDJphCclPseTFih0vV
asdUfYkMsybqH90KDYDAgj9x4HhL5cVKe9TvtDX17/11PfSxs6V6LFUaTdS7aysCiGXhAAZaMC2Z
wy83hsyQO1vodcq47R8lYHW/toFgNqbdf/mSIHwdFQ19A4bN9Pi+s0PkwsGylcKo8jSpSdLUH0Vj
G8m5jh1sUsBXAjG1GBlRbxRkzfMHTA9LELGjPbhezOFP2BtIW84tfGUqjdX3zH9N5BBfVB6VhR4X
IbnTsN+D/wvRTDfwfnv+GSZPqLfCAeutqRKLHxNXOqAvp65FQvKQkOF745Ax3zz7vqssSFcVM3vt
c0QSC2ZZ+4nMFgYW/11Crbtu39I+SuUBYbecizTprizeX/f7cCb8u5YRVjGsRaex2Y8bm29tY9aT
FtUycxQanGu2ZfqeduhTP1XZ4mRRarAe0XN5AF6ISd7/UGYJmxFUeREUwopS9zzqjxH5ZZu2Be29
dIP+87hPI1kLAcdWI4rujpERS5zYFwiOr/YxkYIw4UrW1KTTFy9REOI+T31+fr847PQ4xnWdZUPc
9QVyJPTuI9iKXjLc+ox1R3bRL8arQHJN9RzbQQBYxx6+Ol11q3Izl8rsRj2pcfYNsfNVrSJYYArO
yI7l5RMP/tyQJygTSpXKXo+5hIjplp0MCbeLT4ty+Gbkpxkn1UWVmiXpNVGwI2VbpHZ+GfWuyhiS
eTtt0T6XeQCZ2eF+FVsKDSY3zWcjsuqQi8/Qdzsxzki6I1LKPA8qyPp8lo20Ly9jNxGyEj9O3uA8
DLSw4vDWwpRgSfezMsiVSYDX1XSGR8DdK5ttA6mHrAOD06Mo/M6+eKgcaBUe9DD32aSONy0BNY5m
fGdJ3TbIKlpzS7YQFEDqF2GH/LBJJclaipOSpz8NpevKqPFcI+B9mnytzXJvt7XXOXGiDm2NGx8X
bKq/IPsQpNPk4zUnrBKuEhhYtKUQmT72Imb99lbi07if2g6OGfgmWHPuy9Gt7SCyVaHWmwFUyxYE
cKvQ96oYkbVVu5jD8HX+cIo9mp3ii/FBhJBrS6nCFKSR/cEdfRXg0mW3CmLOtzwq5u3JytcCLN0R
V4MUTsBjQXjd92gWR4Pawcwtih2sOowTlPQwnTjUk6S8UEWc7nqBMwcSKeGcNLkRWQvgWHpRm9xf
b+81tdoecRlIFxqC8MGvzkTS/fe7IvaXo3UBLg+pI0FtQSxjbkC0vgl0f4tZ4tQ9/Ki2PJULx9PO
JxF4jhNk94pAwKSJkBA0umDPOdgcb9uXAUC7rGXx4BJ34dCG6axA1IopZ3+DRTSGH/JecWS32rhF
MdMrW9BszbdlaHN4zt/tIv8LpXHAXjZNNS1iOANA1uOu0zz5rUAx6RPP4lWnSt2QROQtCCbU34J8
ZDo//IKJIyTTgkVBshoUJQuLWs/ljP9t8hs1RNGv1oewP7XCqDUbc7dqY8GGj+9q88Fj79E8rgEo
+fNb0cIRORWq1n0YF/lYoifiWZmSPr5zmRud+0xqYgHD6Yn3Zx4z1tK4+xH3S2AlgnGljYOcpo89
txOYED1dqFLhRVthC13PHsVsi2OAssoz/cXmdwZijpzkNtQDg34BaGSZPNY4vVA1DQHODAS5cByJ
W5IqTbTyM4kK82mpbEuG0lLNwlEzvGNN3PWsiIE6uquslL/njtU35DSsLjouLoNqz6afwqt2NzHt
5jPwQ11U9h3LxNiLyxoXfz/KIsXN+Wcb7oMnxQK8YohWjHU7GxQvfYqNrhG/9AflIkT1IqjHYbTY
+ZvvxJCuwVOe4q2YhhMw4TqPGxCRpcjL65ecWjh2OqOMT/e35lLjCjmvR1JLnmo8YCHymnNlBIdk
vPCW5P3rs5cb3+K2clt8pXGKRU0q3ZUoXBTQJtwK5HPaOCGvm00BzxSMl16TYX0nhB7/HnUgAUFy
FrNk7wyBWoRzbMgVjy8gi05J8dQZd3qB6Ct/GUAWCIREAKwT1Cqvu7Y1n24AV411G36KlNesW22V
TpXozm55MHOgDly6hTck01sbDcHFkLdBA88+kj0c+XATcQPGhKv+ZwPKeSv0EuUXv+2/0xynXd1k
yz9h522qSl1XNWRnCce/FIpSokTz/BAarOuOBXSaVnAaUc/9AjrQKvHn06B5Db5WST+MHkCDQ7Q7
mu6iVNMkGVz4hbe4HO0AudwGKwJgOZNgSv4vur/AoRbbXW0nj9nRI9ogGnXe43VJ9uzn12ChueKo
pMhASTs87ehY6T/5YGZfnIiqn/6BoCwyhHZbHXyHr9B0iluYGVun9BSmhA7HGfO2yLfUgrrzuyBz
cgZ4+CI1gIU6sZ03BCzm/joxUDSioTkXX0jshkuol9nK2sqaPzcyBxFb7octo3t71kLkGbJwC87E
KAqsmB+jYuCJciH7qo3wCP/RuZljZ6Q9EMVbIgASbb7ukCOtL5zrdVuKfcFjLPfgufPuqeVoxaE5
W3W0Nuem1UmD11VB+K13RVAYMLGTpKx/YQL5G3aje6wz/9Eu0H6uOpx7HKNe9TN9auC6wHtWUyt1
sNfDYmyYM4p8ityduU14q8ebJvo5L62dWIvjovpSkX5DZBh9MH5716F4bJM6qgkwImI9wiDch8wO
vwFiFvRDKUqn99fS2mKUR8x9JSI/zADFGntmO9rvr71TqV3+/YbZiVOME6jIMz85sV56cnN3nchq
gv9JmQnF8Mte/QAKq9ouR6n9PCZDggXmvVxp4O2e+mEvIfITemoy1ZJh0S8jgKeWOCOqXsmtmEc5
pSyQ3K+ENCkuk2lGklMeNn33KTc/H888AgnVmdoil9eLXzCZdNOOiKFRuB8v7weYRzRorGwRpXvt
wj1aMojCrFsDqtYjzqyr0FZW1864AX/bRnHxZeItxuWQDilXNF1F3thv/WrfIH4EjtHLOnI7qe6M
d6Z1Y1lz3SoJiTGvdMUtSkgdldtUaxGj38hq+2JQX8dgT1V5r89X1JrIY+iRQuqybC8zN4VQvThT
UPSfjo2DZMa5zrgx9rxSus8KQZKJ60ylxTEs1b0tZ7YLKhxskP7NDq+lyzKaAWytP6HMv5UCEja9
fOkWxCgz3P37G2vdjc8yWHoHXwec6me7dmqgHrU3XldaUsx77qLgVB2ZSpcbdONIo+dZVabMMLce
B2tQTqGNPGN3QCihXV3Po7hRGh483/RQaNfWXEFqC6XuosnZ54pa7kHLft2hwI4uTjaber5kTkvj
4NM7XOR7u07j/ZR3oEECfi8y6ANRe4mnt8qZG4zGJwdgn2+Zt1lsoITF+Ihcrj9RYHKruCrAUmz7
793fbkFUgnZN+mP2+oEEPHJYkVJ/gvG3WTjh/++7AmidJiOnWx/rfirafs5maut8w7L0MqIEcWSb
aMI5kPfV6s81k0oFkOvoFrkwoKB8+TORDKLhq+51fJmeZYDY6VyVp/bzWrUe34Mu1ATwlq71AX7e
Q8KkDxA1iBbOIge/tlbNu8nrmBtyDy28JRcEPTC3K889Q08ikkf81EW3g5rcrp0TulbYADDx70c5
Uuh8vnUOyuHdZyi0/YshrgMvVaFLyAVgAWSbuNlTxPA9Db0OtcoO5kxAWx3trxHigrjmKt1OrJ/d
otABlS8HP9vmU4foVct2z9bIKF197VWxksgnh6hXC89Y9//8WVl+0LzPiCsVaYjg+rez+25uTSQF
biNELbSTODktP5KteET41PVHG0/UJ0Q9Nc3Glt7cFoHQV4bQoMW2oJEV2TAeWfkRyt2ONmXuWALw
4V6OKAw5LDwvK5lFV21QynD1gUYqEiDU6nB22jSIe3+/6br1vLLHXtUWWuT5dEsow5S0L3IUUl2d
SfBK9gW+ECV3Md7XgX7ThgvmU2QSzuonnRV/osWIiXx+FmDNmZZPod3PDb8FdTvubmJVsIT4tsGW
3S5uup3mhhiqDSKj2pTubIOcwHagA6ouAgg/NdK3FDJEAbovaC4ExIBzrUusZXSDQhdy/pRbfxUm
C6CLGdchuCQJh/XuGo506P73KwSXCYnamZozVlAN+FTdu2LP/qRBVoZqOAajrxNfhEnVXuLI5Ybt
AIX5fg48K/BN3KPn2E1XTNtd+Yunj7/QXhjovOeNRlBxTs2mWN8zqeYAe02MRpJqcrrsdNRDfqGR
zC6+lUUYmYnvmLu3cyRXNwg+2F7Bii7l+N4c8c3Odz5YzHdKcMQU88SXvxvKyGBrKk9VKr71UN6G
4925uCSoib6uom8iGbP/UjuGybn19/K++/TjpOQKJonUDqYcpfoDy2UNAPCvTybWE4aj3oq2gU9l
4pd/np2mO7qMhjY5/LO4nNDFMwi9ChS1xTg1+5erczEIj467KBvWyTI/UH5EMGUe2tUyPXg3zaPv
qylqY3XVL6SgTeFy/TlqTgHXSGtG0B9OvREYs/EVHBaWeylVQFAGwG5HX5OYuKPIwN7TV/kSuWcL
dikjieGR8bYURKS7VTmW58kz/JSKT69yu515oL/7f1RPuAz32TiuTtZ+fUI1iHp35fdybjU4ik46
9/fBc94w5jBe7KyRwmHODO2BSJ2lReHC7IFEos0ccCjPj7QpxXSMzn+Sg66fIlM3QMLJxlgmSZmf
jiZWTzia5udABa5ICibJ2iiYERnykIFSpeH40qoatWFP9z1yO+undEDpZbT9W8GCnnv4/ztNM/Be
ivZKbBX8ldW+Z6R11+sBNbUHz3rcWihHyUUIpfZXRgfZVypdjICs+fU9geVqBd47esICnCOXypZb
D6ybRReFQmzPSJRGlvFjQn7CXpFnXdMdpeN2N6tJGkwWonsyKNBkgG/6XGmCtTqvFh2/dfwLU34J
9CH+aRN43WTnCPT7CvnDsCO84+najMbDa216EcgtlHHxMOFDWitPgWFCTXqwyrHpuulbUFUp3ipp
pwyPhmpyFLctPETzWi+4bhzi/N5oDuvYiYe/QwaYufMamd3JCyrSJYGxKPVl26OolBi76AdUokcO
nv7FgozwU4Dc3z2XY4C6r4wJqI4zh+BtWTgJ29yAOVzKiF07brC4+7qGKsjwa1OUZP1RIkh7+1Ew
V12yLbkfHEECBpOcDVgnT1Rh8jpv6X/mSoAbzclpYZX2Y9BuUcz0hKgz8CE+BomiA1Vl9NUf3bGP
e/IEXHJlpU3dYXtaYmKWsHuGUsjEvSLGK0PNm84DdVi0RiCjrtj1ksiQzlLrIxLpUzlVHfOxbBt6
riXW+JcMcFCJpVs9WcMaQuyaCb4UCIpj9KODMlIUGf7eEduGMvnutBKyxpkUG8dWU0gmbhBySGGf
S/tIDlHS0M8NJT2ZOofIATVMSgBCysk+SWtEvDzc7t01pPrjGJLNvdfwUsRvr77uedDlaDaj7FTz
O3oTujwar+wtHjreSFGiyEc3RpABKM8nkK+KZsMDOyQk+fv7FHMvnnT3NkbLvtz9THeAEZiVEyf4
Ok2I46UmfKoWKsbi6WORfKokgJbTbruy9d6eIvEGvgc33wg/4Ivs66T/cl++O/qA4PRNQzKo8dm5
3/Q0PYpDj3VRmVQ9XSdyroV9LCGVhpuPRBoaGZzsrLTuWbHkDiHj0yURZoh29iCu6JI38H6HoBK0
QaSdG4LjpY6ObuqpgKDru2i2X0t8ovA98N8rsxZl1J/l6jyYYpZ8yD5CyZf4C3twytQE/lZLlUjq
9KNXOVtRpUPTuk99UN5wUkwEWTIsBnAtevVpUfc8PrxVnkwDem9DRCd6ybTd1rc0r+LofqadTzcX
kIra5s8SKyVW0KgzlH7n3kNU/G+B+P7BoJt1daI8rAzDcy7ZTN3zTtrb7pM1JpvZLoaP+iUBdf95
1L3nEdw65+JROnzCQTaLWlYSXucxDQhSzIT499PHQFi8+uXwdMa2fNtIwtp0HWKyb45zOEAQFEyA
mqUwQXLBouZorUr17cqj7iFu3I4zTwoZ/KJq6ec5uWX33FCS/JBe5u+iP+FaBgW5ahcc/457R1oJ
yQ/pG/lXZLOFU4YPDQZ5e6klEP+4f045xrBDwdxOvaMJytfT8xNo3Hk5WxxfNP/v4Xe+tlXJHAxn
SaW3Ed961f4JaXAhZGUkVToDb+JHJSImkWpTv5IawNWLa5d6kFHmSQdtsCRm+Kk4+SCqUEAHfggx
V97gvwElGpTudpsmrYZnJi95V9qRh44/eEx9mdrey9CdzTPLxzX0G4lBOUQoaXSPu+TAz9nvHU4S
JUJ4nhcy9hLulu11ZxsvSRmqqFELFTYHU0fwWWvBBaEQs8b7rVYT0dgdm8OmXy6pGxExOAaTAGXY
EhYx04vHsCO0R5+jxJHZTpSwTqY53NMjtznLKUFxh8UhoirGkLSfnskpi2cKlmcnckZxXar8eVwG
TFW17VRUkPurx15SWuIGpTqig4sBzhHoD/7yAzLb53y2e09vM5NcpVpteaN+CZsAG+dZ3x+AMIGa
SoRO9JfASu1+ZCY9UlcHlWcTQTHGQv8ORhegt1OSIiHytm/nJ1ruG0ewtgxqnAe+zf4n2ohIvIS1
C/YiwF0pEv8XaS3tA1tK2zVcIlpoFJEJJNWaxAyL98IdrbjrPTUyKjN/HNa3zNNAroWqR8GjPecU
26wRCHqjWF7+35gNf1WoBgfcLMhHs2CYwxiR0nZp4RwqQ7F1WDykLTo0YanaPCLzEC5sT7DDFl2H
95tmL1S8K1GzaBTmw/MLKTZbtP72UiaPiJ0j507OJJRjzsRVokBx0yKMeFt5L1yQNF6eMtquz83i
AdnyCmTLEPwtswOIaeiRvJdmDROdOYCTrTU/GbLhr7Cx2OSXF6wbtvqZ6QkNomTvJuc++NnJJm6p
x8Tv3QhuH1fEbzxeJTXr85i+pnw4KIy/aZwKb1I48mRdXgD9P4dib0eQR3f9Nm3EYsOM1gmC/fiZ
1cPbYqH/oFS4I2MI97baWyHVMXnxNL1ZGcs7pxcOL2LKlFPgI/fnWZLhofj2dn51BSISIgWCCtwf
ijr5noIzTpqcjv2+ZVp9DxWc7Pp/VNAr+dolP5XxrCeMdWZCbOYkmhBQi4T3/v0/vxdb6UrABpkm
/ecGDMZYnPSnfP2YSxE6t58XH87tjqK3++NTcc8YY+OfZzCcHzUOHiaIscO0Km0rMdT3TmuR+dmE
0kcL3I6YLigNpFn4BeraDgGjYJEQOwz+0rP0B6vyQw8OeKx4MR1u88V7BwHuPJ0ILf19l1E5V0P7
CQxed5v55cnOIUVyiTbYyqodD3qqn0YHW13V9kzChd7U43wetJeAtEwq2eJrOKOLSNao8I2a7792
JLQfbMcN+4ATw8WWBR337f6Fx6iS7IJOR809AObquH8MChOX6LX/SnR8sl2NL32kZcnVhwLsmHwL
peQUiX76ZK8/oS22DBpoizc7InNdodtCd9neLuiXWc1cl4QSruejoNsruKDyqMbdU2E79vvjUi+Z
z7zLTxSSvlDHOfcaaCwoP5LGk6k/Zlr0aAT98KVIi22Pt1mCrIaFX1Zxd69pwMwBhokrI0CDnVnM
EYo13hW8EeANxUQJsuZdLylEl69o1Kxh9z+8EGD9Xi7lmn0dDCsBr7PQ/sD3Mwj1gEndNJTJ7ewF
Rge1s6k8BxYG7Zd25crdb3TTbxH+b/WLXdqrsYoc6LhVTIcWA+5I+gga7PTzYqGsPWDPKFbYutzC
w+MnYKrZ9y+puR9HTdo97H1URbmBgH+8KDHFhq15xGNU+6OK9Ab5HPliHWY7NOLtdmrxtrCGk6y+
n3bRRpJKOXiMABnfOUg52uIBHHGw0zM+WFxXfR5FAxaBm7OBpSpHY7CjVO85HBQjXVYvOlEtgVuO
PpRd/50F7vm8YtZ8u1JTz+rrBPPgnSurLw55SwH1EzO9epwKi3zlLmkLxyO7B0CR3/IkOlAQ0MPP
rPwzsOu++VZcE3SmUsmmVyoRbQeh27SlwROTmqGNNb3WXWzs7bOoWWIgO5mMt2Au1FVUG34vxdmp
QlrD/um4QAfcSdYyhwU6ZkigbQemFMgm5wyUu8tfXZWGY8JyA5AWtywKAujqpwxBM3Imn68xYOxw
JLKINJiiU4urASfEXDSDMIGUwIY1Sukb1rUF8Zv8HurcGSFAJ1/IAwQfiMEsdaTot0NBPcVGLIdv
sta56WJiHpRngfZh5pi4Z9kEMSDUPVHbG4iWzLg88T3wl1jPNM2t3uBtot41ALxWXWvzwa0kY0bk
oQ4m9Ae/olzWnRJ4J8wvmWP0wKsjIPZKmQfPsV30zpgbnV36Mj9jtbGICsKIwoeM8EXbIEtNKgrm
HmHsMKkPm8iES2shuQUVdNmPwEdryVNMmZ7RWw59vQymegBaGOxGUT+XbQQ0nyiWFTL7i3HAMWZu
zu6sZenIME4pv/DBgQXz6rAqur+AMltdWwiB9f9olMxgYfqKiL/EnW9wtjr1urXaah7hGvvH+kZs
5o062YoXWj63+Y1iIwyNNomDydr+GPUsMBS0lydpOMfE2u7HVRTOpwzETAYaRSlZ+RX8eIcXizPF
ufmrkaIS72Qfwu7IUCIDpqmP2lFE7STM3eMXDzzgI+eSyOP0molgdEqGA6pKz0w0xoVuc7zj0yoX
LhFb/SOyQog61OSCwW9HIAy1IV90c8YNtW1hnRwMxFYykT8ozVYuwKsYVKYXJ284xrV6SDPKNB4p
JBmkxvGlOc7K/2ftjTPG4ziCyI/he1MtYkTeqBln+AsB0f8fCazY/RX7u/1ah+ikgAK4WoCM706c
GcsZjP84lXcGnJ2OYcMlDWc0a2KWAyAeFbDMjk/7Ektx3w3y8GSRsQjplbojWeGg+ov4pJScFokx
VPvhc41jmCiCQ3O/jh8VEtWadCa0JpgpZSmERQxIW7r6qD7ErBAOSvZL37T7h/3KJq+9d8gxMMpc
k3SPDbxVVs2i49NR7UATlqZdO908KtLtCBG2X+Ce7TRIjh3CL3E6OFalvivjKdpK6RGJk/zhN7g4
0KQzcmj7U1xYMJORGnYkOOY2V0csDp3ZV0BbLDF7byg8i5jfCQ7owwZ41cMkbgl/4iaBUbhkkhBW
k0CTghAxU0JhMeDzNPAyBlAB5jMzNUnC/sOx28haiC/73WCtE0LgWn6R4YOtS6vhZEfNIUiYWFdI
C+Bt14n5bRoC+hW9jh5/eeqft507HntiKG/6sorgQlBVfS4kv3Wr/yfLqcxjf+mznja93wcFyx0n
fS88pwtP3ZsbiYa+NB7cc6dxauJsTIHr+QJYNQa1X/ujwnFPsZop2Mnn/NBtJBe8egBZXiHO6J8h
ox19emr5iE07lD8nYcw+TIQJ2/XZV6MCoAqV5sJkOmIjN8C5Kdlg2dGgmhzf9atxvPtqW8uL1Tco
ESaJiv/+77pCYGagAeE521n43LAZ+CNjmkSt8ck4kzasUFrTUVsu5UWpJMR4bzwgNm7rQdL4MGSs
2PdHF9yuja+QnVANhcjHfVnaZ+97QsIMBMk7nagPjsP3UYU8k2xjW0IvpkZMd5QGRcWlE9cFjtZk
xRSGHBqCjKSo4n47bFfWlwQHZgvt6MSTxqF/1w6C1HlvbtePyzwlDScXhq9A2OakEXYvIkG586mo
MHLQ7Ft0bXn6J3eTn9vW7Cezc3BIPJUgkWqSmaq6Ar+jnsQwV/6XGnqUzWGUA6lwxYT8LSpK5y2x
gATawoJngwfa0y65B5pZOtFheaKBgM1L8ctk1C4iC/Me0H3N8se9Y+LvXj2EYbKbbLvbkCyrNtsJ
agGEoZz1Wj1PkUruqPClsvWj+Wf/h1dR/Prl2Hef05kofHTqVXqZKNIU9HecNTbZielT/z17leX6
24u/uwpsG5xf9TlQfQZQemMBefuR3HEetxIsnshNjQ8J1GIB6JNvqLc8f0ZXGiSOMyxieYR6eCpv
/1H9OVAn9M2OPl5DRnPrZ9QTnWReg0BLwjM9aUFuUT2+xHhqADTvBYiRbqw11H4Zna2j/vPMUdv0
TmmPUM+a7hWO5DaDw3+kLxzvT1JIajCdb2/QEhXzBlC2PwKkzgvctYOShROVSI/dTE+V5IOJDXXF
p+IEfOyNZIwQchoEAdK0wWL9eusWN74YJL0qH9993IuCagzQEPepHqB2uec0TJKkYencHJidTq/u
jDsklOM8VJaTiQu6HCf8DHFFw8XxjAukzgzkAPKfwlhWal8rM0c2co2LmpwUJuvK1iBkEkO1seMP
jxyJIiuDi9Yk+WV0wN1NoXK3B2TFuyenYzI/BOlgv1hjNL0wOJMkdpxaDLmimTnOx7mBixIFMAUW
B+zUUgZifOj6Hm7TkGyqjuwmxuUA6qvtgwordX6OANNhKlRD/KDeVrMYPdm1W48ToGZZa6MKfOja
i60EovYTt5NsI/+KeGceO6V9w6laF7JgQkN3OZyQsHC72w6+S8tPsHF+mUm8bxOb5p5K/GVjL1HW
ocXu62iKEK+y8dk0yduNmW2yhzwPp5RbjPRWZ2KNq7Mzf73Y2lmbX22QvE4xzWj+1+pZLGHW8OYn
KNAehdcciMY/NYCOG1CijicgreUvhcu1aokXO0oo2uzQY19JeoZ1zwXfwulyxzE6Ps4KaTiOkTJO
XOu4SDL3rEcxkchL0uV/oXNpdRlR0yIR10z6FThnK9lZq0q+TwZyw4JDgqewHeTQvJJnWvhbvTG9
VYqYiS6YY9wPnQYIwsoMc4j5Q7K3MM6DdLOReAH/URnGmDHzBVPS/pCAIM5C3Wsr0urfjc9MJxrx
BCGTElSO/45fFRiIVEvwg1XCKb8/FfzlAiIPMiDHoAmecJ5dCSqIebzBODS4MIGL46vSwHXg8uFG
XoBZqcX++HGK9DXDgeXwse39m2MwDFyQepr67EUNXAfheAKlPYpp/+knr4UC64sNKhSUVJxLUtpE
d6nA8+kXNxgz64iqxrb+BiPv75XPiGb29k0KhTxWqCmFOW6SCIg63cA8yZS8LYpITOHGFtJPhh8K
aF2DgGO2Qq07qLtKMfydafBtXUFBRCmcx5T6+D6hlULvy8WTZ7Qid4Q9TyADRf4PK6DK0o4MqzSI
0GxtNKdtr8+01uIq0DQDE1FfQGegsbkjLnKsN3jJ10fQAx3pszyezijwYaky+n2fIkAuk5SlfBEV
jFlMy2fDNrpEzLJYqBpT6Dx4JboRBh9CZ7IiHO0wJcnTjGolrzaP0f1rPKvaHm8IsjtAxTZk3h2h
HoZ4atl8hGNT9/0NEB4+eDFN66TCC9m2U1bi1dpQvF1RWvQOas+Nv5RMxPfWH6W0rBfReJGVAi/G
x89u8B0oUQlu4YMwRqsXtgzCCsJ/B0xLUJeCWBUm1NK6YQh8P33K3crHeiIOpK0kBvBOss+sgMbt
g2rLTo0FXvUJRymKint4DnExHKjIk9Qf1S/568Vdrl56xvTHB1is6my6XG5qxljZSRW+oEIIu89G
006XnmdBoMPGHYZg9V43jEbvf8yLbxj2+qss5zppkImcJkG+yPaCQAEYgrdl4PU1pwzxdbz1OYvK
QbHF8lpzU9Xm6jFFdAxa+S+LSACHw0qwFiJXCf7WK3Q7AnNnwLOYXvvi9BKvcjUe1CNrMKyJZfQp
tt8Lzp9WHF2iDSGVwFUK+teL7rljR/xSXoqqzuZcuxWZtzfTYtF6lz9Co54MuiAfbKto+4WvLd5j
AuezYWwNdWBPAhkTxrIY3b0zZH1rveOzgdLGGjkU+hIG6bsKdikkmc9DLnemma6PuRH4Ix4lVvin
vFfE/RiJKPxEpihd4eEGz+faJhdxNDZM0u+JPnqiE0+7G8i7Z+RImaIti05N6xmBnFVMH/IMhRsX
pzL9MJmsm7mUrpKqPUwYYTVKeu99ktzNEfUiefxLqr8PpFMKjbgR1ArNDKlW1X9MYZx+7BiBpgs+
K64f/KbuonGDBj7iAar11WpxXTS1kJAPSQsSilYclfm1t/NUnKecDND2/3RPPh3FCcQ8yzKFFi0m
jYlsZ1C5vPSf65jRgHzJ40eKo+ubHR9hXZfp0A0Yz9HP/+9OUyPcfwOVfi+BRnbv0Fc9J9Vtv7vf
xUL/fIsJN4jSztNlalF07SWVltHx4bJFpf/6XmGLEZpF05lrPa79XOePI2J9nrzNXK0P/Xy1ipLv
eh7m9UcxHcQYPRwh5Oloaa30JL+JYFZdSR9wTzry3CtFQ/erwSEs+0Hd4rbnSVoVjY6zJSeMGxc5
p0h4MClD4z3zpbJZAgnFwPA1sJ/k1ua9GAmDYSlCVh0C4G2oHSRH32lNuolVsj4GUHnL1jzzMNnq
pvsuRjom07a2v/hn0ki24zcD7s4NzJ/eMRXZTKd38RGfVCJCVYtlWkLbBW5xnjCn5pn35z/jJSrE
zve59tr5JpqznV8/2pBqMv1XAVySBHxQb6Ix32CEt9CxtCJ2K1mNMbV/rsyTatTEAoK6afnx686s
Xnf9MSVdREPGQxOuV2YW/fO8WEDeQEDrEVQowjHhfjIcLrACHspmGIfjqd/2rc5s2gQBpR9YALr1
1SE+BoO5wlQJ2I8w/ekVT4r+7QRkV7PjmuG39NUSxEGsCh+AifCwFUB6CsJrPj/8y2X3wcVeWg5y
oPhabC2D5Uihaw4Jo63wiRWixdbYtv6wJ/VSrYdeJ4gW/MuQ1q4tBouKna7494QkZfM/KNUWKQgb
Gagzqj8d/HNHUSqHrfMIdsZY80UJGMND2tmy/u3HRZ70oPfuogLT54QmWjx7b/HJZEzc22i8fRh8
YDY4wiAmBZJ/FG6zmSDBT9ykkDrnALXVIY+xZUUbGvli3nMJTMBtBW47yfBf4LMaN/4bI85Z8A5D
7MqxbzBBKH3kr6TiKvTQyPh+U/7EKfsDkCCp6fZvXwZt5ej3xxxQiV53KbuW2JIv3iu5vRSokvUA
ufaqEFbAjlt6n1+fZzaIww/t26DGshBNsOZpFsL2S/coiG7EriEh4far74DNZAVDdza0x6QL8yeX
PzjRjc3fcYWw4EBzX6ilu1lWlcRw1uiiaEIvQwvYvIOADGeixnBdylX5dbePHyzjQq6P4Uu+9coi
HY0aHABxB+is/WBJ6cCvxLThCf0GLqRy6nn05p/bPvFNHTIrEmP23numZQ80IDNBFwgg92vI4t7V
CLQxONWQOXlLgkcbIZTYD/eWdeYcrvlwQTr4aPrIBfzMoeXYY0nrz6tp/0jzMiC/volaR/ZwFJ6Y
CEwL71RIsN3NFh0TXE66gp7cAk7CgQw0BRhuWiPd4nERrBXCJrjdp0L2XObRlYQGD9tICQG7IEFn
b0UJ8DBygjDvtnkdbHPTqxl59opQaTrC8+MlXcHiwgX5zXnX09Bdry7OdlRQ1fxmCGN3ObGx1fV9
ER3ETuNS3deWS1Ggij6hasectj/Z7BSAWri+WYNSV2f9U7qsTSThayHgv0/WqiHHh+rv4upiwwPr
CXoCiZT2frAeNpC7iygkOjk089VA0dvmpmY1wFqQgmlAavhb9T5SC0M9manM7mMXN70u+q0iW2mr
YRovIN7ZdLjjfbSql4CPb6ZBU+ppXeF+Ve0JlIjZpF/PwemK7A6rlJiRQCqmY3kkQcOfbSEMRsTI
4a+CR9wTyVoOhaF4JKB7TV5xGOIJrplYlOYRjQJD2qqfR+VahY63QM+/squkLsdlxuA+/bKBZ3Mg
VilJOhjVwJy1nHVYBLxObp8s+iPCeEAYDQFTO4IyiIsChZCFaPlIRfyy3hvT/vYXj5xV4otgohfx
Yqqnb69Dsw36C2pewPKQ29LzutPE45jI9yFM9tMvrvcq3ikrkXie2UOQLtY/iVHRxTgr9PHG0lDa
sPlZwgjJR7wPsMdfE/ysRq/5WfKyRTB5E/XAufmpCH39QsW/5l+TNtnQJAyj2iqhj9vRB+sCqE8A
g+D8i0l2XRNdAQEEC5uDd0/vLhWBJtp/mlzvUftVaqHsN5PaLguBB/IcbLC1ooyYX/nIHHfu9tDa
+NsNJiROf0KzsPXc9pfYf7WVqg18rFzuyn5M5Pue+Uz15YLXR5f/7eDnO/nc8em7jehxuyTNYiW6
5ElffXohQFR6DIowX+Shu1xGAxtbsUisdd2kJuXzK4kzlMa1++gsxxLS15mVyAow1zCxIbpByuB/
9ifKpGPRDwKQ/UKr9MKIEk0iRWrbd+2ujabplBUdkAM/uQ5fK3TIQNeLCUPoGVAcCP+e2MeTonBF
gFxgSXh0uQ9JMcfqJiCOOp/w+WlnPeIipVgo08v+67Ih48dJVGPRc5mc5LDkBLjsYQpG+/thtJTm
/B8CkX3Kf/WBINWP7nIDM2f2XPckeZ8QgXkG7q8B+0rnEn3/o0RE9C5qW2ABO09zaDPkNKbNUrwi
TowhNhti9vnAXYX1HXZHl+r+xduvfle8FBzbohTXbhF+GXXHaMiRDMp6PxJwEWvdZBgydaWaqtU/
nToxsP+wC8sGPHewruz2UVEN+i8SWkK5j1VnuBiKeLNcP7U3qdokn8QH6kaAv56Ib89Nuuqf3+Di
F7LnxaL+GoVswrGfmyi6w+wWKaKmnYeyXC2KUb/NkluggGJYlpjfXhaZLt6VztnljYRgywQENc3Q
JW/UN7blX7MODCkyFp79YFgC9V8OIM/oTCsSmgRFabj0X+CqcbpDAXDDDmVVraL234xt+MwL5+yc
xN87F692sMqZ8qdvkpcxAVSeswfDL5crW7QYk5JQuM2dTav6JavzSFk9VLpFaWrwTSHsaIOT8OBX
vI3STWULJ+RM7u1duUd9tNAkM8pVD4k27VF4JKPpntb42d2pMiVCNMMAih5dNpd+6ZhvoM2NhzHX
3Sj+KFquaPm0L2JkXVRnTc47cz+Z/A0WSY5xPkUlgaOsbt5Y1P6snHHDkZiFHUWLmmxKPj/e/tVP
HHEV6kMbKKK+3wD3jVGQZVunHjCRZwIOSl7GeIc061NXBJEjAvlaxotT/QPowD+AzpnkC7JVUxts
oKDye8TTXk/K1Akn/jCaUC23iRGdocuio6fhZBlapCW+GYf5UP8ZdAuVKOP7Rkaa71hd5a6/lOvc
6lqrTJHE8fvAEADcyqSRc2je56zFeGo+0dxWDVrHkWeZYrJOPrafyJ+nNYgrov1JC42Cf3WKAIYW
XJhUClnpYJgpyV7ftFofm3DkZmCrNYjQbNbDvdTIlwvi1OFAq+1lQcn+3HD0B3M5EhmlvThIeins
SAvlVmaKD4JnUXjdDEcGAvO2TMBSfY11CQLUaF20SyAQjuyPFZqVDV4mGnS1nwMbIr5PWU8s/y7O
NnfZSVWgR21T752bkifKKSiXQlAW1pTXDbOOrxyG5N8SocJE8635ceOWUcSb35uQqi2IhlhBEBwL
KCU0ZlBpwhqBXUpLpUwkC5WCM+bHwhpqYNB/qcH/IM5FcXIR8T3NMV4Ek4ZrDqOi2fSNhTmKQxAC
4B7TiGyulB6Ni4X19ktt3x4peeXNT0KKrs6Ra6fp+7wCzpDVMqqZnshRixCGd/XvW6ROh7+OQQjT
ZMDso6Rz2357KAmix2TIx6hgXGhSjbMvWCs7PQEgOVg3AYfwaYFwyF9I9FBehvENld3dwJTdmPBE
ANusx2+a7qyUzmgK6BBmnPBf5mrYabvhLyb3WwI334QfGYX1IKeHiOQFWJLcXkMJwE5c6z0M+odb
Zj/TVfQOSfnbIiFvkPa+CSn3XmcMIspZRy/zUq1ZafZW+EPihPJo5jjxamznRZ0WeBRMtRBiJuXl
M46etoOgTcsihFUbzJceASOEvnFCYb/DSvCAd2y3eaabtIo8hhZtslrtg5czry9kXh1s3/GwRaZi
HxJOZOADVz10Hdg8rZo4ESsPXBwg3N6R461/A6aMHBE+pkfGULQXiKvd77MnI1/ytWL1PmTTkShp
j92BQtwaCl1qp3zj4BWH1FlAAKgBGEjhdu9OF+7v+IHMWUrXsCrznSViDz48/GY3l+oKxXyP2vuT
hnSlAB3y3sykzBCG4gd7VFBRu3Lfw1t9fjqG/uhY10ufMAwwPYAfmEXcY4HRWd0mGoewNjO+8skV
E6LsB/nml6AM0zdha2Ekya6X7nq+3kexAGjhNTo8Cw0gbCVDrHWiM+3qqQGs/FgjTW2EJQyBJi07
DTNvtcbCGapuhrj8mIp2bit8htUte5RenxfOSCLvlho29CDeAoXWa+fMnsAgrcmRMLwXPLdpvK08
8Ab1pEWDvsRE3wlCGo/E82k4qizXi9LjhZtQkiDTOvLqlA/1auE1wFMhbppDlnyqa+yrTkjq067/
OrOwdyMhU30ia1qZuBu9NljpgkZNbWfEDxmjMiUhGC5BGvQnmLWeGGR6XEJKUFuM0qnR0cU5iW16
W7Jie6wAe9M8bWaghd5nNTMQYkG/1DPg7lMwUPIDzQ63p+U4g8ARZkldesbZqPiFCuhW58J+jWBZ
yNdxenxYb9Xdw1r/re0NWXBW2Db+z5MdoB/nhGi5XI1AXiFP58Jv3+FlGWldFK9U+73dU+6zUlDL
4JQByXzDuCcB3fGS7DJAxzuUCuT+rvYYrp74GAhUyty9IAYeigXJjaYvWHWMG6g725DBFWaf+lLJ
EO55G+QfieUaHijDbITtGGTmnWRBCwhnC7Q3NeKfo25k7bIvknqLTOEM9vEzicu0iaiI4E59sPSf
hxDWBbt3Q3ErefYvlNODqFBk8HxA8pieFPMzn3TWmclLoHg32MEYXRLZVp4RQjm+gSmEpeFsa9Ay
LcAPWRIA26aYGCyPMOMw2vVJ4o0ApPrBhZhp7Hg31l7zaP+w5Avb4ShKOnonJslF50gklTK4Jyxr
aIAUUG3y5FM9LaRW/njQlxT6W3yXqN3TsXhcqAMoMUmylLIrFVQS/eOVCCr0lahkgy23TSfy0dOO
2vEpVAumAzR6I0/aHQVes0nSAt/HcfQDsJvU7K+dERKD324KYT+tdZJ4L3+KnaKWENUOePau+aD3
pNz+NCTOrZX0Ymx0B+lrjsctcfG6MHAwJXRN3qWGiEXyHo9Z+90PGwutPiWTDMLsnx6523EajEmV
W6J2ZU66TWsQ+NYOA5N+/3tD+tTMTlPPTMKXaHrzjz2I08902753qDS9aAU5nrfdS3BIxkCE/Kon
jfO5UQ2A7l0gWOqpXrvjQlreW2KHNp526aoULr2UDgwfXzd+HFavUEMrtJpg41oZe+29fKm2qhH6
ENcb1a5BQP14o74s4mcl3uFyTpi3mvLxMSlQmVRj51pEn2EXxePUQ6kF45ZydJyWJl7VxBCRgJy+
b1U38HQcrEwxS0+C2LoNtRS3gM9iriqEcf5Q6hJpV+Mut4KonbqQ9zYqCp6tuzJcM2hi2iY4lW/A
d4gTiOzJR3xWGoLDJEyjux+VqCpnhB/y0IqZKQ0EEKGsCXA6TO+oJqWylYqD84iZwOcLotiuRSw3
Th7H/i77zrNm8am5Qz7h+/1wzTCWopaS/jBMkxbWiOxi9+r7diXqJCph/VAuqUYolBiGNSS3GA67
m40ozwkBcJ9PZtwcvHfJxE73dTlzb5gX6LB/amIAiEmTOMi8KejoHDyti4QN0sVeGO+bqunNuueq
X1kTAyPwmnXse2fQ4Film7ewAiEGqmUKHuqRMwlAX4FIVbCJeJwqD+gKC8lS1iWRGvBmqLBozr6t
Le+vzcypO/MmSa9b+//5hCU09c9b720qRulvZdur7/bfyc97Rn4YjVlvjBvpCmIny+Q+WWG9j48C
bMhSwYL2dK/uFi2EWk3aJLFspVqPEl1IzH2R311z3seaUjxlmhOfypBHAblKZVM+eK/bDUC7s2Iz
Xt6kYD1cCM3d8Yasy/AaVoc+ixxrRlYSz0gbtrv/GQECyA4/cQFLA2NfbrptWDB4VsSkMtF4lQY8
SuCUVBb1R/poc/dBy/LcXkVsNkiy5vSFciuF6/ZcINzBS805mQko4p5w4iGWJ7wyYatxigdgCLWA
bP4PFWeft9IEsEcVVT8V5HZrDgEV8ELhMkS6sujAYFoBio7gO9N7Cqwwzz1e+678+oGwy3K9GKr3
/d494Ja637WurVFQ4tOCoYgaLQPTn2j+xWi7UKAObgyeWaQdZhi3KhjE8RrBmXlrSm1z/zlbgB4M
cJv+K/wKNJ4mtSy0ULEEb0l8k3487RYkQPMCSjnWh1cbz7xy/lqDjf3Et83nFaeGDrdZ1CpKIC2l
msNmnNL7fGLLmPDP6PdzdLqqaThyQWOH3xg0YaPtBRFK+1c0pmiC94p2g16fRvwYAKD0BEOsTfBV
WAK33jbxNtD5t2dj8lokhwY6uor8RyPzYsVRuGTXoJ16hWltBGBRItl6sxgOS5QF53ToByBYkcNS
IesXGkWSZhtPp5IwFKv665nWTQb2hfhWiNkeCbmThrSwG5Cr0tQHi5rP/tE+bFkfmqZem/rErk1y
DdplfHnM/SZf58JYl/GhDZcryvIF1MJ0qBn2zODexa7P2PYGkRaSvQg09gS+nIVIG4P9AstG5GR/
APZzTrRxpVBZct2j0jfk56bwMvi4S6GqmOgKnvj7LMYUJN76rgSDaZqtLgctMkb5hb5hIhLVzqvp
P2uRdxD/1sg0Jp2Vzw+XneBfzlcXMlB6KA+q0afruLt33dwJHrmzulvvYPtraxNuFyYh5Gp+yUHT
BRA1475TpzkUxzc4EamUv1iUpKi2QYLw1Y2B5TpiQCSwDa2RsJcKqSi5nd8v4wK3xOAEXY80GDUu
vh/m7w2vTdmKMx4M7xNkQ9SO/qN84xO2fokURwtBRkgbxJ/nol3R+2kv0kZBySErQN882R+ms37R
JAyIb8lfiJv2xkmJbTApgTZK91YG/nCfxGYwrY4dEAMOkY01hQb5mnNVpN3wYxKUR93J3KYr/UDG
ckOKT4rCRFxOP/vQLj78CM+2k5teT2YoASuGbVCxQxAIVsovocwix3MV5Xe52UyrYbolpDEhPw9T
calQzy2dUtp4UK8lPEB2Oq02JMMaRmo7yWavHkQs8df+0+EySDQeToXnfwTPVjyCkYvhRlbVftej
rJKxIY0mODcivieBOxxCpdwFaa209IwmTNvEaduMdM1CHK4CM7qcy7YVX2+cwXJQCo9hiAF/dUI2
ILU9jMYBlE+5eVIGNtcWvjGgwHui1nxHXRMT1bVx9WAKNuTc3UTLxzH1TXE+JgUFi/Jkaiav3EQI
H3QWQAQ5Qkd7BUfF+yaVn2MgAbhj2Vi4D/rX1XOt0nIHGKL/gUTLEc7cKStAraYqvFFW/HOWsWFn
5E/q6rEuaAtWPYu800K43f+sLGexn+kr9Fukcdx2J16bqn5kjEaCMp/g79PrAZsFARWW97CpenN7
KIHILexZnY5WF2Bij8fXAbELC3c1zPAMrH1MyfpjFGBPq9lyqwoUSKCpj5XW1n5IJSuRQUbnRtuK
4VJ8sPrNINsxCAyNaH1Ze5G6pbiFqUeI/eRM8nOuwssvqh25Podj7pXs67UeZGRXlJnNgpmhByJ4
LZ573YaK9horJyQnD7S6pIfB69fnYfXj7FTM1MlQQRwyoM+NZkPzy7Y6AFKSESWigU7/nGjM7b4v
0CajsKwhISHPov+83np3voiAXmYwkeFvpF9b8QD5d0LVicrBDMt5xgXCdQbCl9QN3QCmnTmN+M8T
KA+I23IruFTF87Y1ETk8mlWq0u8kgzpqkFOBIt6RsR941HUjHYZgcTW9VVR46EIpm7EIqT1ubDhP
/VSp0i8lBhasok48qPbE1aIZnOHyi8oqH+mvUdbMwUrxqWvYdK4vDC2VMBTKVmiAvLmzrezOTuDP
BGxW1E8eCupAsU8I081cyjCkmU7latx2o5y30knKltlnJC0L57eu+Y+DZKh75VCd9P1EMBLn5UD5
38/wOnE9cEr+WeB0riaQ9vVpcAIUZ1llBE8ef6mCdfbrRpnKU8FYC16q7CrLfOR5iocwMQg3eQdf
rsnNzGhHToKIYS/qXiE93fUYNIVfZC18OuNQPlmm05abeG8wp5Nis7KZt1h+LOXoETHm8fgPc2Ax
PCkI1JYeV4jUGZv38+AqLrOp2QKxXLYxnkGat3B8fH3sY0axRz6Y+sjCwRNyqpnoEF7ecb2JIuoc
FESfI4M9NM29En2Lme5KPqgmSuKEOHuLlUUv+C9MVjklPwPOZGz6WiRfqCXzapb5+1MUUFSeUuBu
OPdVti4gl/j2zhjyQa3WDmcpsiI7VnzqYK4RBAQvzg7Uz2XxUZkdmrjQ+k0yZ8/zDjsJbQAMkC6s
nENM2CQFjcCconJTigrsOwCsXvv5K1Pz2pbo80zKS/8ai3KaqW0Wm35WzcY5DBUmZTOjchC3a2SS
CkBkZ7KZlXO8OMLm8NI/SuUkI9pPLaY6yiSsqiMwCO6MEAepNtFmyWkDlWqSgkplYmwECcHvk+Ta
AWD0HUD50i3VxU0MkJ7Ne8+LnoG35XfxdyYV4H6jO/X+NYfGeiA4jwMesgd9EFQPInCWEGG/2usv
ZUM20rTcYZA3SRnXCNCLiKWlLBsg5EvGlekbZfxgu18JGshURZPz1QD5zfi5DZu8JvshgBnHXS1c
eX1Wuz1gI70QbW25+KsL8U7Atc63Rnyaiabc9daxjZVruoqii/ljeDFa4plu6EnqtC/Tou7FYnac
MD8qoLRDNG0H0M3m6/eLev4JNmTvmqNFxt2cDDT9D9n9vkneWrsVFnBUr9qq2XAh0AxwmuJhe8oO
e1QoqdBB1m/QfQAWCl9W63onlyeY3kzTBjK/hrgf9mcyoWWDnogt/2ChzbT2J1Gx/9ML00MMNDu3
643m7hnE01qf1vJPD4iixKtKPoH5tZdxsTpwta8wfueGekxdK8vJmi5amadXZhSOrvx38hkYtSou
8+zxFH+3cCD7+huaSU60Or6VzUSnlMKoK/UZ2ZMhDAXYmIsIjIK7KjOK9BNahORD8o6A7N7ofXRs
1xjdLqMxKcePyIIfnhFxFMixC8ej2UWQ4k8kkdvUYTsIGjIGx889wLvvKKryE5K5SxUQBAqT+FDN
7qf6ki6UIlcwkxItFO7b31GrrkcgxaOcuNNtZ/Ih7c61OrFUaln8o4UPT8SxpnweXYfQwn26b+yn
w4sobj5MwR3VIkGAnzGC8hLOPm7k/xbWxNRfmKgcr5iP55gCXEndYir1S++CwO5XPdEyX4YKDwlx
CzOxTcSwvxR6HX5E0JlmYLAUu0pNVbZI/6svonbl8g2ZMG8SOCBkB8vKvVqL8q6VWIRNOZk+p21J
YS1PjODcRyrbvSg3Xw7a7YZok3wzCXHr3pO8GNFLqIR+NoVUOdXlcfu8SsnwIW8CGbXhqU8PcCa+
OSPFfDM1CBv8F2sDs+cr5qD4fNlrR9Z5eXOs1wSeqg59cF1AVKgrKU03iQv0jF41J48vlTawRTHT
cyIpWWDQ9zG9kgTZvODzIamnfQ1wzNSX9GEMCEgnpa24b4ntFeJQgUandLYSWQ7tCj9pww+GVlv2
yLwmFmiw7mBhWHGITwrUoBGBeJHNkMEilrBY2HnB8c/1tpWYNMpyZFH7z6XtTwU3tdgvq1JXXI/g
qtBhUfScjm8YqAiwZ84zFeR82znd8P+NadKsCUHwB9RZmsazY3sWjAzTBd8jX9f/nZbCGgUSds0m
zP1Wv1MExlHfXVuZq1B2ltWdyRIYVa5q5VZi4IGDyaMCka34HGJ22/bWhNLL1P/lhFWX1iqWeAmK
Ipo0oQ72hUwYvpCuQxEnhWyXAlDkTK7z/q9OteF2oid6BHeEMpH5T0iHzBKZmjhCliPWtfy6pWQD
crnl8JuN3w6TNIFdrgYEhDivUySNU4xSvA6v9IVXDCSc/pUdfuePRdAf4SNPBpCS95i5zcEJdsE1
meSi171NXDkYLXr4QK4revjSj9n8UilJ0gqrUHTtxW4Se7zAVBFSmVk/px9pyCo/WEEJj+vShlZP
eerJCYPKdiYOcsmHR7msVhb5Z+eVN+U7xfpVIv8m4PxedzhZmhdg/nErXrwIXtvEXa9UPoHiDmOX
+MaZ+juE+1lWm/RFAcNB8+mF1mn5z0kWfq7txoFnNGR67erCwLA5f0mZXb2rZpZsB1E7uEnjiLbU
PikLodRyd6zbRWMD/5lsjrt0aWHxYspqjpidGymcDfagrwn+2PWWhem52wgPkoIK9c3duou7+Lz3
rn7Q5Rvm2CZ7k3nfl12S9NRiMHyeN62tbNfEh3EAm4nwau/jjhp4Uc/SsOXb0ZZZPsZiNVmeeW+g
F/FiiJ91zlgS9jOyjR7c67yXjWDpo7ibYAKrDCWjNrrn1OJKC6MZFUoq1Q3NAE8piikPA8EZCPAh
0vK4RxTBpjwlH+H5DfMTu6I++zmKRNYmmEtYzxk9a2FKXdsk0ZHjBiAXUZdpErvFjCtxj3stgY3R
paCoXMUPrYFMwZovkD00h5vmytHTeUIcpzOkGMCow+gCXMadZcQzBBUyVYS3n/EaNp6O+rRu0sb/
QNIEKBumFqBlKiNBeDWRexx/cXJXvZXzLj7Tb+emBz4Aks0C1RIRLtuUS6P/lkzttUGvzhVygSsx
9GPoosL1ezqzWu6GBYkfnqRJZR1F4FBJdXIFzoUd+nPfgaM2cwegmMhfwNN35L6EFv9AsjJH8YCt
52qUj6PNc5CFBo79/+m6MFJ1eCbAYdMRJB5w25NoZa2iabU7GGI0eJTIeT8Zt9gCSczXNMbt219i
dAw1l16t6CiEwNeYSqdRMdsO8mNrEUZ0bpAjotPZ9KkRXQO8i2GpgUxkJjQJnlg3x8IrqlCveHV9
X/fN8lTLVcGT7Tb05vs5Wr7S6dnZ1a3ZMfMEiWuhjJ5wW/7zoFIVIUL5fLlMJCJzGqij3BC+ru+r
NeqBVaTF+lUXQBeP2LmZN7Y5uD8p4z9VQV/LhXbVBSIGPTNwoFfQbAdtHHcX6VrjhuPYYTGxVUJa
RaHBK+AYMu9llnu6KoNsTspz1S6DLM5rfWNHLPzq6CqCXZMfeB+wzmLVmJ36bAZDWhRm3apy+iCk
vo7bRUGbXA3Nw1O+l1MEvBEw0TIFn0CsF3n0pu3WzXgYo7Wy2o5yQP2YZEOF+uBzGo0QAV2ExZ/1
5sNIvGI4iMx+GZW1D+UBEKm+xe2pAXxhPpv8/ByeTtInnqCjqbxnkemeCV9yF3MD5i6GyvVG8oHt
Ns+4aOOvcvxDVOySE3u2e9on+PZBePhpV3vv83f4qyejtQEUbmDHiV72cr8JVVvum4RfWQLej5MF
xcoXQ5liBcSU7/zGz06Dz5RyaRxFIzZZVkIAMr8r8E7+OuD/Io2i7psneaydmfGJwcDwnlUhjBQF
/CO1QCvvOXibT5UeC7cJkyK1fg0rSVIfxFyPcQspXTs500N5F03LTXQSjiT8i7Av9HyxkGXatfZe
rLgi0BIgQ20IWxpytCjjRkONdn7TtxCkK0zW9IiTZPZ5iTQ/JUvzvFh/guc5J6p/RoI1QIrSdesu
e2ksvRV7CIh+vmmsCS5KgLSNKk+uE5vHaTbIyxppIdqazkcnBmfuIsmRIfUPVM4pqHqKkoPIkEKI
ks+1yn2B1Ami8xj6U2XAZtyGXdT4OONQCm9eU9F/PDALugoQ1oHJ53nY8TcBFHKAepT3W/FfqMdV
pFLvCGDZ7pqgq2HbFua4k3edbM3t7Ksr136vyMBD8n8xQor2t9N2nO6SS9n5MXKjfBA1Fx+mqDpC
8XR4/h8rS7jn0IjoLJBeES9wv0JCkQfOVRWWchJnNwp4tyBfTz18zdEaKndUg5O6LyFZ4c7MM6n/
8KUhDanAb59R8mFc82tiuIFzOke3lTaMYKCtpYKwdZim+GwtRQjbnWJEUtzsT7+nA3en1oYAqWcj
VNCBZ+1sf5tdm2ErBSB+GsQuNEGLMQjau9qrfq/72DSRyAE6AXp53G7AzxLlhKtw59taks56cEXx
kgMgp9J6MvV/zGkI6QNCAaW2q0CPBSBQDaOgI6u2/tUDRNamL280wcusNk6nqMPQfa1OVfTtdAQT
kxjk7e/btAmCn+IiQ4FPFr5uS4NFugyQhbV1YicjZGjGJLTz/j5MnfcCmuYSu6aDKgdsw7WUHe1w
GfjVeymesMMaDcePRGxOYdKAVBoLxrnz7Y+O/mTT3htuk0UxVlw66idDTAlYcv+Sx24XjvCNV+xK
s3y68zBPnMSc/YkcyPT5rTjRzZ9sJD2Wpb4wUgHRWaW5fwtibRd3IsgSmJipZe3Szs+6UUv59cXE
FUglrfWVVCqltFy5xhE/RsLWOl7Tt0s0Ns1rhprj+F3DLdOHOKaf0R1q7umpGXj+4lYetHWmDuex
qSMkVMF7oBPHZdj/QPzYqujmE6mZquN6PZL1CBric8efoEGYXBI6XCYZyhh0Fn0KzWdczMPDFT5q
MRb4PvHbNnoMyQ7oCHXOzs5IGbg9aYTHpAAuI+cUvGmOPqy/6WsnKTaRtEVYTgFgY0nXXz3Iptyk
Ei+4NRzxlWPjLpCKz3sWD3TqBwrnrctvgetLb8Tli64Go1+rHq/LGh4QfjxGGGOVKwrScMHXriHY
yX4dXxLhdR0ekxWbx5Hd9l7maQgZ3cSdU5OYKTxJrbPKoemRhrmPAKGjyORIhu0czZl4TkgtBcbD
NdvkHNUYX044xkpARedHf54EVWLtVIBuCGNrrk4x1qd0cd6xaXAJcbGj+/KtTp1DJlkMmQPOGAFY
RDqo5i2ZYxzNfwta5vJV4bBOUoQnhM6OvlC239TVtRMYOVJq4Pky+CPLCRn3BRlM9kvX8R49wNnD
mgRPJTC1Ogt3jhg5CLOhxI4I7vz5/QqqpJb2JqHdkXIpS2YIGADY9E1qrcIfbUoRs5j1ml9aQV6/
iGAaLT1bAuAORubvQJLbOZCSOo0Z72Er2m+H0UPi1nHCGQ7p1QRJhG1byATy9RFYx4ZqVgUQfQj4
Vli35CiuSt8yXlDJopPjlLwPfh6VrMzlkcn/GVqeJW+n5bi/Jqb+5ZfP02oqBVNO1do0qP1l/GuO
G6wyMNQQu3dAsUi9xvuEsJH+GOW/DwvbNYBhBFXMIVHsiNVmUhxvssvNmvkHqZsJRF7Ld5qBBDWV
b3pBG/APZpkJm2lZQ49QQJCy98N//2xL3TPtgUPGJm3qa6sNcTFw5A89SqL2wG6zcszMwL/K3NAv
xZFXsYC7IwwaTPj4NSTIeTXQppEoYAW7ksRs3W35ToAlP02LO1Zxb+/hTzPU92DOyCL3aeyT0iPg
M3sA+A19GYmwKvmabcxlUNLDz6ySQ6jgQcI708FzPpOcsIxkEt/LQLhq+8UQQM+qzu4zoV8GWDEp
Y5uYdnV9QslmRKOxCZEifv6ptKyK2SEin+p3J1yNPwV8r5j8S2nDbcn5blA3pPNgUFJ7G8obk9vx
TvUtJ9lLneyTDsGl8IBvLeG/ddu48R36VL62S2wsSFxQwSarl4dYZMHVttwtSJ++DHwNMg/aQ6SX
jdJxstzRvZX0xAQPIEGIY3GWx2Kxu5yPoxfLNRKauaeyanfauizoZ7L386Jb9hYJfvrhcToHFhFv
pjtQWJyyhyJyZZlOXCEIiq5HyIRPgMSmL8EnvCG/E02Kx6xwvnzOw5ODOtnSkkHyH5iYSsNxu8Hd
0Hln9Ow/oPXPI7WLteMtvhZ//iylFvxbJJBi/VEKfpvpxE/hWwLSE359mfKqrBtS3jnFArI6nVIE
93iqbQNJAeOqLBrV6CZqs5vrpv44uWmLg8ZRVJNAMGdhCGIzlIYO6aPuW9Bz80zWiCKnaRADUMiv
wV+4qpbAzUseByHyVWEa+ZkN10cPI0I3SAhj93ZLmzWjbx3bSlt3bRt7WwMkUsOgGtzKCtOq2jrh
VFPX9ae1EYclAiSXoaKC4fDbfgpv7nIPsnAXVQ7X9Rug9gFz4X6DyjlZvn+B7MaUJ5yrmoIfBBnT
kkpIGYgkxrxSzg12iHqhmghXRCadAD0BD9gx+Sd39TGNGgfCA71m41IY5irD5+nR8REP6bwiaL/N
x1JaEyC/CUiD/alQJerYZZK2aI/m6o4Nkoasq60+ozq8acDj4wS07YWTbysiMYpkRg3x2qHqpWkW
PaEAU35u0qmH+ni133qzOFbTb4rYFcE4XZDJQAgKe6nuVUa5yhKb1yat3SEfUKu9LRMZDuISivWb
e9Tx4ch1S1Vy6f2ITUvOaHw7vaUJQ59iEEyvjexYx1ZqiJ6T1bYaHEVKTtJnlMtxNblY49iE2P52
9DTUKHn3Dsn6HOs0rWZtt+LzQEq86DHsQq4dpMcYrsbJ/UT4X+msySj8m6FcoCPLu6/Uo59Ien7J
lwWPwJoRWxBQQmjySC6dXFby75+FV8+umsUwtgxR39+qE5s7Goi9JzJCEavl/kJllLl4vfMw9TGL
3/Z0p6PPeB+4Sdc/PVI3ZrovjFYDWViuwgHWGIMD3crtgJ14YsFoQuGINLH00U9RI+O59XQgThRq
XL8ZYyn78PFcXKr54P4E1anLTGojn0LhHaCJwD6UtnYNtS7IADXV3nIBClLZdFziWuxoPAJKzbxK
WxKsJrWFJYxQtmpCfi9AxfIJS5YOzEleKGLBJ30cKx9KvN7bMtqF9jHMofdTn1grJeuWXJQKB0Xf
IXCOUFUvHOFLJG50dIjGhcMjQhcd3z8lkLoTKVXyVBl+FWp66uJaZvS3gsUpJJN92Ur3P5xDDnTV
/K0LM38j+/zDZvI3DYx1w1deAViK6MOh8w+GO2I1mOx9Z3Atf00HTvzvn3A7RlzQJv554ESrc8Vu
lmoxSwnJehH5qkSF5Ou3JvKV0utMvr88Xd2NsNd5s87YfrTjXiTo5kiy2ufGdiwsgYLS4xAiZ1er
Ys8BNPUzqA32KQQ5bfKbmy5pE8NTKdBC1Ul0qmEZexTU/Eg8C74gsIRwbtrmJNnVbv/PpL2EzUAV
vBNgNcyD7zE79o5Qd2finRO3E5fa/p5Rza9NQiuImPNm4TTAa78l3QouWh9xf8UW2mQBhLjMdLoP
fPCJW76dsIicOVTG/CnMQnaYb1PLZP35+w4KgLmN9wtxDdKRyY1bLgx4mdwlSyupcwUDcWp0aVGO
UXnfiFCQVyJSJEdxHsCGBg7nfioJvmRc2uYggtufG6zeDlWel6fftVgJeV9XyxMYxVwatkLh1+3f
+4OfB725S+Z66unThiA8gSMNMwd5qEFfIuuKSyLSHDgJJeCZf00Ec+G7eVIPsdVtvInOWv8QXtW3
bXOlc+NQkC7eSuzPKTRpYgJgBw0xq+hQi+QzCvKGQcY7el8T2nToDHkCQSDQUilnQGcSOQLaysk4
Bl+115BCeUfPKldnbz8rU6M1lP+LqJIPdghPXkCTOllLU7PS6IM9PXlvfkQpnIrFmKCPYM7EPKQb
MnLHqqlyiGY4ln1ezPcobygIk9nCQ9hNnHNCPgkIlDUyi3wzntHei16BWXGKArg432vqTQby6uOR
pxEBuFLwXkLt3tBtmEHcdRDrVm+JzyC3ZUigf2w3vlBdn3/a8mBb55cbimcOsvmn1z+kDaEAvthG
WN+jMYrsCD42+bPpv9HLuUf0iKDR1Wzyx0ztvYmcVtN59aD1AN9qzMoeQycieJ1wxalpiSDaPdvD
2ztzcke0WdHw2dkwUtr7KuaSY80aohgT5FzYJDPW96CaQrQqDCdMCSEB5GAIv6akQqHWBLqQC4Ql
51Bmz9w10NQz6IjGRa/ImP6fNqjvXc1nAL9hRr1bLUuDNK93XWGFeZQD/Ya1tDv6wk2h4C4qu/Sy
tyIDpX6+6falQco9nHy7GDTF1BF4xtXedcdMSx6EkjZpHO/hpU1Hty1aGA9jV+MYm+bS4T/IHvgk
B3aALD98pJzAhersp83uikwdVlMC519FQe0adwD2+v0D4xPUZNrWfaNsLwIxlWSIPLb4huE1h0S9
RH0r9RiZNXQbYp6WjIO4WtBI1vXlGzhILgvvis/zITLdHVnmxzODYwbQXoheFsdL3oIaRZgRpZdC
A3LxslQLgLVgOpZ0fj1mNafsUdxvX1IaQmt3c8E+ySszlWGtgzGUffSNTXxNa1DWqhxJ516E/MJe
wDLphP6l3t+AxUG7u2c2ClY02Reft/gjA3yws324Kmyw81eEUaGmzF7P+GWq2xD2x+BLduj+jTEV
YQ6b292MQGqIrkF3u+zNIdewSJor3QBxuJxtdA8BcnRUvJSZANupjyWWZlzxvN/m1/IXO5lj/czW
MXOgHPDP2J6uXhw6+JjdCNJhfYEAMiT8eHra8Ym6FizEY59QYynnf6BUXysKy89j1hslmbVSLmur
/TOh3IuGWFlTMxXOKi1TTJlBbz353pJUEYAn/NogGRPxCXwzR5zhLw+N0ynhO5cdFv0qTsNhUIkr
vEKEthUdauhzF33hU+mNCamUBy/fSnY5nIRFV4BEO5TTHKQb7nU09+LVUuhyzElA2X3Q+vPiW9wW
JBftW2cQYCjyd0cw+jrYHk44DGGaHNVGAPt08mJHHgM+kW6WlGG5hUDM6QPQYZ3pV5K7Rt8oaMMm
RGVNZISOQ3tkFpkHwrDrlahDT8KF1FrozNpkIxy432tkmRF/DBwwjCtQImeKIAfhLy/Xfrzrvdye
v0Jm7rORZHDbepKX3mW8UBNcCh9ZWp2jsJiMBOX0ljTpmm6RvlS4LrwTNsgmwxwpVCoEv+1/Xun2
UoPkAj7/S5bXHwteG7QBEX/lIKw9zD2JVNKKilM5EEJFZIIP9ybsZL6fw5JejeI5FiHUsVCX/jai
uxMEcZa0BZYRMgrNIdUtc0GTXx7UBi5G8Tfp5QKM3GF41Zch3etE4lxfoLwryKt7P38dsFfe8Q7U
++OKZBekx/cWBuUZUyHmug100UjIbwX6pvexf5deIHioVV9OapMAmqzesJKvxyyR3X91qnDFqp3E
7L3UOFk13GxfOAKfQHBpqZ7Pr6h66XF5qM0+FhRHtPToj/oHC4P7IytPVTDuj+A3Nb+FopWPSwCO
1bWs+wSQ4ZOs/d+Os5LKXPREgcxM4iycye1L3MqPL/NI1T5FRYSZuIZZFW3AYusoj1iTtiTDlLIW
bTSUWR4qAqz1xmGiexuScplGqOm4FXN2cyFOfYsBXSzDdhIs9cjURIkDMCXti+6WVwmvqW+6r98+
BZRnN/TePLwxWFKBxsemJhwSAgZgjxE0PFTN7UOlJi6yVc3YU8t56h+InbPqEqzb9PmbEGNK67CX
P4R97LgKdWWWj21NPDmQrqEWrHFGoKjvpqq44nsmimkxjR+jA6EC7CUVyDA3dwJshm4RzogDeM6f
/g9lj2JnDFMDvIY9Nf92DYeLGxqpOr/WFayX7674h1Z23UdeXcB+m+fgSXH882wBm4UqifzzgENf
yLg2Rn2MlBdDofrDWGqB1ZwzCT5e6+70mqMTOOPSeOGwwhMQUG82f0e0L9CNES/4S2kJ2BlWKfpA
/iOvL49zVlps3ftOaF3uHaCXN4RqEigXJBLgs9VoF0IADzgbSeHIioHcipoyNp8tpl0EeLOX37TV
AC+BeWlCDixY/gWonyvT5vzLX8WEJm+WfoFEx+zIx7Do3yCWz+qZgInaOhs4QIxr3mFZ6XGJh4E0
SjmQVx0fmkbAkH1E6UsuNcbtx/U6S6Jsk/uXScN6m1FaEPM9DUO0Yc1uc0pAz2aWrv2uLlcGjAOY
pADvFWveJIxyuUwEWLwKPq9VCDBZfHsi3lCTq09d8+bY/8Ir6pLta0mDU2xCc6lGEPuVQZ/3eVQ1
znPvxGB26I1bacTCwga5cLK4ulnJuadWnpviqhkacqhuDxsstraZQnB531XB1w4QMp7OZcf0nOSv
0DUQ+tim9ve+O6s5eoMV/0pYvEHnY2qyxEqyoaD1LIBTka6h0OkHjyHVT91A0lkWlZusqqi25e2l
qYzoObdWe7W6fiDefNYcODrzF3TntDwKq+irVaAJxMbk8auxyJ/qsECLlbXdjVhqzuYj3EbuD0RZ
jZwg/aabe4Wf9M8igOerwTIn60q6rAgasu+bpEBeheSYSMYd49VzKB9fnvM03PyGDMGwhZdQ8Ooj
s72KSxyFz08fuTmZTLH4YIqIqlmD2D31AoKvRbm69Gp0c1Q41MKqtjDGYEtEcUM/CM01svVNYykN
DMaFiYERzZ5k5qjmu3Y9ooFWS0CI3RV/QZohCBBOar5BHlNrz+fsEVDYWWPsCZlF+phtvgai59Cv
yKN9EBt8hT/434ccXruVcRvvacr+MQjTdlgfK0P/tzZd+CuRBkNsS9/pPL64cDUZmbbf+v9SN13s
6HinLlA7YNi0yYNupgVeX7lKdxJ0N/mE8fK+x6mZDCkheYo5ZA4WYqA6NCK3/er+Ga6AoZO154yh
7+s4eUcG2aLu9fydAHLHr6gR01pgjHXfBn2xCqh3v+i0CF+3NX/ZVAoP4O/ibYCAkZnNIcYTWEOt
v7IeJV/lufjApE95GKgW7OD//mcGbLaR/OAg3HTwuF2Vyc9zueDFJJi4kuiNBJczJj7S5qu/YHWh
+qI6/ZAQ/BoM4CAiUgBmABSi5TWEO8pxIC1CabKtkN++rCIusKRAv+VA27Dc7BN1zXT8/PeIR8zy
RSgSLmVVK4FlSyXOgiy+91Z39d8vg4790g7UL3kiF2pOYdAdmPavZJwMsjpRKe2AfSKHzM6pVZnr
zjlumLhrEaWq3iF6tb1Zi4EuzqZJOxmBqjlc9nNtVEmm+nU7dF6F2cxeppnPQd6TWGg/YNhzUKN4
x7A4wR2SDTDZZmtOWke4SOJgIkZPSsOkhwU66g8h/VHjk2mUa+BZHnphZDeRmZ4D9tZjgqseAEQx
MYa+/F/bPxpBYZO1bf6DWMnDg/F8n81RB3cuaXcnYDk4KO/gT/a1YVRCoVOsubwYzR7+6rjMGTX8
KIvpd50pFfExevb0WgV0IH5FECL3nkV2so0Vc/+PvkJl4Xbev9g03g2U59h3VPjFizHdH9RTf4UZ
s8ilqNF0yd4x1NKyFs35L0nokZX0l6S5LLEj0ojsf/iWDYfQeI5/ChU3dFysdhs5nbljrsGpU5Jn
A5wjXFwb3k5ISUM15tN9oGYKb5sOQfkFNMJvjeez6iNv1QAE7JjumjwnixGw+T4VfrJv6dDX7Avr
r2Uz/ahcOXrbqIupoNUD7eT1agVgPP3Ebz2I5edKB9tJH6HDGoykD+EcTlMDM3OGq+5/vcafQN+L
oIa0MPhNCBM+KQ/jmuvvkn8i9Jp9JvTN7g0riKny7AfHw1m7Z5+UU4rmpbriYhAFlxkbXqqjrVPT
mzN7iaIwFJSxBBmSGBbPYMKe/xpXDeO1GIrWlCSvAaYo53mG8tfc0T6fUdMGnEqZzngngUPRxqaw
rMIGvCOuQ/1gfakOhdPKTgSuBQ7N1MpwX7RLFBfy9Fplf1IClAr4LsHS8bTtZbtihise+ZGpXtLx
5QyQTGyIzE0i8QiK5fB2Yhw80yMljACxI8l8WKVT0Ss2R/LR7hCqKTjEcQTxdgK2Tn8S882HraKD
JI5ym6tNx3Jy027pSLYpmYpjZs18/lXXVdagmPvN5Jlwfek1zYPZIOXtY9vLsnPyknJW3PvMjn0T
NMTZL0Cxjbsu8NhiQxUaU5Mizh2aAfl/hnzATQGs7wcYbA6rsEyj5iQEFn0oZKGEFxWTepFpLgZ+
OfI1+Qczh/SCIfzBm+UoPy09x9L5SI2vCizG1Q/xdrtmT7lbvvAjrORU1BAi+0dfneU54j7RsxY9
u41sBBiEoN51R6Usss+JUVb8UgJ3WuYcacjzcjKbEgdtlYJRQrt5vkcaTXarnJfcg8PbuqGaJbBE
KDst1islZ+GXnriBDGEnAQ/xYtOApE9uKl4UySnXCI7RL46gwV5gCB48xAjBcTm5Uem5bZp6FRrq
nev2qlJoXbHfvxlES1vogxWc0Lbto69/gStdajCvVMwGZZE81OzYEEkgu7OpMtOY2E0z6na8YCUI
49buPEZTG7f6gouTrNXMivUEn5GDqWSVdUaPw7KEajhRDE/USIQgOrgcPvPFowKvbpHRCLYmQIS3
27pej6E76zqZj8BLwvbt7+W3H/kcQX+h1aa7VfW7vWTo7H6epjJVG/GintCZGlgEBj/CUGHR5DnR
fargoOURM01+/T2Tq2moK8b+i6sz4/g/dCYurzcI8UJpDieARCqHd6K28jEMk71AwkY1GeVco1OT
vqqWdNtISFWeIuKdR2BTmF6Y+vg36efu2I9GRHAuKY8LGc1mbcVT4qzzTS/xyGadnOFyUKEJJ0n8
UoiGtL3ZwUiryzpiY/h7nyZGUzhbQTDDWDPbcl505Y1TTxnFLG3xbxnk+ndcKNPWikwCFbnAMyJI
NpNffueLY8DhUdG5xaHli8inYdQX7wKQLcC/GJzcBIrA4OK13gtGNTANLMcaProo0Qf4uL38bAN5
KIu7iROgTfs05hcnZVs3dlFgdDRj3bMljbZyZBlRSHWFTfl8dPatXfXa0Ze7pR7oRIoRGm8bJaHM
NED4jlmwuy/Jf08tG/MYJETnC8aU5XX5jAmsNUdfCP0Eog3z3971BKSZvOImyEm+Ba2XSxnIUpKS
S0uBbonins4CI5Jc9TqPZS90PdDT7J4ctPQVtWyHukT6Lu5AG+T0q2kI+xxFi60rb2YSDngwnlfo
5auJ4Sq5j3i3EiVHaaVAn++mWS859N/W8U3/fvYaafQ78b2crvlBFOVa59ApYt5NS7iTcgYEKpqt
VRtcYXRJeTXK94KlkPp+u6janXKWmMaGPkhnojuqYxCvmPoZFaLu7nwxi8t7FkI3oE7Y+XfmdJEO
kvTzSGXmEHimJ9VS/T99jjdxiZ0e4nP3TbQmVw4K2hMW+eVKkhIZyg+GHGCHDJm3/3Npd3BEVB+Z
fZF6EKB/lZ5lGVepwWWSACgwCjhV7D1mXEMxnM08cH/DYp5GhwxlmQ+Rqmh4BNFw+8od5BRkZ797
sjz0Thvxex4u+eSD8fZ8j6BRq10pcVhTXSMmRTFYHzDQ0sCYSvSQFxrEoICezKcuQa1J/BoSwzNx
KoFv3kbPp1NSFcKK5VLGwk7JSfwa4Hgtm//fRhfHlbRj6D8w0PU6Q+9xTWtEBxObUmTL6/K8fiOX
qFDGR/XoF7Oc2IfUQescCiF8DijhEtrZ180mY5qdDaJoUlNny4ASGcPRYoaKsCeciVrierLd2TWY
dbpVnu34O/+QgNsvMA3paah1iRRA6q2Cas+FyDE4FK3GUJyuy35bqwW4lItS+Nofunv70Jx2pPVG
cHiOcl/KNJhut9ppb+aXf4yxb1lb3SHZs4X98M08sMkCcqK0ga64NLMmKUN3BUIX7u46WElX8lI4
t3GXOuKLYg8NtQ977RhwmOsEjjAVgI2f1UEkOD/rr8hSSRS4RnZnWuAviFFA+15DtH+ifPbXi3lp
+aw5z1/rF35lPsj6d26FTPU3PLOxR6S9OYTukvwfrc4TvMKE/0d9vyYY5OBV+HXrd1/SnGwwau16
qatdOFyzW2MhvwwedfkK6ce994mNd3luo0vksXTMNUIA4GMHNJvq7sDfi44Kj/xIRqtZvvpo3B4Q
m9GzjAn6C25s9MfvVitY0yHWdGr8B9NH9HlN3xzaSYs91V3klXSzwNCTCpu3p1tBpru5b/Phm88o
AM7wS4UFGPSN3HMb1QZqYBw+u+1EIMEpICajP6uRmGFgQiihIeNCC6upaiTOdl/wpSaDmP3C+3ae
woJJRiddGBf1KLsesxnj1LFzebTgKW+hLuQ87g4KV3rL3zkzyptZduQbD9esGZL2Yn1OEBDeKG7H
4Jgkod3VeNgMGQwsA0FNDr+JPg91aerC73p9fy9uMMoOZhHPe8RlBgGMRRmZucz80u5+frYbs3co
QiZGEdh5WR1GuTNF5avhoduk4rmFrkwXblluCLquYxmqWFpYCwZ2wzxIghmOJtJkfWTpJlwnlK+3
9sgK6nApw110FlR1ZVzR4DLdFHWiAdz53nViZ9oQrnMPo0H/HDSvglBeklLJBi9JOmnKNoD1AcJQ
ZNHpS0T7vmHj2POs7aqOLI3F/EfCUw64VFPMvqzGzytT/tWQGpUzFTDmWRhDWG0FwPPdNu9cUZnx
nveBvYxH2Ul050yG1SsSSJiar17XU5CZRfZFuPBbdcemHsmZ5uFtMDmjeJumVSLyaNu1Nz9OyfHL
MRaykzyASSL3hhh2b22ofRAiOHW7exLSMsmnpcNrRSRPDujBpp9RppJ69a2UvFuxFr4i1OTD/Ezn
LplcKMPQMmzzi0N5UnTB0WVSUw1uD0Q/9yLSFUiDlSeImIhVonH2I8mATr3TJwY3uCtw98WoJ3Ix
yVRPID0G2EhrJp6f8B7l4QhMuKMmP/68rbkDbvj2IARE2PE/sIZrf9dXc2CsaFavRL7nqnc0i938
q00sCsFKsEh8m2UZZ3kNG+6jmQqbdk4aNms/RV4ZqtDTPWoCnMFvVCwGqJfGEk0fKXw+VmobvpDc
+DCgUg45zd8khGE5w3HgNFg225Ts2sb19jEZBHvc9Z6FSlgLJQw2h6KHvMr64ebrB1WhOKi14YF3
66D2sIRGylXtmw1R1aMUdRoGlnvUV3ngZWLm1JT0Y5D3xKilJ0l068m0XvDc790Bapt5YQGQXmD/
rmPtjKK/XSY0aq4i85KTYB+LYuEgFdCk1NwUTJZsgYCzVJ/TrJRgOyOhCfMb+8DEyKlvekVJM1e7
BDj/fUWuOJqCkLURIbJ9nfDVJ0/Pf/TATV7XVyl8vOWaWsHSTrPZ7rz21RairekjVFzsp9FGlcsr
IdWa9uoOIJVcdMYmASjmOrZWKc21Kn3huQSGaYLg9CDXaFZz0XLVexI3ODdhgilmRS84DVgy4TEW
+yGjQDcrxz3bg9msVpJwAqzQPzeS4K6lRH5w2ZBTFyRUqHkt/W3HcVs+2YiHm7HCJ6IuLRI2WcVu
/iIUJI7g+9OfONIWu/lO+7qMe8TXIRD/oHP017HpjxjLChI0AFigTE8POJwglyndetet92l4RmQ+
ugB+UZveZU3QC3jj4DjJ8DA4BfHyWqrMTGs/OI+LfUlr7cmAjk5EbT73Lxv+qI3EsEwWHZmXg5F5
hpJgSIdmYE2XvzYHJ3567XVyclOOqfzUyqgTTBaP7FhUNnbZbIoCmjnZAF4CKQiQ/D7cheKes5Ut
OvzRsg50ZmPH+dJ8KPIn1MzRyHhXYXCMOa1kR2UvjpSFXAa3CM6a4CvmPff2+0Pxjhy6sDxoQRIl
+wK4WbFFIby33pUpIGjD0M1sjqjwqGrJLuF04UMe7spI/3QzN0zvQkjQJLcz294oQTQRJc6fPzXb
jZQjQxEqjHb60nU35C9O5hWPT3zs0Bc1SWV2Sm6S5nvoTK6xzf3rHqpmn2kd0Y/1NBDlS1J/lY4V
TGecAjsG01cXFNTufqfuiUWh7aiCOozbaPnH8Ra18r09uOlb3E2gVt+r7kE2bB1cDZU1kcXEaUQv
No8bHgkNxiiWPnuwbDSZULYxPiTox6VU3fsgErzq+90Q8nCly4qDI7kUBTpw+O9n61xuMMoKvPNS
tdha2o+NBBYymEhlHpgYlzNydMial8VNlPgldlW6ACULygyhytZDKZL5XZu0DNEVGHzS2Cq0RKDw
yFeDxhJQg/KEofPWyN2eszjNJ7Qt0yhF9vafdEtrzYH3SBtKjUTeutWxr6n3qzHUJYe1faYaM3Aw
L5UyEsw6FTMqNSgmx08CW37JiWKrNhVozo/61WlVsPmbfAkK8kWKIXznPyX2QVMu5B/NOS/EmhLM
91fvs1wjBDlvwDUcGTagKzjOat6jCsgWPUH8b6Sd6N8OVXZvshEShjM2hP5VfD4uhm5HXQxF+BUL
f9ZtVhffca3z03mQ22f0dZGnCPNe/qEeZtlgj/tlGJny8v6TJl1kxI1ziXYyECa1dBFvJb122o/N
UQegPQPdPbhEPiGNI2xLRnjekS913B1uPdmNiEZldwzm74xYM+2YAAG1OQgsVIiSLtIx5LwbUrvw
5JoH2utCQiGSXWscmjrh2bTvC8dBT+TOOwI4R6r2tlGpT/SoTM25sAICLtzyw4S8S+0QQxmuhKMX
Cet0+gDixyFqErIlgCwrMDxmb/pSv24EVC2oiL9i3PrPu+7WdAby/iiqGdj/aQRxbQ3f2um130UG
TLhQdQsHykkbSMeezcH8F5qi3lncvTnMWlp96FjNg9HpBEf2JwgLTP3IyXsbLighIdPu5O6/vdBB
3K969G7ny504TQLLgaRskvrCryA+2Co4n8zHZbMp+gvMTvsHVtSV+oFjIQx5orf06WfU1LxzSOsT
HrUZGGOldJsbETeiL+XwQzuP/skpyd1mWT/89TfSUAPgYUo+BcBe/X/pAEtQ15Bvnhi2J+34tFgX
Y39/qCLqSLIAHt6CD8N5Hpzzul0WN725Daw2YxiwA185yTfrpmRWpRi7eTGPArQqfHdkNzqFxRF+
rPPkH6EM9dp7THcBz/s7rpL1xFLxs5nYHx7QdfsBGLO1rD7dKKrREex+s0lZrLgm7bgQua4lYYMV
q0HKMffIjNX5nEFLJCHFGILRoyZPAmIJBkYHDH5D2/e1hpjUxNZ4kjK6P2RHHNGG3BaqBKnoxc3+
09j17abOzjbJFBTjqbHW/LjHw25WaM3kh6Z2vLaWA0KF2uszbeCFz753cg+gn+Hy0ogqnFuHQQ1z
DdBQ0hd79QyrTCaV1qOdOeY9O8UbIUtCUKVJ0JQXmQF0Gzc5gBzHkh2kFwHp/GuzE1AaZS6WcG1/
UsiahI38uxtjpH0RtfcI3tlvjiaa2Yp13rDwWE6sv5ZHfxjRHqnakONBNNXAJeah97Vm7mpzQUB9
AHVrJ7APmammdMWOxa0/8qyv1ekPzTyzZ1nq/7IZWtKWoUjLHOkEBXEHyFH84bVBVsfc9Zr43CIU
zt+rck3j+eHZdHuy8aToREsnv29ynJtOWX3sMiSOMW3Fy2dL/+AtM0O3b1i3sjsdDgCFahIBdr4d
nQnkVPkDR7QDBGkCChSINRsKPcI8yCeZ8il8Sn/Qr7Mmt4EWsuYTBNRcWcr5ZxBgr1htDKZfS2aa
g12Z9R+FYOr8t3JWnIv9DRsak3C5v65clec5I8lEO1Ib5RsI6XLeZ0YMUIF3uV2AqZBjhQfD03we
J5KCoeZFKPsBJ62jpiF7yc9x3ylitzMUveAgpv5xPxSl5a3VftQRxF0Hteh4ufhKuPQ7eqKEWYeg
HELZ+e4LoKR3J/WxFmwll8XhwiKXGxhkZ16kmXTW1jO7cHwLv6smKi09DcaaDqNuh7uKU11FdBC9
HQQLxlM1gb49Y7kN+kZI5/C1BF+hsos0krut1kUHyVtx04Q+nfSg6vNtLLxI34wokEzHrk+ciTv+
011um8rBWjTxLyu8D65NCuXURhFwYZXtkkkWr20PS5GB+zQoaPL++A/yWsM7aAOVY5Pubdl64z19
Njt+CXyB1A0OnWbVZX4j8DUTV9BjR1IK/9NueJ0eOAI2YND1qXRXgAnIstScl9xcJ7BQBKK1CL87
xGm/aCeX64TvByxSgDe96ya/CbniHyLDrYkomd+BoyI6qISijoicAt82Fz5j3MOChdXCa/UzxA46
lMLvWfYIgj2HVfltj/s5AqnZxBucFBPvjWxYkXspYyzCXuQhDWzm28Tb9xflXPQKmtqVVfpYXlh1
D/afHETOmEtsqdPb45KeKn4ypxEdSlRYAFV3nY0CNcJFqkv9pf3TmCrm8kHt1y0yIQiH/56PuEK1
PxA1BU+q9SSn5OdHMEL97hH1LFcm3etSpy9dva4FuMA1bGuVZYBsmObwFJ0AXw/AYZcbgaQ1bwMx
Xr4NLTeCE0nAI7jUcF929eJOBIfkzf+sphLm3SXcPw0x5m18HdPpmQNpw0RrZxXxnGn7ls7hKM0l
FrIeU5HlZ5YkKYPgQNpOnAI09+XOJ+9loJwGK5XWhAd70tqBsGE+LDGNZWsrL4n5zfzviyBAVqBn
nsRtXC6QZEhDIGXVbj3rSn2iwIOH28GTZ9eWqQjMlDOspHbYtQOTdnXEImuI67QNOCHo6y2eArbN
LeuZxgtryZ3fTSOVET2d88nPxO5ZNd/bVRFoNh7X+Fz8wzrZBQy02dUuy8ldiVCbl35GopwRmW9g
kBzYm5Wn6DrL4Y2JLDQNZU7k8voW662WFGiuo0OGvqR1pH0Zorhek0F/lmyBvgvXeeADpnNDEs32
y4Xk0F11v8b44kTQJ5pTmr3wYEm8IzbEyGT9E3U2No9/iwN50NDX1qrzY4zuA3NymWxEEX5dlf9L
jJSwSTQv5NXjaBVtLcZnvaV265mOwouKfrgfPKYts3+VTyHBPbXTjDfJSuuSyRLSU2gBX4riNKEc
2vUB1gFA3QsWI45eK8ahLHP0q71gR+rCGrSSSTJnnEHO1A7a703YQpzWqWU5FJg9zWX+6poTGT83
ErtMh1FwPB6zPy/WC1DC2yiezuoSgZhdTBDLn6lUuBaw3u9eYx2urK5wkicOY2ygWFdARRoGHcAl
6IGoLCqiG0wfJBu5STDCwHi2pYxXSYuM9TmoM5x7+hLmqiiPZMta9FptKOSL3vHjDPUkbco7xI/o
IAf3+eQIgqN1pxOVHXmDqUa10wt9senbbgBiTXWCG+x2cXx6uNDmvUWgMg/QNDbOyO+3BuqJoZFW
Dis1az17S5P10FP13JUr5sue+CejFnCKPrAvM0/ujY82JfX8b/ckdwviWeFZvNo28o49VBMwVl3x
zSVM6GAe5zK6adwxqpiRo9Am87plQpw3+eqp+nTOQER0bmHL8LhYvxIS1yCHXY97fiyPjrHZDeAU
k3i1YIxgMeDbS4zYCJKEFx86EBAW9dhua1o78SMze0ebwdnpPfFvck9qm+2+GMh/0WtY3drkeOS3
Xzt8Sl1EAPr6Dtu5wIG4gWn0W0zeqQua85TCV/TaGceGHHo1qi5F9h48jU6uOZpMxjBAeYaAa5MM
fkLkbcyogCElJAprYpBKZct0aWtQos2BBGAiJIKBXrFPlc3ZH6jj+Ey7MjHx3RHDwwnM3mbbR8ni
CYQPLIeirXgda0f78wbvLXM2Q4Q7nsh5OoZgVT0TojooPA7SB4LeP2AuHaC0rY/ZGZ4E1SGAM3yl
Md9lES2lqL7dWyHvg8c5RWIfdItzuHaFJV07zyGjI6UDDIHNW0s000pyaV1r001pN1tZpM4xA6ug
+/JI682G9DTZmQOz6RcUV5mCRhJTxKVQ+uSaIdawrXu/Njo2PcpI81UgP2gKt6a6FKGRDoMksnfi
yIt3r8l9oaN0Jq7Ql53fIJOkoGt8hrJ2pq46IXznVyQ4jliGxUCj+QlARvzDGPSNv+Ebi6uyNrso
6qPH2GljhEROYjiNC0E/bLMclEUmet7UTZk5UrkneBjG1M35U1IhIJHvcF/orusJchVa1q/VNaW4
zxv0VSHXGiM3FPBXBXImKrEl5PaxVCR3evG3x6UvohEwh0/4G0P0lL4h9GWYZf1ghSzeKYIUU/QN
BCumyRbdKfRltzoHO+GLh+9ibX6c3N+wZfRSCN5Z//NUCZPjKjKtxkAeWz0bfaGc8Nq6UzXxtpke
HxWOBRI1gLBpHRtjzhpKMPg9+pf3zPe2MhRhGuY8gbMvk+Q4UQswlnjTRU7cNnQEGOMLv7TEBOiV
qvfhlh3zFY5pBerCp55jvXhuJMYfI1SbQCJpgQGU79QbhyNEQipshfwy4MpF+ZiB+n55AYbq2jeq
SF83lxHNZGyZSBUB5N4twlkxA6ipwwJBO5C4RvFtzTEPJ9LwAugWrj9tYnuemLBQISaxvmFXcHK3
PvGupN9PucCLkhOsKkAmIaWAIdlFWuwUVSueE5It3La8p7ClLvY3AJQQvs0uzn5doIUbGwHhdxsf
tKhcVlOniwQKbmv6e7adZMfT3Hud8VBv0p5bzyPe5oOGzBid+N8zBaBj6glvGXYKGRbJbLd41UF0
pbYyD3FzjVTHUtTe2bIbfCF+rqPbPp+fuYhGtkFDuZLnMtZw+wShv1N5/wyTjegJOA0CFL+yY2l5
OEsSIvMG3evzNQkmoGP+UmzqGz8GSbhp1l/8rqFChHvCi8gev+74rqiHsy1k5bFcGOWuf22L7Uqz
xCPyFPLgACslyhhrlurUvR6ccnUszTi4YY9zzySfOBAoyJRGaM30gSGEvv4wqNWpukL6ANYEEfxq
eR3uIC7Izp46JNr2pO5pl9yF7rMaMcDyZxH7tApeqaoAi4ik1rA4grXdRLY5VdvdaI8K1zDfnSWV
qRaWu+N1CkLcru2svVVO3tMhlUlobN+jL0dVop5jnK0vx5UPLdMKqw1/WWwY2hf6xKGN/GswNuj7
ECH54+UPr8SHNXHPjmkZmtMhVy0BNQs2lmO37e96zIc6F9wPXO20h6BghnH9YU/fdnjO1Ty0wFfu
BVZ6/9aUkrU7T0dAvCIGfzMnqYEnfFCZRO7iHfgZKUe37zyCgyUBMahb24sIYgrwsbBEUGI4Fivq
sEcjXG46yxPpoBh8X3amqg8C725emkf1W7O7BvPbp8nePCX6vcqdWSc6hJACtGJD9Cb50Pw3pryN
CNodHxsSsU9sBgw6JKgqdOi4Nzqyd4d+wJDiaZbF2UjHdSQXmK2a0GOPJzUqrSWIeZEGslN0Fsdq
XDVhzgdDrZqSR6vGd9YIKF8QTa9/mcHzcqV40hjpexHNfjZcb6yK8suRRSU5lJUry0Y71E+wndtG
SLp/ReoKo+zzneiKlALt4TTrQ3lKo8K8e+u45r7I4RBEBbhQuYMB3OB7XNwUMISvf41qlL56JMuW
xfSXfY2+RePQXhXTXy4gLqI7r2iUbameJVW3D96FjVz8o1eQlrCJPxN7i/oW6dPLPaftQTD3A3D/
mnOjqDwgmixAWDYirHo+ititXFz5uFHMimtjtLfQEBg/8/wAIEk1fz0gXjIDt3RRIj+L8VgMsySq
Sj6LwCaW5TUAXalcjEQu08Fhy0Pgv33uDMmTsfCDWbdh941a0non+tvNp5ggSJNuPZDDziiL+He5
vPDwILwo8QUjPMnzqn0u9EHQ+sPg7mAtw9gB0SK691Ew72gz4onYD14rrSfikXLjqYFNp/kYXsmO
JZE/HhJYnIXBeHyB3i7TTO68+4niq8j44Jk6w6P1+FBU6yrug8mWfe6xtjeWPkYEZ2zQ0M75nL/V
Of1QfKcE4TPN7Fu+RRHhaMsDrxSKzqYOE3PX9XqnHdszOGRVz9avQTl+zM73Jc7oCPhGck94bnan
Q8bcPY1rIw7dVuE7P2s+eb2FqsqouywnyI3C5ORNvwRQe/dROadakUeGL3/uPgkWj7/oYEThGeBI
ug5NK3gUP5DJwBejtLtdtiVbP964vUiQcUy77RYqJJrv4N9bJuV34iwgklOUwXpamadTzBc1smjA
OJ1vkfXfRHZhIzaKfNKWUU1y+6kMwVUKZHtP2Gg4a+snP+QhsprmwQg8SNqC6HeDXBFLQsqcMbNQ
OAOey0uiTSuF78sU13aYctC0lV1xhN/Tq74iHI1ID2sTQdrL6+iusFEBWCANZuJZEaC6gA4xvnzS
AF2X9BclEN4pUV+nNBAsBH5tntzLmjB6d83cImKyF94x7Jy7/9ETxHN9Q0uZV4QNbei1u8mY9Oft
nva+8i46e3Pks5JC+ZusAPoQhRTwVJrmS3S+D73z0ud01T4+fVArUGnoUlzShT38gDh7gQ1dsQZM
hzGTH7JlArlxb3hGnz6gfq2ND+g8jIeERQEcRoAf4Xl7QsFtCAdcJBAanIXpXrZ/m3vTxvyskG9N
N5mg7rIjMfFdNbYpqVJZDgsMRw7RRq+SQ0SkYSH1Pt+d7UmBz/IY/rfNNMdzkRfOycSLpUQLcSmZ
+fY3bUKt+2ookqV6L1o6oUjhMKqNwY6d8NPOCWGoHQyWQW/XeCGVx8vtzbtBrNuqESB7o9FKFTZk
JRdCBGT2aEnpRfrTY0fcDVud3LL4bEGJkmJJhiyDPg0NtVNfP8Gy4wY6NkYQgT74w9GMB1RK18yu
Q9xXF+pvzIK1/vDmPtVRQH9HpZqB4TFuyVhwjAfCwtcg0OmS1DCpiTnHnoTHtvwCgD1nC19+T3cj
ttCm/E+ae4CdFejfltA9CLfUQEcu2ttoCVDEt/CqHiZ0nqKzD1gxzwDMfYxMn6FaUmr22Zsy2x6l
hX3Y5mZuiZvP0fKUOguM5QdQU+Q03szHNOd0SO0cuAtTpN6KScSKHQNs0VQJfybSbMZvc/dvQVKA
H9+Hwz/x86aZ6L/HvRJDuzYr2D0OpP9aMx8DKh6gO4ql5oUZqHxCkJGx7r6wx7LSkqrUyrIeUrpG
eQLPAHGPAi7l1N/N6N7haLelAXftQuNFhg+tD7mkCI+wVmnHklhdi9NuCSTh0pdB7WuRfYiO87ws
N+1HaCCLfyvzX2fzaTdtCJWJ6xulRnTqTBFceKVm/VBsEVo8gK6zKcvStJUuhoWLAi+gG3N9bP60
9Y0z6Wbr/nsqQPgobn1lDGwR0XWc2g3VUkxJzF1HC8/fCJ165J9ukiqmMD7iCz+Pa72/ypS6EG+3
gDhzOvDIYs6SFhtCteGzQYcxwp1W56jfVuvtNdj+NzjLzEcFOKzh9GYQ2niFuwmtrgxArMn8xr/5
W//XUw3qsLKQ+xKsIFDePpQS3TPkJB/mmjeGST6Zccg84POvvFZz58ngJzRNluhIyFZHM45fkfjz
pdfy6kshasT3Bu2YveqDtP3VZY3m5LmOrNeTl27H23BnZWoxA+2a54xt9XDp4OlF3MYEuCvTVHSk
s91yqvmKpXYF3psaPOmisr6e8OPJ1nItYiOCdF+PMWaOs1L19BkcR7hTxeCZ6z7uUcfmo/lo12W3
8zj6q2yW1zJa8mc9oLF7Sn5U0/fm/jTQj1S9anUUb+wUqAKyCFRVEFAIkgHBBogEIdnox8WoD3Z1
PqKc45Np/ZnDje8G8FUqeox33dzmy4/RBoF4VLJzvFaIBDy7BwiO1gqoCxaUOSZpqO/K2A+fCTgD
S32O4vOC/A8RjUi2jFs3x/szl8lVXGuVlXNiPr9zQF02HJiaPPxnptAfJLa+jWblXJ14utB4u7Tw
sWXP4CzbAci3eAA/TutL281YKD/6Aol10EuhpAsUVTqPiXFinEcXle3CwwCXarJaX1LfQZmY8ZVz
3TDzheVQx6uKoxxXoYGM3V0eOPBL/aYsbjEkoqrHLwu4cWvhc5dNrhrjPVquJYg4rIDAzuY9tjjV
OPTJpnpxlWdZZ30PDTS5MTq6LhG98Fo9gpmdIdG6MRX62ww9pRY6ynurLIXr4ItsNP/Qs6CF4d4v
dAgTtkpynY5tI99NaGOi/zPVDabZBS1gMP62nyAwk6VRcMiJJeCjiMyjViff4i2Ol4Kxxx1+tYKQ
8UpPObrC0xOEScaf8ehau4aRclS6OKeoh0KzK07P+3ghI7lAsvwreVgeyaYclsa3hxoYotuJV+Bq
OFe74LA3qmMKBROwNwX7iIXRF/pvjgdorJn6xQb/HhQ+9fffGQZmMyXQsmTgcn9U5IffZPd5VbVa
h5uTQgybreIYgsM8M8GlQ+aD6jwwda3Zyr9qimUtZcXHtBICSFDMBCVgFa3n5CkYLo2bP9omZfxe
lGraTHQEgOktgJa2LZ3tep7z22uKkvHJ6NuJiAFO8EzPyOdn81sennFO8s+GBzvubg0+JwZf6gIN
E6WKrlDJoKF8RsFTVlLerRqQEGcU05NVM7aBKl47JtJVq9ZM37kCtytsTp/Y3iq40CGF1JxUjgJT
eFv1RPnIAvglIMxaAQYgFqaUg96blmQ0PkYDakJ0le2WWqmNFKJrPSfS8w7+rDba3nZHbGEWGKPX
FREMmARVzMvVxU0QXX06Z43eWCl9CssFJDZe9+8jgCrB6GYnmYQtPtgXyIw6rX4ASTYWAo4RfBIi
pxx4oYedfKe+JinI+ReaA7t3muIciRIleA44eozX1i3+pmbPs94tl3sIuqgUgSUErj0HehHWPYxf
hMiimk8KNBM/oe45W1SX/C2ms/MpGlIixJyfq1sI0Q9z0V530cY7kmyT9fn5beninfzsDAnz3+0S
zr2e86h/hmxxZ7/bh72dSp3IcTS+q/s197YrTkSMyKMlbB/OBJ8B30GnW/45RR20CD/PK/ALzyRB
OCNpWYP6VVtQiq3Vyaj3c4TruJ3iBrfnuCW/oHz7tLK+AyaY+T62dut0Wll4CI1zgMXrzAcfmSZn
z4m+ThpH8E7d2RwMpRFXHuw94IO46uVdcJm/H4z1luvmbM1EFUBWAhJE4NAO28lMOFCNCcqtPyLD
y6hgYA1ZmdZ89lnY7U0ZgnW/ZjnwYY5mDB66WX4I6WHxDm7xt04kwQoD6VEIYvOrWRX3lJU8clNJ
tLzXGKDH6m9vMcjcCEfxgzYLmU59gKSB5Mczk/2O3mWn/nhKqJj8ksmHow1EzeIfr0ZwZzglGCHA
WR0AZ0KvDTNjW3S8VrBOgiXBSjwKwul0HYreIx29+OEjBILfh2rAQlaE+su1qoqLFDXF+l2GXvRh
YeeuN86BCrrVHQNXX7JfZJVJk6fd0Z2EC5Vs9XOX9Eq0lg3ffu3Oizw+lZNXNT9ljNWEAZ80DDvS
aJCQ0QeIKFIZIHztEY2gBq3QRDfrBWW0z4lYjIMcFiI7Sa1t5URI8lAoCcMQ9Ax2txmsBdgJmJua
q6uGfbsQkSSR22ztzwMHeoS6jLbvy7qGFuhjWkaONW4J9kiNUgDOoDS4wNJKeW+fuL46+FPF+zq9
AuBKQUQeno1loBz30Un1IpcBbhJ9XxgoEa4kyrcgD617leRXMzlwGmvNpUzQncbJjPQk9wG8mclT
IiRyDX3fotIhS1x6qPKdujmOsyL0bnZbFutk6/fksed6qXnn5HTe5ef4bNaOWWYlaBJEw27DlW7O
HxAin64Mq+WBYnMHbh9wIAzzCTcbNm/N80e/vjRdQOBw2bcAwZKwx1o8z92nt3IGvc4thmN+2GnV
Ig599oGhbZ9aiyxymZROrEjopKTmzijeZaWMyZ3+VTIVLF0LkvdrAwnOmJM8RbgU5ArM6daR0d1d
yl85rRe+RnMBbWwhKqdphIxxe+un1B1stCZZU3mBdjHbro3ferwnOJYesfzwoXa35suGqMZESNKk
1BEP1YTmb3VR7ImTLrQ6MdOaYV20qQKVICXY2s8xDpA64bgK3yIcXIyIP71HREs/XGYUYND95hUs
lXphFTShSGeTd2K8kaD+e4CfLOh4DF1Xk6PxpzCJHL4RD5hdYH+2XQ4tJewBhlvIg5++g70AFa7u
2NyQO4gdVXceyKu0EKc1S6RupDo/HAyF7rgZGOPb3WAjUN9KyTWymaNJSFGTcIrwWm0bIYM6Y/2h
rxY5XKW9SUErdW+AQM5hlEZ0zDGpOwpJHbuQv8XYuX1p7uzSLD5eVApRY7rLlDBtRz1dZyzBDTEH
emhqfis2X1sdkiGWUsLRNdM4EIjbzmTpCKADaPCjbZ8GP3MKDVY2jVd2jtyOCMn9n+7OMVzcYWD7
sHhTjveq4qyn2+6snSjZqj+pne8/FwTEcohs4/Wtef8VzPW9vPiCiPcz43lzEjAS2RNg0LKnKsMm
u0sU1CTLa7Ouc/bto6z33i3OzZbJJkPWwuAvmP6DyuuEIeY3iQ7wpa5cexav2QvCoXH4AfK7am5L
GaG91XeYDPRNr5M/nw3KUsbF2Mj5tXHiqTQC5tjBJYW1nchZZJxD3qX11/0BgC9GIdZN1zC6iR1S
BYf5xOhJ+offDOexIyMxgj95eqrgC54ZqYrjsB30Bs/wFqRMqsrCnqk73gUfcyl+GMRifuKlZKp5
AHMet0hYpDS3tMHYotwwIHYzq8HYCzmyrB2STKJ6/Hl8hHR2G5Dph98LDo4QtDZ+rvbKPk+2bJ8Q
Y8rxY3si1PhaABNfEWvcLSRS6+CaEJGtQu+oorerLfBnr1gWGX6z+0xJ7e+s2EG75+EZ14fmzaAX
uhD3RDiE5/5l8udjdnP5yKyAVwxkQTlD10yKY+oTPF4f45AcdVzJXwUcm/JzGVOXUB9ecsy+9NBE
ZwuQbwrrwWTduk2ykxNUhRB7YUNZhq6UoINsRC7mcqi/zIH+9/cdn7wLAmt1NedR8INWzaYU2gpu
UVAXLUHYE8H6WT8PI5C6Vquawrafkd8iUacp/Y8GUwf353n3xQy55+DDcOpx2r/yCpVjXUopFnKx
tTyl33WrW6IqqxwCRVsV61lXADC/xeKpm3xRYqldxTPd2caij7+tNjEf1ASOnEMJdYQDXXusKbIg
OyLT1PNcb6KTa4sx50XjayT+UN+ZXJVOzxndjZdEfC7S6JL0qsUWe7CZu+qKof+rhwY3IcK5b2mI
i4cNTARG6/GAwYzfVLxFuWDz7UFBMFgNmgx4zdS8aOkBlAvlxls8Tc3nDpTHxrLCRziauxJSj1GW
qWCqXmYnoI2t6lp1DfEYVCPZXdkkY3Xd/OaDKlCwC6AQmKJH80muUUOpOTNXH12G7hDxR4na7JvU
V117Zfkhxom9MBkR4mH3WOukh+sVGxdnezBFfB5xhh7MIOrnC7LFEto9CgAl3MuaCpVm64Ff4kR1
T4XkVr1MzCMVV2zpcoUUrCnhMX0RgfoYFtdje/WBVMBAbIvWVjrxms9hOb5ai0Nh0DDqs0h4dHg6
BTjnwMqJ6Hr4JLxOO86FbiW11NFWkQGCQ4B+CE7HHnO6Js1L/nxlgPe3CElpyEofdnOIyrtHoj3m
OlqDsyIZbP6tDP/Mk/jaLlUlwwdoKBmHOTVkbEaiBObtpsd3Znm/yZnblgFOEljaH11nR/u3yeQI
NggceMy109WORSduKorLWTX2VhiKJgm86j1u/1y2sikjFm1J4LYbEKrGXdVeBnCr5PnLlpT9jCO9
ZbPDCqJLrpg445ExD5fX9BHe6fyix9M5Q53RIHtxpt4x21K2vE92MqduCV0u0+EFbJ1JDTN3DUGy
NB4cC5V2VlW4iUaYXUhVab7rsWLeIqyqtAD7Gh2FtjpWo7y6NbfxS8j7+nEhMdUT/XODxVdztPzP
0R5V0lXQcdBYGjyWN9fHZMyRnqgyt847sygJISDrNVkmOXL/Eup3QMKPr72A/iGuNu41znbk/864
VSY66j8T5+Wl6f/hXCTPGyNjN29rCb/EKKehht1NqAowUMW9R80bUAw1J3VLWclK/5h/SvN65zNj
AqN+2XUs67eWOcS1rkwt+z42FqFKvdOii6Rst+QWwpPS3bI6bZ7B7SYasM/HqQQVcdXsg63ZFskv
lH/x//xr9chAcXVR61Aza2Cb7ASP1ExmP2XjWnV31bbx9bOvr+uaYvr060cJvZrCJ1dt1H5wOjeK
XBdcmMHgcgPEKOTiZ2f8GaVWPxcUeQ9hnlRFT9m2VFdHWVM20eSCCNOHvU2bryBsELrQ57Wah6ub
R50XEy56cc4LgH5Xd4acAQsA3sId++oYRUDrVn6vc6KgdABDSfZmvae/DKFdHg35XRbggDRLSBOd
GxnWnjByGCsjY4A8EuR4fxeUhdm+LLe87pqvaY3DmvIgTmLYKcKlI6E8lhTZQGf4XDMTv8x8UUTm
+UwYDVVw4EPmMSf5kX+l2nyHQ1Iepkj5xmABl2rCr6JdV1svTbv7iB6cJ4+IEwi+B1Y0FsSq20Ss
SI/8ZXn8l98bX+8Kwv7d5y++d15u81a2hCSqtBH3VBtQAYCmHhfJpOkG0FiouIVzote0FUrag7kQ
1SuDS1uWgECuwrWMB9zJ7kSRmzp/G3DNmy2BtvN5AJWja/VZe54d6l3ticDU2BzX2X7ZQ08bPN4V
us0lIdTP4pfZ9zAUccch2ki1ZDvCkUY3xM9pItk9KE38wPESGci5+FgODAsSggXcdEjVfkk6uiu5
D9VPl/ED0wCAavKMwRpfqw4JVXyfaw6RvMVAQ/W/n1X0CDpAoGbWA1Pr0XDCf8ytVLcN2hroPiGT
OV5RXaFq9eoiLQblRpDzSTgHGCjvmKvuVgZcQhz6PTuYN1rGjEn87sSrqvMWzCay8aoIJboW/rko
y3HME3DJBsoAjHIGCn1+mYg8Rr87hfrXmG5e+fUBmuZYJrL+Lsr9jY6JxsesDh9WMvv/R1uHPAAC
YUKLngqh5MGYlJy39iN7divge/a7xlU2l8qtrACjv+CtJ9n/qhNrpPTeFGAQnSTxzmazDZnvkVzb
0RNdov4XQPB4/oRGaYoGET7sMy8SciVgKUBj/zlBab6AVbCmyj9dExf0Gwkm/YxlxtLCLdThAb6C
dIz170ntI5FXF3XQuCyoXNNT1J/UM6UqhIHE7EDeTs+EDH4o6bchxHO99ldY7bw/SpZiNG0n1OKF
727fZd9JcaEfJ3mCoxvE9LooXTbIcTm3L8L3vJxndOPRphABLgWCaF71H4P64zoagMTbVXU9UA94
UuBEbUv6NjxrRXgMJgnEirj2nNOmNbD1mgH3XWW4E88e7I7LfRjYRBomAlll+3kwDE0xHRJrkt4M
EsUf/xCdXN7yRko0ttzoef68GqIkIM2YRNuszOcEGGMLHs7c9a4YS1FfVkiVKtmkGqHYEgA3mrip
oy6q4WvHHc37bEoCw943WNKuQ7SDE3eb9Lu6OToQr+OyNw3yKXI/F7cw9iVbf7icyMXNddMB/eKr
kGmxvdvqr+rGViDAjYkOyHH5RK8Be0d35LrS2sGYkqRF4hXKvbJ13FS6XOCGIjMaKrZjeJy8kqi/
jkG68zGho5TCcPMfY2KZCmz4lH3Z8mPqnJ3b/wfn/F7nLCL6gLRjMTYWgOWWXy1amLTWn7jN66Of
YzXp1YK0gCkzysNBrgrCOExPMF3MQtp9G69eU40vC5XPMoOUcu+eKcQSV1BD/QLTINpcgbUyns0D
2pcLfVCZt68CJvG2cYlEKXKOZPYrFyS/90uWpOPPh4yT3cR2Mpv8Nlay2sIU1V4LM7Uu65P3/HOe
87xS59fI/yU0WzveNAJS/bpHdOl3UCRvjQ27ModwfuCfQ1B6q2oG61j9Dd8LfY295FegilgksOkf
+mK8juf+3tAVk3Y/rZXq6ig5YF61iY9+GYRiFklZgjYzuzdzqrVxLNFAkZFSFozOmFVVOb1UP97v
1xQLImA360jtALKt1urdwfiuIQUx17oYsp0WU/ZYJx4hyrBWS58+YBNcxaS3NFYoTg667ZIUiOCo
sKhfw0D/1BtNSBI6DfxOUJs8G5PsJ8gmcDiC+lES4iFQfNvF8k+LqqxDHTimzMTEPRYKDWwpQBYj
WVMjEGc0K4zTtgAP2YFc01B6LYcJw3+9Axo4kP7c9EpQN5s4g7uuqfH9kj7dlIxTb7IEFNH+Ism5
N1aUBY8tSH/8h8lEMUyzTHAA3NVH0CPeNT53GE3BVlNhk67DWRCvc93s13ahGzFYcQUXVFehv2u/
TjwzfQg8xfpnNrFJhmfG0GRXRZt+t14bOe2/qk6iIHdAquNycsBCMwfKRgjfmfbqoAbzaSZNqfw7
1f0ce73Ji68FFtRARlKJmHnBRCeLVkOGpkiI/PraVPxu7L8hvAE5GSwJAffDc9yR4PITz3ECC/Ks
rC1in7VXwg3MLuI0fpcv84rho1SYLypLcfuQ15BHsf2fKg+4efknLY8ePxGzEVjs8Mvs4XWghpfm
cAQ/sefKj56V69mAsbj0TrnUDtINkRvaor4uP8WS98IwX6bjOjh0n0AcgxlZ45VMXnKjY+YrtOS6
4i01V/enbOju6Dbizr6bECC/sE8Kh9e9XO9UCfNh+mM0qTKz44XtKMBE1i5xGUx4os17+vmku65A
0T8ImcAb268yMqi0g7oCYMOue1R7vvrGUC1XMKxJJP7zwugMz2A81DNCZzxcp5r+EcvAjOu91O2o
WlE957+58TudlRAiYiRS/1wr3OGPU44VHs4zfqAwwpHZNPLte/iVF0Gu7xMandeLtFRXMvXkYdAO
NbdI77Ki1dFHjexEu1KpOjqRWq5H7bsxcYqjuBOHr/m7ncqM3DayYUInQ/WW7Cg0rCT6tmnzuExx
DcTs3HSGloFXCx8im+riVCcjoIA0zlEQgrHDT181qseZkQWPbwhLF4eQ8mahP7fY1Jz9NBOBM3Q+
7j3lBijgPOFU62EYw2UL1HvH96sbuLBTAWS2Loo92gUyZg3jn260q6I3Dj7KJs0ADhSeQHVSTN5l
Cc/HqphZcmMzu3vjohYFEygUtdZiyX9Ww8ezVT03nx66UaRfEGEW+hhGzUxeYyz7H6ez1uGeOvmJ
n9XSuCPr2DXCCPaHEhxu72EF/lm5PONAdhcmjT+LCMpD9fQysTMoDO7WRtj+DNQvpyfWxyXp79N7
4BtLBe8cn/fBelGxsS2n752MlIFDaOBEfj/ObSf0YQmuk1cbhHeRDYZWD7bN7GoXxcQu2mu9SSqE
xI0ry8z9E4N5D6AB6pANJaHriuk5F8Gv9ySvIfybtC7tvpzV5WVqFINIx9EgKECTXyKIc2/WlqAC
yUZJo+aqjeJjXYpEBGHQm8LLZJCPUwHa7dA983CGl6r1aDGGhWIbDr4vDdaFyzokh4SB+XeQmFh2
tDzGydYGLGXGxwaY/5I/G/QxclrXxO7hlfxloZr1d5iBpKXGWMyxyFxrMAhJ5E56Stg3GI8enhU2
QkGGgQGeX8hBCe1emUj2y3PYrWSDaqUuWV2sg+RnyWS5h11AP/V6KEtCajqONxYCeqOLuuGgYasx
Zj+jFGNcq991tPhgS3i688Q6h06+1qw05Ncy62mhoRcEE3lL6PbUciz46txoQu1zx2LgG0rfKhXW
3luUAq5fBTI+ysS6bpFSulICdwqg2sySbkcTWskvc2U2PS/TqiUTfnsT27fs3s7dKqZJId3mtMRY
uPAH+O/76+1k20sux/XBSTnJGWlsFHSxcIV9PRfOiwi4Q/7L3PjRSG0A/lIKvFqr8cCEcyxpqLXc
nLW1mGaNHwL8+HTTiPlaM+dpGO4X2fWbgay4ulypML2K0Qz5u42ughiRVUbSViCKluHDPrylqg0a
7v9J2kN5cvC5O1BX3s40n0DXxDF3zL3xZ/avfNjExxgqzJKB/Fg9mX5iK6k3uqYptP1rkUiMB1bw
gJ13+PI3052KCCqx6RuEPQrOBX0jK7e5u3sMeZ3HKITNppKHOfsQbMgOnzVqG3mC7GzHh4N9/hmi
aPwEUB1RHGpccA3Cl549CVFN8D3n23eH+ANmpIVSF9ymd86DxRpF3RNo+NIifSA4ZNSKzisYjKTD
Ad8AawKVv+6ruXJuafQ6GFqEr0V4zdBVktLMLOBljcCyzOIeFVsD7cc18uPpZj4i9rXUmnHtiObD
Q41Sd7gHfbrouJmFuujIycG8qR3RspRI6lh0vOzTGkV/y+075q2NI8icyEKYWLqzr1ovgqxtF6vm
KWcmeUEPt3/kiGDc+eWFU1SRfRpSklC8henR9N1StYQtA2QsDnQc3eu3qF9xaSWJRx/8VL0n4R4/
FWXnDSG2zXw/3/2eA0qfbBDsYZ4kky3PqCT7QuhZ6CdGfn0+dZll4Ydjvw/66fd5F480JnIbN3sO
g9gul8qqrL03lrQHfxh5WbXOjk4p+aCXBH4iESJhcViGw2nagfnzENnE7OuVqhk/kuWIKa0Ue4cE
YzrFbvyZ2DvWmgpe0GpqM6EPmC/eUjHtlTkZb0se7dElnId0I5to3ieplGlq/y/4thGy4zOLqAxP
OQohvyEhtFbQ3Y2gS8+bIpGeDf18hwmewQK2TrLxRfx4EICDcA4mYiY/4/3So4XM5P2OzZTXco55
ztQuuRbFARClBuPVhE0pGV4SjAVRPjT03m7awyPrpzBLQXo1yu4NQ9ucaUcDEGD6YZsivqGLtK0K
iHTaFCIZPJ0j7hMS/rmFaJMQhBWbqdAyWYCDlQL2wcEHnQ+waVf6HZruiGjUixZxTOzr8/RAa/sI
SlHhOPvG4FWc6wZnxWhRmc1Y9OopCGcnqtiUxvm2ZW9V0AhxPLlxzX4ItUPoJGnl4A+tz4Aw0kcE
kYdiIxMdJTM7VlaKj0BBPrgcnUKpag37FCQEhy9d/P2hUwmClQUx5Ad4jYUzffD4PQIvM1Hmh8ZH
uWnmZRJs3zSfksLNnFPFT6s1ZQrpAviqj4BFpHQNw6yOPafsxiuhywIaStjYuAkbDNRwqrOqRdwh
nA3RtdnzgrCMJ+0QpF+aA7GMfzJ8sisMVt0PcM7cCBzC0LylHDMIJIJ2AH0JPMI7ZNTLgL9P8n5z
4p9LEve/DHQSGoErmFepwpTv3TolQsxrZwNQxuUa/BdbIaVIei2oZlpqL78yH2f4nUa0k2PGQwa7
0o5DoOU4hTsDmcNC528mK/j34GA4mV9v51jQ6nxiWYT+vZptPB1YUeKkxoUAIzRjg1Z7a2Q4Ss7p
FwOwBEXUT/OsEDjYjFs/vuZMdHDJg/+ieK+jdFxr7+gEIoJyZLZ060VsQGEQ47rSdO9ETd1A/NYg
CPgmPRvrqGkba30pvL/sWaQ96G0H9/bHXIJEVlqs0fYpR8Sy1/eBD1Cd9KgZ5qh6z2l+XBOc7/A6
6c92LhGaxbh3fdkRvutnvp5m4L7YF6pf+4a11C/GGt4tDOcufvTWQ4CZLbiBdn5jy39aiclu5SfS
TuX3Os6GOggz40blgCIdWYSG8PUzj7tbs1YPEgJ9H/qln9RoeKOYyrMC/VXDsz6wGT6P8eJ0l1nz
7B8b2e3JR4xxAtuFjMb4RPFAnkzxhc9IAbZXZJp9XOCzMVW8YtWnGoI/O4oBdd67Mihlo7SzHiJn
3u0wOQX4ngohkCMnwdzY96oQuofk+LhkVO8MagOjkN0phXAeXwjNEcVT52x94as9itQWRfzBTGLk
lRRFgOhr77osbhrNBHE7xyj2l4DnsNtv0ch5CLo2uxYTeZ+hGc7WEgHXczXLtvxLfFNVh13COMUl
t6C5FIQs0qMlgfUa16hikh4GBimj/0Ubj4ZVRGErezIzwZUPSkIPi1NqJAxAeazEcPS2fhqRGHzI
k7Cwt99FJEX0Idhhr/o5yLUUpMNySIJGfy9GcX1SeSkN4+8g1TrfIVHbgVSIn1zr8P0d6JSFbcPQ
LZ+DfLOqa5RnLXtYCfMtp0D8tN8hPGZ9xbk85zBW0Kb2t2jthQ8mo7HwOOuSPd47ypj27N/tXvJ2
niEMoChkqxuRh4OFVro9a7g93b/mTOa/bl5jGxQaMTRd6Wi44OgBeUMYLPzHrY0zXZeBikfsVTjx
yJECAo+cBAuWIcYLvSsZ0o5wehYt6GDIY7iJ38YbF/+kEJXSU2qJbTY++Bsi26AVtfTdTaC2kdNN
1U/6983vaBQgir6PJMJXYEtSKZWFoigWCrXWMqfE6TgjEo3n9X8zrmajIxjkb577jNizvSIn3GDo
ziB9Ya2JS4ODZ1VavJLMhlG5vE6gkMCYL8HqwiEAiLLLWZvdCrISjWMtsxCr6VSEQhxHs2T5nxba
g5JafkZgJ/XrNS2nMQc84fJGNlFcWsC1J69ubn/zKJrHUE7/U82xbqsvuraYRnTgvxSAIIv0a7yq
jt2VHw/4R6VAdj4Ew4bsXRew8R6O71bfymOzeo7Urk1wju02rJefKaYbVqmCmxhsYL6n2FQl2UEM
Oyh9xvdnQHXozLCt7KiIrXCL7N5a0iILXOM9b74rfZDA+61nfqKJShUuJXHtDoMuNr1P+T4s38dU
m6w1As99j+QmvE5i1TEePC6FZMPeG1dPUmdMw7YEMAewXCctwRpOM8GjvlJoRcfU8tBCCcf9JFX4
nwDFx91RAiFDjgWmYDrkPUS2Si70bp13NI41JQshh3w3dYO0QlM1bFlSR6z63yEzfmZDjlOs4bHi
KHMl6cxyUcQTWKkU+QYKC/261SX5dX4kDJ6jddGOWHEi3Tc4Cjy4Yi3gWXOTplCCiM4TOqqGbAf/
fGt+Ct9tOMlUjrgbmPKxhGk77aF73LbTMqeD+046UCEmzIb0nXOaZnD0eeqYotQs1Xg1VPspg2Pr
uHsrmI/lZm2RA6OVrrBWyZ629itT0rENav2GyVxR6fn+nrqcuEQZJARE/uSj7sEkLRFDukJUwxuG
JNd41JHDT/K/0+qJKG/YDXTjZMMPAA5pj5RHdhm7KC4ddNGERaqBii1URDrHMFDZTL0fo5WsbyNz
YY80JEFft0sKnH906iWYbBCfaHTrMaudIFgNE+FBc3zzAqMtItAlak61aE7R7+GB0xF3WKgr3O1P
veN0zmBQSa8sADYJnG3LMd+yDQ2RnHlLdrlHC5ehWklWpOwbFmpadJhs5PsfVv4sK57ucpeG2xjV
Ks5NA4oa5ypvk5G3+Cfg3PIsA4PV936DNhnjmJsrn4iAs41j+nvEo1+B8Auv8UeiVgibp/lextTu
ctU3EKTJVfWEdr+IugNgW5T7/Np38vDY/rSJPQu9Un21Wg28f3AiIYx1XJdpcv2llmGK+huFq+u4
PJ44Aau31W4Khd0LdWpl0La4akc5kthT/oYVhpwWcJWEImrFU4LGySW2ZaiyP3q2mAgfm0PPa1RD
KIg1L3FAFnV+8pojSCUoA5jqwamipMviQdsHzNJw9wRseLkVxKXVw3y5L2hy+/TYZWNKefSL7Ls/
FjjwqNySF1ISMQGkZO6C90T4SdkZNF3x/Lj5BcxflcxU9zx9mc6M4oFHrpPZr8OaqT/94ww4ejjp
eUYLzCzxopdT6i7Y+VFxdLnsULeDD2dSZaKN4Dnmye3OeMxrvgdfDrYVCx50SIWFn+Qw/W8RA/Cr
NwrxLJ3R7uyMfxWVadn2UKJhohC27m2K9R2b9sG+pBpxzaAjoYdCq1jVS3wQOWaqZjphnCadDR5D
otPcOhEgfasGC1T/tbcWjahooxntzOtBMmt5p6lW8MEy2MMetCPjt7irvavEb4fVW5SHxQHLt/hB
js0oKqm4R4a5aV5rvFihPEqGrEdDFLgg1joixaCukPmuC+vTtwhZGizhAoqjQaWd/EQFqZH/RBaH
j4x5VF1NxlB3zpqOZkNdG92qSUH+le6lVgNf65WpCabuUWR2NoXAXwRyZPd8uKfh2EP6xkBapvFv
b66Bgz0oGpJLXMwuKBEcmhm8lge/fynqGqdA6B30RE1njnnM9K/h/HJFfSmg7yDeJ8vJ5Zt1nvMO
5tfoQEAHSbpBqnTHbzd6Zy256HGoDiRYYQf53wqWEPMLS2a6ESv4rXXzZP5RXLRVLtYKeeE+59hr
3GWoS8VaAcb/6ofangJV/GBnZ9gM8UipUmopcWCwRzF/jamTMNW+0AAAf86+zc2tIm1WBKFUC+5S
NIUC33iDTx2kID7VP/0/ZK+Q8yTNVdpJZjVWWniMv5SaxuVkJrvnCVnMGZeNyzICAONGiqdaFX6j
e+1g+fuEJDbIjvvBWh1luEc25rhNls4jdPZMfm6QzeBWn5E29FUdZ8p1SJKrwrzSmoHJZ639E9XZ
D4L6S0Ffhkb1OXk3y1WLGDttYk6wlrSuhMRFEMsSg0aYkVC6CsQSGn4Di26VcvJueUWx+LISPzxd
gYcNIYbhhI5xGLmZHzEqhUoETQiSuy6z/9YriaztrryAuYcKeaIzKV4sB7Wwpp3z4z91r8U1p4oK
ynoIM4qPPi4tGfV3LxHSM4qcYCOw89OHB+ERSfDW3gYCvZQRQnuf7xq7NiFyrboMX5id2wZYm0C6
VMyyF2QNFPI8/wQsn6o9fRow6/l/TiJYIQAtSlptRIcU8cwd85yANEuGHTZWsFGvXxU5rzMeeCmX
UGmEE/mvh4KJ6yGXfji4rTdhHsAv/cg8djark8w6LEpFF9tNaWv0XXRzlb90iiNLEGo6rTZYfbhM
1eaAygcoNUVY9VKzaX1aJuNo3zpy4HevrQ0L76Dvo5eFik+bW6meDLL9AsCGNw6KnReqL8xzoU9o
n6TYwTVWrEHsNZOPfGAWlCOtjdNbZAfex7kipt+IFTsRpXXyqC37izJIng9mkQ9CiRls8thSmYgz
vqNUDSYM5LQAKyHk4EvdiqW5XyCwuiG3XOpTdip2s9gmlJmeVs7+3wJu9NE6iDiy4Q44GQZIWrk6
0N0NKf+5qvhRu+EcDt63P/KX/Ubx0y8K3gwBHeBRo2cMrKiI86W6Xq0gbfvAXy/EvtZqE1s9OAIi
0d2+Ywe0cX4g7B02T2voaglqn5JDQjMMd9YqXpCmdh52mMBCF+cdt3V5uYEYjTLHXTWiC8UCmgLa
1N+8gkiJQI1vM8h0p1jG/8hFopHd2Qzg0w+IsqWIsjdOFdn1rTfoy4Du7YZjH9iVoO5gFdAjFo/M
2GGn6aV26TUzQz4XwFfLTDjKHQY7geX1wn//Mc5PpPiYV2ZcDLTBbinndy0mlTAVP6QLKmHIPLCX
iYKitInspbhKULguD0dUF3qFUbnPctU0Y37x8O1NAeIbCpIfBgeyHnp3wJiXVPBaEe6wfbIArwT9
lRUMsQxFkriWZzjWVHc9geoFmnxBzbA6VYpvbmj1c/nnQDblWx1OQHq6/gb/Isakzk4HkVjv1AAB
W0EdtfmA6PNypdLbQtbphmNFB91mCiRjr8nzLnHFc3hPKlAE0Ipo3S+5DKzibwjem97xjrTpyJzg
ka3OFdSLP/F2plzq34dzTdKOkyMYFbXDTKzAjwBdq1KH4ELYCJH6qdNZZLahYfywSbpEMU4p3Uc6
EiND6+gtmumQ5BOFE5bwBg00piOZCa7c0zIeUWPHxIYwG3dthInCzyZTIfcSpdLZXOemSQt6E/Og
6mtlQwFHP2Ummty7IGMCCqIMW7iRXVswDmjDrweDJb2i9o4bXo/fnKcTeIiR3HY6XBV7G2of574c
sxMq9j/bc8KyNhvaWqiX0Vr2+JHaWgJRtM9CYGSnBw7RoSd/PVP1K2YZH58s8XEWnKLwWA/conAi
p/2BuBGoD6Pc0I/tevosYW0dITGRpFAJXiSYiQ0GtqTp13lTMLG8qYKMSR5b9lHWBzqHjjTEwBkl
CGLY28GySIeoujF/J2jpJij0RJeWiK10qNeofHRg3jn/Fmq6OjRAnpxVJ9pohYe7fxHtqV5h+l3v
KaDb7/KFgMKYd4dKnmlgwQ3fgmshgq1U37Tn8u+6FFe7VA3IvE7TY8JYJFdWruImbPhaF62KV+s4
TY8pA17xJChvjv821RKBv7MNd5AG3IGtiYJRQ0ctnKcpY36bUaD9uJSkTJIzaKoSuRy7VJF6iIfc
NZ1K2hYEF3vO+jV2XIAvr5RJmpCtLXj3rAAo6V3kYrEPYuT6wOzErbqr6M2GhXmllWxVXoFkGI+k
geps5G7eybE4u+N/X7XQ/V4xQD0AOBPFjT5wMXY46Ww6m3sWXqilAwiuh6XRjctQseXoCutlS/ur
tM/rHvBKCQtNT9nJj22LZ8H2kjE+De4x1dag5KmT7jUzpK+ua8rg/bIK//DN74lPh47gCEo3UxOr
Cd8hvHD+oddACrCl1/GcHN09iRRRBTasPtZRxY9Bd1+aRJHj27eu8QTZ/pNVMT6uk23OBwt9CrCs
XzNaVDF+SEna0HswnBwLcTKAPafTi7m7kEBEqP5XBeKbH7BmpaHe//9vw1ETgf6w/bgQ6ZRhlxrq
pP+nhQg68qgIMb/kgvUOFO5TljCbGc5W24JJetdMpv4ns/HuFUp64T8tFrV3mUWywgt9YNA8ovCL
D5QbgVujkWPH5nWQhzm5J7PcxA7pubi/E5FyfvmitMamQR6LD4cobfYyt25KpplNi1C1WXPMaHZH
y77fvJAkLKLrK6NaGcw/ov5UoZ0jIyKouTGNijywgbF8iMa9v8CVe2hnJ5l0oiGD5GSmT1FQ1B5F
XfGs6xiEwQAed8xkCGm8Vui0RKglvXz1uHqa+X2OgKEtPNuJ7ICohPEdpZDeLQw6R7DIlTXwrOfq
5/Quba/aj6Fvd74t31iSCrj+NowtF/QkYNuoXmbCr1BHkPsyseQ/F6YsCK9z2OH+l9aLrudeKonY
ECYcbIUojWW4KJ5tV0TZ801UbfRWxipsyHhrYLVOJttsTksxWHomkNhYi8o+Czc9wGtxmzXQ3Y/d
lxaxiyoFyyZw5cGmqZEkhwciqc2pMN26tyP+M9YWeNTEdq5A5FTpMlrsBeUcNmqpo2CI7gMbRJDs
2S2xGqKqMcSDkQ16NYEsUgOQfiwf2qXstT+9Y5ruGb/zAKNeClj7Nl9JSe5KQEEQ4NR6ycSkPjs0
7mxpeEoOc4HUN2caSg6h5pPYrC/mlIDW9rl6d8h2G7pkak9GeMli7Yed5/2bORfyMc9m5PjyIajA
CxoRUaidhXLfuMLuxKCeJzgv95+3V53755dOWeK3DuuVVrMaA49hg9cvSOD6ZDeunJ1S30g8c7R5
ClQH3C3sSFbs1jigonHkI+BhLf5CTFAQpskIMU5SbzsaT14SGeKjYkPmgKjX07SPKjFLKe43VxLQ
staEhAcwkvDxMJ67GpFKMLgSmpO5YsZ5wc/B3mrLmAi/FQbLMYxBT6LnTq5U7NgimqLJxhrp8xVx
kJWcAU4n4UVIKVchyxP61F96hb+8fXXa5FXRDHlaD4QCTC/8LnTC7lqFlk+khP2J5U/lZfFrgfs3
hMDmAXovo5WrTX2w6iXjQbH0gD8HhJ5K25hVH7YEfR7NfJlJoijaHZn/2PkqRqq8ECbBHCX+0mNM
XIWQONAVdE0gSP/tcJDNM7zbFaZXfQq0jMOUCzRKqU9GyThSGgTUdvmT6nc7xHEnM0KAzlu3mtEA
QP+q9HyRxQvSrai6wlM+qVumW/LJ7Wmt+yH8k0DoooEgCOi7sqdHYW6+g5ewG9vm8a+V75OeL6KB
15dwK7uZsfxfWeES0CNJeOMwxHPTCcIoHvDB1XUapZ668i/9PhdcRW+a2w3j9xaDMX0Q/j2FZH1i
2M4q+uGf2j/5FlER7OeNhmg3g17xg8MmbqrZ3ET0GxyHn7UMtLzQf6/16hZqHoWo7Kgo7OaUxcq5
EwEPakJECoSpJo+lL67Q3WwM8Qd62h7UVXqj0rB8ZmnR7+I6EglQz2Im4N9PBeeI5UkkDctlOvTp
4OozrDykHPZd/OFU3rOjKHBMWG9ZDtH18aVksqsaNLqAV6Zs+Vc196OUwV9ttUleu86/URbag8WP
CyfM0X8PUDNt/b3ctJrGP9T1DybbTZiEAn2MYMts1kV/EaL1n0vSNA9iG9ZJIrp4kFqPIhnQJTvG
UCmqkPAPAN1etMuXvQnovhbfYpk3YRfYT8/pGuFwJ3x7hzYPkv/zz5am0nPScwjXB+6eh7l06kO5
oS6JMFHhjfHAeMEnuvPp0bD4SG94x2jKfK9GX+JmcGimwiceJ2hWiHwAXL4UxNjTTKJwOnIODqC5
Q99sz/QV/DjACiCb/kkixY+VTCICW/IT+y1q15LOMO5F1aXrTA2b2nEcR0ffIPOI4l5D9i3NsxCn
+EyCxXw2ZxgvwuYNFuHauaMJKn0caXds6zHe/kTWWmefjPWPrzYIWzrnd53TP8Si1XXJISxa8ZQq
xf+h7YIve3hGLlj/WY6IY2kxGKnbHBg1KgVViyq5xv6OCfkJpLq/tBvJN9JE/rLL5N4Zp353hdby
OtH8hWc76bbbh9a0Jn2jj43zb6b/k0QwbaiK3Mj1rS22MmUxpWzO0NXgx1j+NiX3W1+/2KGjOf/v
H+uqIH0UDF27x2aeSqD3RF6PvG4rceMqUJGQboMPvCh37Dc30S3vx8k7RP0TIJSsey2eloD+EEfc
wrTGNCW/0KfUC1mU7RfQhIkgkeEUM1cjJAajMkN7NNaazYz9vZ+2Ogln/qDdFn5+e61uGfnkWeD7
fogDeNImm417tY+gTWUpcyhq/JVSPXq30unpAPW5gbVnUxnBt0rLV/HGU7W9Gsj35T5if3OxAyDy
qhcOjhlZa+xU2IIS9Fj/Y9XiDpmFeYzx+fdCJIZ8TciTCKbAN4H03i88xhiGVues60l3//vwYkGO
i1eupjR6hLbvXpkIGb56qV/jxExid/h95zMYgxHmxI1qhhwObXSR5DXtArzrBRRfhHVl0SE3yB+f
XfleaW1SKwLX/AAjiXgI3kdkgEiXLhelfWtH2yNOEOzuW1b0bAfHiY3gr1DSCro+mut1fRwI5CVk
NEZjhWPreQ3hBim2Q3iziPrZIWFERvKBTuXNC7zJExSz0wjwyhisjixk1UQTggf4W6E8yxkJ/gGJ
mTTehftFSKd6/CqL3rrGAMiibEPADIv1doRaKsmFpJ4EJAoYqsumrnqXL+wrSrXtcKyOpMk6IAph
UqA48DSCNoMFmmdLrrDX4+B3Fzep2EAR5Dy+PJu5EQ5H6RZ9RlHdxdNocmFkedzCU9Z0ZxrQsIoS
9xrbqPYZoEUCxH+jUzP1uqK0eBXXJneCdakR3trnPghvmiIiKKOWjkqoQeH50mh1kXiZ4iBks6FP
rLYwImk+98raNPfaGnBuhNjRwn8WsYGUgFBDS06jCCwp0IpP3uq66LRIF4DNBI97apNOGopZknul
uxjIBBkkdN3DHEHEmGyEgBdz/belvZAZN0paEJ+YUOqCds3zu+jozInS1KJeLVAzRztne2Ed7aKI
VNXeg99jveMVIBeegkJJbTQ5TcChwpwu4pe28zz/xvc6yztXEL6EpRbNRh6RM6BaQ8wMhJAbL+OP
hM8rnYzRfk1uZwVTnc2IEBydOlHm/0ICI+HS18Qu2SOZ8Y9Pk/OWfIuLOjG0RA4avxHnndM+AAJ1
fdc7CUfAxVeq+4fQ+XuXKxR+i7kfFUqixQurMsM59r0hKc0SA2ZnuITBNhKadZLu2MxwIagAGj2y
RJJ/oKyg1QMB5AGyqftEpFwkg2LhmdB66lUazvy/464PcTJpC8dJBUIPWA+kMAMFJA/gzwW/y34Q
011qylQHoTJKwrl7bfntCT39Q/HWa+k7I6APuvUPlp2eC0bpXBwXAClxFf4DmXkFhaCmmYLI/L+C
ezH+hnj2EvPbRinROKm5wBrmdac6WJbENsoOOOdiTdtQxyiFh1AhPRCGr718G13a01Z6v+P/fSRN
CLX4/Cxwi+LaFXbZBCSYjbix4L+GsBQNp3Yh9FuN9ESxh/3W5QOr79qni0gwC82u/3Rkie5ELBtc
kYtlBNvsUKeZv53edlkhlZsht/a0dglavX80Hia901usVU95kR3MuWinlqlJ0AxMbpDM0IGSo0FN
X9hdQBWIM8/OXs4SXUQw42oZcAyKpXDt434NouqTpCQhLLIC3EU0ji1D1J061zDSOzSHEsOM0oUg
23w9UbJAjEG+632rR75FiXqBPbHr0lZWSMPzEewFqenyXamLxRBJ5cWG2dxpfHrKXs40W0QkX7Or
+6ylByjyuW08LJyhZk487oeE9lQEVabm1dG28uIYLiD4H0c2bPmMVrs6KFmu3bwWPOWnsZKiHHkf
YeElJAO8YRi+ZUz1Dwzy8Q1fkgAVMiHBPPWfnLNqTw6YrZn8XfambBKJ1iwUfMfIlncblAbTREPS
ViMHcAn8ggrYgbnDQdNfjPpMd8h7kvZXC8e/DuiubevoWQauBodvkJlTjsc+SUnFzoyIzTO0RIty
E3cH34y9jZfktW9zhjWvOBWKsT9Zuzuv+M1XVoxLe41EAiVgolK0tjEkUGEl1uXRbWJJx0Ik3tjV
lm4PHFjoThqn4ncULxkGCFtn4RUKTydBuNcmpODXfKoyp5CnTGbbiv5stYo2wUAOS0ZWuU9UgXd/
60LZqkJI1zZiaAdZ5Ur2PpukBLS8q6lGBwThFFw8tzjLAIL8/O1bdNZs1kgWS2cgEKYtr922Os9o
/VfU/5juLFlIGwaZClOgVDJkuhruFMAUuidErutrO0qKoiWCGOqdcYzLpl952VIfReapYkd8jo2q
2RLLjPv9axdD4tunHiZiSEoa03BnXQKWyhVbAAv2oSZSoOEUMWi7frf1VhpTBRHBWMcADFsa+XSI
32PVTK49BHNndne/oGvSq/vr/HZxcXQmfIdotXicy0HjHgHoTnaB7Q1pckOA9TAJpO3GWPlgoZWF
rmupbn8L407kAf8lmJ22TnkDRaoL0SYjQNyCklIeaQVTmC84Gtnj2vUQLyjEXKKi+oTOifHZvHQA
4iBHCy5KgDQhgT4l2cRfmdQAFw20i/5RIaSVwI4yKARGMi3fcwx1eqVP9aPx1M0KMV3MQ/nf+u2P
gsFDPyZU/JRrWV4McUbAKz0fBuFCw8kH7I/lVyRX8LIdE58vyJkd2qc7DYXp6xpfkNb/zOtE2nNf
1wbByqVARxgudDxiIvMhI3j5dtZzmFqxQJWiJvmfbmG+mQwGQ1i1it47fc11Dujlq+Tib9Zl9FQD
7N79qqPV3pOWNmt5CIoOXX6K9tcRabh2zcEyHFBbiiSptFPSuucMnFEELdbfS/kmHE6eGJHld6/z
LTwGgmpMbRsodrz2CoDcjgvcvQV9bx1Ha1bVBzhCL/yShMUjLA+EysZqDcpyDsknpAcGUuVhZ49J
1BlxEwErMiNZ4+P9/h8LslP4VcOV8wlBG7Rf8C8Zkit8LGoyJ8XF1jJjgGI+ZAZ1FAxB3+cvO+QN
WfFiBYqQftVakvdBcmO3gGRPIqcES/0sMHWFaZKvizpQtYNcZf7o7G/IyuxcTVN9tJmGPUZmzPJA
srhGxRJqr+OvDHnNC+F0zjIUgsRAhHjiiZRfeJAQx5kZdOxUeurYOHRcQCJqdB0aKLCDondSoGkT
e1Z6+yHYW76NFU4ug5v9tcAptrQWdyU+k4uvo8EPcBHmbdBpPTNwG/4tQG3Iv+X6w8bKP+n50c0i
4fpOj6DeTV7cBpMw+XNv+/Qwz1jjizLgNnthSSDyA786JakS9vQQxeqFJsxZ1Ah2Sb1R3UyISFb7
h75rf8oic+Ftm8abOnEWxt2c4C114GcW3jz2t27sokbKcqa/xtMiIJAa0J6X73T8r5uJMVdVpT1T
XO97ezw+wqmEh7oOvfsjH6LVpaIZj89N/HDTNmGnyXLwqwn9soib5RgIXASgHN47dwXc75ocpfOh
15mOeqce4uasnmt9Noulyb765UYY8/Zds3XoX3Ts6TI7C/Um42O4I+8XvkSmooh1abnW1rAccJKl
3KreVu1gF5frOd1b2HATeMkmMqVjLVZhlpl3EBvQ/hiB4KIbNLiB7Ee9wHuTuy120PVoSiX7/BFE
7Dgx3VwzDpXy/ulV7wA5YGk3BVgQ9zwy/w8gvbteEp/qElHvMblYFvEyemr9pedhrtDJRhj8wYD5
fe2IuSSGTs8b6q5HAsDQLlsivSBypOl5hpFrYjYqmj685QX9iU3BTAaUTu0W90k0RlkJHFSBXXY6
aIaSL/pFwwFyQIsTXF7PFT7xXBwLeBCVgKvH1SqEDRz0NWk4CQ3/LHPtxJBwgwMxrF8OV8605WQs
Qe1xMHhD8r3+hWvly9ki42z4hAwzPMEYfP6Sje5CIg/34Wr511KjEDLrRPi1O0xaZBxFeqEptgEw
8DhqpXj2SMMREA/lkX/V4NgiHEYUVc18PZCF7yb5lJFKv0HyTvTnxouwM0BSErKNdJN1yNf7S09P
yf8DZZxiKPObCdNApdSwdDRJTu0D2SVsc/bLiH1C2+t7boSVQrq2WjIcjjRqoktJS6bgOhZ3PD88
+8Gr9ac2+SzxPgVvFA1BOhu/Mp2S4nFJ3Ji8Up207fzh7RxT6LmxiEPIDee/Jtlu6Cqayt7HbDj6
BtCbBDe1CNudseYbeDWcvyA348e4i0vfczcnAf4REBrHwgyGJc3nB9LUtQgoDQ19/qYs045Dk/rv
DQx/fBSc8QrfwSlFNGlgpdUV9horE192l1izQ/6cI2mz5S03aYndwdv+yH0WxaaEvVOSiwA/JJLy
AMLwuUltqmvgxVgzrwF+5JTLEY22NeBkf5GDxGwj5cusDXHRvsyetvC5JIBRDHUsFe4tn79GjVmi
VuQZf5ljNQDwBDhGWXV4sCua7QExqgtfIxayyZfUzKSTBVrDrPRQonjnZe2KwCZan79WOeNZ19G8
Yg0rW4M3jMrzKZEbhsUvMiVWna8DYZhrppShnNEE+E2wVff2xZDrHU8xPiQqHv2vc7Y+hI6mzGmN
DuwDjbWefRdnjgUMKjTDOX7IQ4OG3tnMFhiMH4IBPcS/l56M4bihYC92aMkc9ysYKfjoAZeDnAEl
d2Urg7DEZY6LDp3dZSZNWr01JHHQLZkuCO2+4ob74sZpReuZOTtp6cgv/t6C3xbkrdN78cJk21zd
s3KM/Dvnjadl7m5YtF3lrUyKqNNTfzvnI12EbO83ViBapoi3xXlqgvD7xIF2s4BbBcJ6wtgw/bu6
qBM1wLz2VRSHgQc2VvcixIgWlkeyFYi0SU7+bESRDlNKa0+areL8nIZAjYwCu4SNRjrTMTwA0Riy
yGL8uurnTO3W+vHsud1LGnUDI2ySciA43k4YVuxPKihsC7puKPrsu+y1xDs4Gx8OEEJAX1nyZPiI
bVBSHUQMqV7QHhZhhNjIeO8a4WPJjpSRHSI8HXIys/dRMsd6yFwCiZct9B4J1FqXsevv7Dfq/W64
01N19/5ZWQddVrJjqO6G5vpyjPu1+o8P0+qILyiR0wot8nmFjqjQ55BLx5bOcelB6wylCU1HBlir
JekQQbO5702geuryTjZi0vYD7jZHzO1FHjgX08dhrmkt+PetUAPhduXor451GArWIbjnCg84/5ZO
fGS0RTlHh2W+A042lmOSsnhdYufCWXdjhPY+tdOPGUNIklG81x5ZELfjdfErLTEwPiIfQJiWD1ZX
pYAp09R9L/ARky89ok5kamelZXhpi4+XJ7vKPBvenQ4fg8tOtc1GApOY7R6/hQQByeRYJvMvBqZI
FZsrY+0PEPp0zA65otP9gxl5wDZe31uNnWglitAPPSXzssXC9Q9nACOd56OJ6BmKtIgg5rq0hT4S
oKWxVemq5YhOjoSnMSAQIYvKZq4T6556pf11CqMW13yTSHxdMHlM0um8hHQGEtI7tdwapXkT12Hz
TVT5P7PfoQUlCWTXUFJJEhFJ5Kyh/koZVjhI+zKOuShvWFbluJFiEaDX2sByeIBI+YvbOaCzBwUP
ca3y1k5ZXh6j0BWlLoDJGWoAaYc4NJTxy+GnmyAjjy2a4Im2znRTU0XV7z5mH+H1awaz7wKpXb46
TvwamZ6DarugxlkOSBFfbaR+ubilbPN9jwS7F2CTSNpmhx0X4FIQ4QZYBPbC9BbjhAG0nF3D+bIh
2UilgnV1xTRGtw/SfWRDJdKl/sXEansk+TpuVJgpt+1SmqKTEG8SblHRWg9INWY45skcOxRmqEIv
snIxOeyJ23RlpffKmZVbnCU37dzB+SkYmLHmA1BlhE4NdWTtyXt4f0IEahXMDoEjZp8laRhkwPqZ
8EdXEooSFaZY/iCqMcLYNwFc8aAh04VC7Q92BxzSGuScnHdMxDKb+UtB1sTLyyCeNybHwt79UefH
cQdxy6Dn4j3Sb1qpE2EJCJ0J8zgyrWpZjByvpxW+nmEDoHDGUeJSm0Hgd0g/MtRquaUVjFOGaEs6
n0z0io77WvquUEWA48W+zwjvVvHOXDITrENydGoouZ3H5052XlP7hWdOvt7sEpm27daj80YgS8/B
gDRA1QvdOKW0CPpZslaQlPkGt9nYIlOvn/fZXyTJJ2ch2C4DaeLzre2V4eQolg2xosU/QbCJ5vgW
hINNl4lQw46lA/glrANaWFzi19OfumhGqGCJkzUqcXWsi/abK7TF0WR1GBjRVP1j1vgK+yvsKo5z
yHorzLLxr2n9IJj312Sv2ePpvH8I5SbQZsKf1xqxZdZrSEKORhyz6zYb2vjDlvvUbqBNIZKCvliK
JqUdNRj9dDTxkwphmI/+QVw9RUIUIPoRyacKbagt2apuH2StBFvphuerp0TX43MnOqePoWdCAvZS
nwbdfPurtTYg9AkN7wz579GxojV6goS4ZN835GY7mFjKpP5y10JYpL/2v8D6eSaVBtRuGm1g8zSy
fktiDC0eGR8aiHkoVe8NF+WHwrhdKXp5o9SV67Bfw2zrFMvbu06UHhQ5d0W1oC8UbDC/+62Bu5Tz
H9qneZQ1L9qt7lVLnie+yfXQpib2LqTTK4OyL/ttjkdC0CRWQN5X7KISgJC/oT4F3D3zOqygAxMQ
qiO/EOZ+xCZdcc4iJo1Tawy9HHN/TXZXA6yxXZ7o+v8WaVX3nHKbu4VyZYllVfL/aBQSBp1oJJ7w
AK6SzUE8RerQKLgCccX9H0fVFUknEZNsyu+jy94Vq/MndOgmJFNvjcLee1VSfxeIw71/hj1QTKlj
9eorr0I/iGzycDJMEHkUog/4TnNPfr3jsUc2N9+wn/Ls+DeRpXLzNl+oPZu+t0QxAYFHXdpQ7YyX
FXmzJ+MZZRcZjuD6YDbvQYQCJIs5o3GF7CShBtXxc19YP/TAUMsU0ju2Osr7FAzyf1VT6t+zdFUD
LiNbxr/tZJZkNMNcxiafN9c3FZzDHOYzlvcnxbM2Vq8xZrJPAjc9UpvjDxlvLn0KDM2POm6bN9cj
/Rx2gz5PB598jwtVCU5n0ShgsvM8bCg4kAmXZJirDbkb+O4cJ1WJe8jhD9HjQWqHtZ21ZrHjgM9y
x5L+SyFz3x0DbXhRV8ols/f+p5jHpQ+lMfGR8uQ6quPsv6OH3x1dytW8isIPTqtmdMrJR9A9dKeT
yIKTMGRxGut0XuiDnhVy8ETyENeczgxgL1ka9qQUwrU1chBGAmE6yeQXNvCJKUkjQn1DhBeREG/m
6g7aDmXP6uZNMHm9AYjqygvfjWW0Z8e07PlM9REuZDw84K5aAqWBLGRZ3q1cOz8SuUscFSY/OeDi
z/ytuEnoQhlvqzVWMG88W2uH5dhu63vb/VTmuHjCTge95q8fTLI7J4Bnv2ngrXl8ihurzmeq85eP
tvPFYNjqs8LkFoFUg2MMPdphFme2sxIaFD7SfK64nQgVtlXuP0Ocg8u9z7S2XoHNjH/6Aod7GMv3
C/Ynw5sj6jpIlaG0wVqUShItpZjTgS+AkM5IR1qIy1E5oX2BvXfmQzcvab2PQ8kC+Y9qMBlgp7Eo
ZuZwkWDI1eUogIbzsTuvdM/celFoyt4+BMP3GNB2qxUDWQkNCeuPf0xa5aBjGAIpCse1DaDrf6jX
ujvOACqf1UO7xRNKjwOAEmZ0qYpUDT2f51iTH+RJdEq7YHUvSabLm3KNTKeHOlIRwlzrZ4VYlKMp
f8eB1WcWpiRbFGahlm9lMgHbrYoNz/6BPt2jITk2kuzaBB6vISaQFiZllmYy6YGSgLkW70S/Xdc7
/smcwyaTFto3s+HtY5cQB8K5umOCF8ileWmoL1DKp+0H92hrNmp9HVbx6Cydh0HTBHhxoGFIcP1p
ON1V5gwUKSfkiAiYausPx/pDUe6qiqQwtGOW0nUovpiGzPHxQlyFD2xREKRLjOETrEpmANm2u4nU
XWg9x7nayx+R/4x3trGNLuAAUmUcBQSNY+fuLNgWnws4BMfw3m+TOxCwCnk7m9dzuZ+Bsh/z6eaS
/amfzLsSH6AukqrEG+SOfsAiKC2v7B1GNJgZCcuCxEfJLnGDjhFXTIfN66Z4vJTiGLFJI5NkQ5n1
WcK8Z+AFRadW6UTQmvHSSfUutRgU4hlAhaXYijVoARlBJCXwIzpOcsEE/lpifqftRzTSZ3EWseEB
nLNncBQQdZGM9J0OIVxyhAVRJ4RXiQNpvqTQLLmU0757gP9Gm7d92Al6hxKIdlznrq7EFu3Jytcp
g0/EP1foF+JAtob8UfsjRViBrvtthDWSGJtt9Mvec9es2lzE5IdXki8shTUR8q+OAbrZ3nlT+484
TFe0QV2e3TKP4G/I85nFnaFV4tCvzIfEJgDZEK3o/5u13cbNNYzlO5tpGkulv7EqfA/NYjHYrl62
WjENBOkPK35yHzdrwhY3VcJ6D/ouCw0silbxyUDQtT2J/GpNWM12eELHWPa9gt4wAjJyADl1Tlk2
SyhN5bJlUsLz1nDNYRqZjW46XGaOdEiqcsCKYLrKvJTxz3xeXl47FB1kdWB0cNXXFzaMvEycD/Eu
CPOUMPCx3Zo8fvWRfxYUXYMTTS7Y/XAug5wPD8qWd9UCzP6p59N70Vtw1wEz3YoxLWsmudP1wa1h
R5kGvAUfp88waUgZL+vBYx/dZB+vHpitY0owEDN5vIEUFnbN1fsg6scMNoinySrRYboobLGHi0vo
HQLtTn8gapOKEW7A3VewmPbl7LICy/a7zLNJoFp+aMSAg/Kb2amf+S56YfyDiFx+ApZWbDLFnS+E
W+4J1nkgRUSFsK2tMacRnx0k0VuJapbJO8WS/OwgvIEimV+GnmNDWsECHAljx0ygqNw0pp/Ro6PS
rj9e8Fur6ivBQHp4bHzaWvPerh4aDlpzxxNuavdZrKQBd6bZ60V1tAqU1Z4KVLVhVeZIk4gowEeR
KO3ZnXV7rlGSBrlVXvTGBIaDT+i8TOIZ5C8XubY+VG07AH0NGVZOQem+t+/Ow+DO4OhOlyz08TdA
PP/zdpaELn2vJ3xGfZTIhO6uizYPQsnXC6+c3g/Dbpe/liu0BZayh22m6pUI83tIaaxsqbfbO3Ns
2nN3WR3Zn7g0UfbCe9In05A3VWuHsC2pADiiyG8YTIT+wXt21ta8vovWMoTT0D2gE5GIdip54d27
JBVfQ0JK/dXHfgkfBjqJdF5w9Gg66JBKvIL6tstmVeHUw6U5iIf/7EvvVwpeHiRm4PmfXrFY5pLG
S9oyHNaF7IPC7qbRcKxa8H7+sRj0ADb8uiH6ola16HD3euTnM08/pz7XJ4BkQBXd00tK04hDbW6d
JCQcb9dFCYTOF0mGO3cri/kf4tCyVYuwhEgEFJqBbhD4/FKjEcKmBCm3N9wfwBqIJr9pF9tWFwWR
kVDWF5v6fSAWQylC8+fH/e5l4ZmvDf/UPR7TgPnvymJw7I4X299sgb4lOYtruSAXQekVs1oPkAoj
NmDS2wnfPCTZtKTxGLtrdmeOOhtjVjIxX/IWNYy0s1vlUaHPN2GmjIsWP6k/lCfksaTaiwS77W1C
i7f1RyICfSiZX5tEg3PkPE6k6buBBYi67qBVPHMGiJvHZM0KwFvjZ6bSxxWcE45ZUf4xQF5kh7UU
ZYnpERsMZk4ejNsEmgUCg+1sn5F+V9WrPD1+BAb+ODvVAVUuiFnh5ASA+KL/6L2563oygYNIRIa9
vdjHyV9ixDij/ww/zb5lPwas5HuIrg16dO1nA8NvJtkldErSOmFM2mStkR1i+vsArlgTmA8OuU1W
J3l+hkFoEXdd2O99p8z5/b83Y1A1PqxHCcwOX/zOQaHp7wFgW1o2uv/c3K3JdVTQW2fN0eRPPUgg
GeSAMoB+zLkwH0VdvHXvY97mpFFrWFNhYxoczpJZRK/DWCaGBQhpkxCwT061jj+mCWEL1VDxD3RM
i+D3viHMs/M4AkKhZMeCpqK8BQ8srtZydoswVY5gSKYvQDhOOQXUURsznM1UY2sbX4BSnsO8NaD0
m3tMK3H7rdxAigPFMEiBGq9rILb3c6CN7cNnFcHZ3/bqOH8pVkQz1/i+3zBAlRfcRc8/XCf0r9My
EIIrU4J0By+qBrE8IDyS79P6V4IZK+L1XIG0zo754J2hf0hNDoUuZkkIJlOAbAOlKK8k6j4IGp4i
MzP0ho5FCw7CWbjcHXG4zFWCxgY/h+Sr7I1WfwySqGRbC5GACyZusQZT5UPZcYDGCQZDWdJrBWQJ
kBtUAJur5NaNZvjlbTLGhcOcwwuY/1ti3f55rFnKVZMAqSUZ4qYPrFEXhJXCkct7k2cFWBpRxG0E
usqcwyq8tV8S1GtlRJ+NTHmfc6kFqHZnSRGL7QKJlbOXMSRhVWdmoC8Jwoi1uWEB0OoOeOmglksN
++k8A09va7mll7Oq4l5kQoix+3yv+YYL4FLduLYXAAE8zzqWhzqnOexfyOVVZMgAaMesEAzRa0Ab
DiShFrteYZ0qY7kisaZDH2fZpFfH7SeIabPjfx5HcQKyL3U4znL00gUk7Ki4vz/YVRVQbwNH0XPl
TeIKhRZArOCdAjfJeyxC7Iu5N4+s8/RKbG+4nF8sIcbXKgQKKsQt1TAzXubg2fVYqrsv9XlYnZu/
V0si0XAEPDRa7pOcJoujE0tPjo0iKEyh86hkr9jqPgozZKavny+TYe4HyZjLygusPlOfUZog/ucR
cJnJBOIs+Lawk/BrLBgaMjJSvRT7WHmdGmuf494pVdUp1pkbGL2NNYf+9yMjkivqbSsUN4kebLtI
87RaZ2jUjTSalLYFxQRmgnobhLcdXzUzYro9cdL6dkeE5xCU2bWZhHmTulg8Wtan9P0wwmErzSHG
18EB9oDKhOhw9w1jW1EkTQ/6pyEh7uGc49lEiqwE7LYYAV5juAbIgjCUnnMWsKKH6pqysanuEYU3
YqtkLOkS1A9VRoYVaCtmi25T9tEW5/jdj+os6SMwdPsEzMPtPYsVeiNsLLfZUEyiVXTvCo10HEIO
uX+UzFB/Uf9AZyyevM+KAMCgetSM7TR6MGuiSHU/R7vaqxmo1uY1M6y2mF6YXNiNqw0ON3HqlL3c
uv8oyX3m/H/EZRiL2o0GXnhWztI+UkGZHHN/IwK4k08l1pB8a0DEo1BOKk5mA9uSYH7z+VDtVANl
Wn1xKrlVAWIADTKObtmZ0xXC615ACc5trOh2yRR52dvtKi8jhNX6jwNtURfDEoAbFvFbK2cN56l3
lEOElqJDhcB8mVskQ9UQYL92/MEzR56fikP0E3fXPqG4fKvyzuhxyEaCU7hCHHXW8kvlMqbS6mDw
pk/0iAs5/YdChLX3MVV8QSPILP9Te+1ETpS0HDjRL5pYLW9RJ41HFvSHLwsxOI467U2ZIF3dSLZK
yPxTHnGYsszPK0D+cdussChtz0t8fMUmA7aepuxK4XquDMKDjSkQqY0bHTpS0mA56Jifq8ZtMknN
K9sI+GKffiepD9L2W5kZleii/OXROjZRTAK1ifVanvFJpC21oXO0Kg3d/y9d1wBrm2Ff+KtBz/Ed
vSYcnKcUex5qZ/bYkvGqwozDNmCf5rZRwtYWib5A2RDIITrXuBHG9ImcorlQtiXb8n0aUgrvPEQj
IucA/tAgRUc2G5T5H/oZE9RicvywRTSDRSi5x8Anq2K9z7hMl0OLDQg2QWzecG8jjAtDnu52Xugs
0lBOz6pJIRodljco5Q0wzVa0mmrQdKOSi6bri3lLTPfsSJXsweVg0rxyim9PZF6KghiFwFTQc4IB
3Mmo5a8rezNA9A5lmaBF42UARcaRxHm98dYu1rSiAHWjePgDkpK9scj2wyVdVlGSu1+1OCXJQGxj
Y6MhW70iIeg4F2+GMf/btOoNknEDT/jTTr4+scpteucoUS5qUk1SpMPIgBw9D3Nr77sytczbpxUX
XJg1XJDaTXVdf3y4iDk+Rsa4Pw48mfJpwiUvxzJf57sVM0lfRphTwmkcF2rxbMborHPXcZ/b3kNP
ZfIldQc6IOy4oyCgFKjaAkC8XcOxf49doH6Iw2fqE4V4HxbxRP+n3i3Xodt64Sh034dHXt99EfnJ
DD7X5YnLEQWeMt50+nSLHM4QZ4HSniIZ8STSwRWrPkhemu6kjPPBU9Gw0UBNgyPYYpYdQCsNm2y8
Rz/vSnA+FxOXUqrDtdasCjyolrgmUF2wWlD2JLfgPgHRCzwhZVvJa+0SME9xBURdsx/TvQR168Rc
tTMdoDjEPnTRaEnKGrc8f/rk+dfpQnmmvANmiJtcRT3Im3K+4eKIkRy+/xdGBQCDY2R0K3zh6Fak
R+F1vP4vhH6CGas6UEC6mmibegpUs1PM3RXBC38G0eS0jlrTKeWSYpQIF9XNdeh/G5BZvV7OuFtW
Sx5BXWd1TLGyBxVEmmkPyehJMb2XIglcsUZ8e5XA281u+PEn6sMoI79W0Xaj3T9vumD8qUEi8c69
iSnRHmNTaU+UDB4vPJVguzOtETcTQ7KdJ31U4RumtSP1u0E6USUgNTGBMti5gUaW+9AsUZtOW/ZL
nS7Jo7RGD0R5uFgqdRP78jscU53bdSfe7Pa46LXXiWHfUyRbyrwNVqoMo/dc3aO+0G4PJPUVjHRk
T3XqNrwdzswoB1vSFAJshLwtp92wrFCH80Q/m1mI8DXOc5QVWtS1aEb4ARf4qZ3/JKE39y597IcJ
FAalS6eRipXyf5pXYd9iMVn0ZYyDwuIjq+sK+/1nLGFeqBMwoquhFhh4A6EchUXN+2f1m4+l9a+F
DtBUvy0Zfd5rwyape37QnOMAS7aZjJf/j8Kc2rlpfI6LC1LJbSpcQzpW4lSbefa8hIL/VfI0EOuH
6mDpt+pmhlZolDWOeXx9tagihmiVsAZPQFCR9+J2vxT1ZKK0o63nGkzDDZEvW7ASxigqJw/SystI
NvgWK4rFWWmcqXs4fMKcxCxyT259+n4n36zhity9dtKCkvWoUiR7EsbQ2i4Gqvd5zow0h2Gcd+A/
lJo3Hn5Fbvzh1T/g9jOIABmVSc0RcUFVE+q5EgE8XjzvqnqQ2lmxlAHI+F143xyXmXV1vRr8yh4Y
g880FvrUQso0TbEVBaiHe5qfy8IsS0Ruh9MJh1nrmnVLQNWbzFBh9N8vXdjrPcQMCOD6fkR801SB
sd8REvu+0cZFtjGcHj34/D1eqXOTUIy7mW1SRX6a+kqfs7ojVGX7Ncgr1Ob55FZh9xzs+8m8+Caq
yuV8M/LnLkv9EXjzbiYLFLKsWed4oJReo0jEyRFVBF0R9UYpjMaKHA3VYaC/hbi34BA1DTK0rvBb
howPYL20KUEE4Zsa9St0H88FvR3JpUY4KqegfUr84qAKx1L+ZPx+mQY2lsQb/03ol372uTha3JzP
KDHxWgB5KVCVm+b85W2H/sCtiqM8oDO0cI14x3T6YT4V41wqC8HZArD30LbEk6301oTtAiPqTEOt
FwZZZ9VOd4/EZ57HP1wyhU7tffznXtxheXFZFdREiWmt0LJzdRC+jdv/SVj4HUvJJIaALTyXY6e3
kPMx9zuckP8EVnlM6xLGRlaLW7GavjlgrK1WW99D3UcyVfyoi5dc83ioOWZsNio9NM5Phim/zPUo
7f1Dn7VeKA5DkmALIwNC5cE5FJckAnBj0w6/9oCt4pAx2A73xrLJtYBQXiPfBuu6Iln/H0QkCDvS
KfD20iSbAeO/BrKYnqTGTeXEB/cYgi0XlA69l0S+U7uh6QHXARngEdIklSuhl6CvaFKUe37AlpR8
9XRtV31KtDIeOFF/pDmiZgeBUI0ArThw689+uXRCYbWuNKZyxO4g1aCqEGBLAVTaTL7/gSH6UU/R
gdsJGY7CX+1STf6xnFXpdHffMI+s9uuXSVf2CYaCO6WSl9SyvvwTL7z/VxJb7oTEwGMyEFv9z3sg
vSrMf9mUpAWfXvZEFds+fn+X/AnUMly/bf6Pb79Xhf+6eIeBQOMtIAtYIxW7+NhDN7z/XyXqQYxp
uUXiLURV8oEXpGPGdIl2H7voZ4ADrJ18/Nws3PCSWN3FPloF87fP4GijVDmkOz3+ssSByCubZftU
KWw37MQCU3FI76vAskQE+YIpDfOaulqe0d83DNnp14Rdr8lRbJrUSMqMnM7iKZWi8oUmGGbW5IkX
+pTqM4eNAnuTHGd1qthKkNgmQPj77rhdDKR9FgRLEOQ27FF9KXGyB2qgCoR3Y7WiBB2QtjZgMbB3
loksDM7QcHVX6AsuypNXCRTOCV1HWLLOQ9TRaOox8fdgOr3GO1Y1X+/+s85KRlhl+0GqXF5TzAvq
jELkKrEf0BvHa2tAWisdFQ6q6TSHyUqAPI6ETnmfn69HpUPKbbVo/uuqN0vgq+xYGHrUv/jpe7LY
EEkscnQmTaEba4jifvVNVMZ930AJFZ5yTdUNA+HwYoznZBCxx1nQqINFXtVa9Kqrw33kaXg1FmcA
IurTWlKaKN7mhsaiPRfW81SL9ee6klEwbBIf31u4TxGFn9cthnE1hz7G5dOgeA/qTiKH+9bRLR/S
oriqEJ5lfjfBPsPFd6MsF3rgArSwudFKWiOEJL1tPQgxiXwiy6fv51hTeyP1mxnGcnZmeuM3zlhv
9i0TfsdtnV2kqT5hNa3YpLRHkZ/m9CB68JaEgNgGJgO2asCd/St54sz8sSdI6xcYF8NWKzb9OG8D
cfs14lFbBvvmRp7PZx6l54YDhCzwZReuZqEMlJjicIIq3gID89Fe3P3xRSh1o3o7SDcBWeEs/n2a
c4OTMo2pfwVLeTCdZOcPlB9eXCK8dhNs6mpVuU3Ua+UptY236nFzFfBF7BeXkSD06y04W0zwMQFF
hKYeaYfriL5hOZ9awKWwfTuI93tr98MhULh10WXFleNeaoMklRCfLgSjIAKZBlN8ZAdpMfFtk8zC
519lhZ1p51/29CHsN1NkA+2oWenu1KQarQ42Uno1gk03VPE97N4IdXRzozfOuzforTNZEfTOzChW
PpmGSPjBPsDe4XZqnd8NgWok8PuAnz2H8+R81dhbxZHgiBu3K2p44YWv9fbcVLpld8KXMtijm2/t
DmjQvgPM1/p81yAzURMUHLsafvmDxIxNUbBh/gst4SfOxY8cloKTunsE8s9rdbQugDLqR10M76hr
LVClWUrUPm1RGc/LCjh0QcZ9Ix52sNwj2CFaF9AB4IsmKOEo7Sgs2HYFdES72MDM9ulYWwSu2IFV
Q4CXCHDBfAAbzcZumsyGI+XhJgLCNQTA3deR24frj3mnOcFxBKwueibEL4tHIfmf1AlODGHgdOtx
DbWOiRf5gn3iTyiV24LPMmjN3gPrH0hOY44bf2khnCt9lA4X//A9uVoYXN1ff7M0PmBsYB/h2qDQ
PQhn+eZkiU1F3+pi3q35LorY3stcDb2sHdbNuhd/Qf2aqS4q7RBT4/GSOeHwTfv8zGcRMVb8V5b7
xEYfPWN+GxHMQKtTjVXXEAf8I5x1OQNHnevgldyMTcJacxVw1kn6/JmN/1zzCzyhg4t4RukUpZcp
8u5tfM+eiMZtUE4ZBrnRYRHtc+kKPhuPOmOuBLqF2UNfzkmFyvNR09DsxqHce/M3Ox8Mg+CkKKNg
9Tje2IWxog276SKJ5R7UML+Dz+LmWskz9pWaEnQVZJfi8ssyKCUwDQX2x0Xgln6KF2/WiE1D1Y5t
DLJ1M+dbt+nhp5wjxlKXFeXkvP3Wawcgoo7nmytElFyIGlPIa8heuj6bv+CzE/g/HMZcN+/bWvSr
Y9+pCXTZyMI0n6xpnGcj9GO8Crv+BYp/GOb4c5g7l/dmh2tRre8lj+105MxoOEn4H73nLJyEB0ME
kMqe1rVgGEPYsU01yM7C0cFyXnawt7/aRGt+B5tyx8PejJVwfUflBRS6MRh7RWdWgPm6XVoX3TWL
6vmr/dJzjBpIDn306nS3rlMkjHNxsa2cEfku+KaFYSz3PVK/Z84cazDF4OQLcNJukVXYR5c0eTw8
5yrEvGuFF7HXMJVv4lPZ/Tgt4pnLRZpCk47cy5atfH1yBgtybAwX72o4++CrItWK/xh+szs6ILDA
TUs4Xve2L3LkZWO3U7OP/G3m3rC14T+RWqfBSwGHzIHSJr2rPq5BF515uwKu+ugclirxTBnHlmy2
RqvEOxc628xuCezdw2O6Qq2rpkF5bfz7eUkLcXWgMg79A7dxDe9QX3AdtvuchJZkhUSOliLjhip1
jP8X9TWHWfW0yZz22VjzdiboUHvxoAZUE2bWiFAVytYizhIQfJzoE3sHIV3JR6fUTBI8PoXp2b/c
ET50pYjWcNnEKs4rAly6jRiDMTiKVm1o5FtfCNqcOIReqBLXu89Hb0AxUFNfBVUlgl5akZvH1K58
uYkHbgB8yn6UEDLUSBNse39D7eF1GdUgQatAkP0UVScNQDS9ZBFe3s6kiH+2oQogObZkE7DrSFWu
H8Y+cGrpoVv1wCYNqt8FHHxq9rbdE8GrEDJLf5oRpv8HTVRkHOGYJ3Td1ZrWzmk8gaC8SSO/3obp
+OPSMRqBBEEvBQIerajdTiiT0OsfCdgqSa+l6wroMJpIf3nfgmePxqgBUGLa1MgTObiqY+xiSz6L
bRo2DVT2jW2341jgxdCUNKpbK1Va+NZqeVFPUNGW246eBmdHwfl4/Yz/GocKLxBBfCXxfQr4KGmv
qCTYb6Ri1+nPve2AWiaLviaC1gtlPgY8Tk6LuKGhBL31QJP3kTpxB5KQMb1ZXobInREAa8qEAEd5
nou7M+wN17peQG48DnEXsjbve6EQmc/6QTq0LOmffVcIcjIWffwQbuApzAD3qqQaedS13XmRgwW1
7dZNQoPFYRCKqsPz1qhk7idbATnxgNp0z2L70WHad+p23J/KpDTgn69BXpN3iVQe84raN333iCpa
y8bqQqqMlUL/HPzD+cshSDPaPuyHg+8jx/DvOILsDRAyVFaM7Uqu8UywLLxVKrLxEzqqfVoZ991R
jyiO64b63V6gwvzxHiC2uT6mHsB0IAZ84gx7zC2xF308i+b0RH2vJhakkcJZ0SlgSqScRJa2hZZg
Pjr6cyHU3QPDf3vVT9BBQEF1t6ott6/y8z4s3y8o1vYl8AE0np87RY68nxELiJiMC80kTUf4TtTr
eE4bLOUykXElurHJ5eG/FNRaZfLAEcOiaLe75K2/34OHntlk47KUPQ1NkZd7yQVpM5sEogLj9E9b
ciD0QeeAfhGe3ZM9prEoYdmng/dsn4vD8BT2akByllD8PA4VSfswrBVlHwhAKgOHiznFoW7PljDy
9m8ei2ljWbeWibGwF4gBPFSF6VPwrl1R+cklthH7NhBYBadIhKuXaL3lCG7owY65CQQ0mV7J7qeH
Ug4Z41n+x0V/SRS0apQQIc9zYYcjkqsM29v1dqvPncHGrwNZ1SBFDudmOi2PwwBXaqa/HfiWbrYN
/DVBhCGsYYXa67gIQiWpcq/lUXkNxZiWHrdXVXEajOC6G7UvgC54a401dyRHvY39ny+600/h/Whw
V0ipbxLNNfYBFNhv+uPK2pAXh3VKnVOXAdrOTz0Q4/7lUGvRu9aFpYxNtlUTiJ/tvmmHns1Uh34m
aMm/61k36NTUClR3krSDqTO+AWHJyMJoO2UjHX8J0JWqeHILmle53ZmL3B6ZE+VP2JHLV6LgyvsX
YFmNxvZlCLQze1YU1C8Nrem5ws8z4y2rr2nYeMNQivGc4QqdEY4pFe7JWgfAULiVuYRk/r3fu2b+
eXL+4Xzoly/HvI5KoKg9ttPj9XjfujlM7Co0A4nJICO07flTvXAeQ7kM4nSMWFs9OduwP6tJsZGy
50+WY5W2y53eq9oxVuBGK0I/qq9Umi6XaGpv31fbyJtR4Qi+RTIgsnd67KoUuht60h2lK6nPyY+l
OiIHF4vTOYgl4WM7LQrTt2DKAm08vlroAGtoqJVic8QsHX2peRH0PQ8A0JU7UL5EgEUIl68MJ9Lr
qMVihOMTcin4RxUvYEDZ1E7/rNvf2/AOiCFPJDZD2L11aVMd9yegTcN+WKMIB8deLIuT0LNoJG28
Ainr6FSRBJCkS3gWL/kdbq9Jq8G7MwKppS0XWl0H1EzXWeh5QuLTgjntn7+ojsrJ1C3JaDZckzdW
EilWRscR73zyMyhN9ZgKRmx+3sZDCnAQPKGKtu81ovmz3WXBAOTIBX2kzwXqVPoPxkLmDdVKv6Z3
pxOtJQUa0Y+HhI+wf21z0uFV3SaH3u0HZ2UXxgOTuT1yPvhbouVItwPoAvhV32P6XdKAwHI/PNd6
YgqLqrd8oTqnQ3sosxhph4zF/GAkV5w3FfUm66J6qdB33xPNlnEjzQVg1NBpbeFqkSV85QP1WOVF
RQpM5cEjyGFYHUXp9RtnLAiDbRTLfqst6tWzyH1tbQukPkLUgJjMIum+J6+n1TQoT861RXmP2gZP
ueNsXLxIT98xfvoaUSZqhzkGX58O+DRaOkEskgOgfbWyeVuzHNTAKy6p9roCNfs7YUjEDMi6RdP8
BiRvS34tZg2xMn4hxOIvPIFZtO8GcfhXYioo8LtSv+ZlGOn8fwGW2J/n9X4BTfxlKMmaS6532htP
2mJBROHZJ/Uri5KMpgb7XYx8JDPGneTxqBZsR+nDFSmhiRWZMtgOAWJUsbjLn6+768nH2n+8TLa3
9r5I+4A2ZhVsZ5wSDD2qe6XGaS3k9Y50gtpkIX/kNZZwVSwObqNiZYR70rCNhqJQH5+7acwtHcMr
XznPMxTnU7s56CSh9So3PKXWaN7A15n2Pe4kTfSVfW80yDi+ktPMHIXRywf9xtt3PXzNSYe+yRDU
PAefz6RIGcdckYIw037lquvi9SIcnjHjqvD3PRgiT8LRnNTQatfZI7cr+V/0FFayC9Cq5BadBqpY
upNOgQpmfs/XQzb6QXwdK0Sd4jDJpkWnLihHl89jYG9dkFioPjG/XOlkmgtxo65KJNQA85fRN9FU
y+wGQKZugFz5hXs4raRSuLsZIdApi9lDxjH2UuLzxC0gK74gLR7p0fdGzZNsj1ECgxF9ZJfXOU9S
NI0oqWyqyABhpFu1HsU01B5uyvU3hC6xSAReDW97DUqV8osXrYNJWyayqbsAjm+lJ8Ru8miAfCBi
fDLb4e/8GNXyUDJiJYdnEsNocGT0iiuG21ihgxK/3EGlAd1idx6kwF+MhVBVX/pZdyyDwwPaWMw6
DiCuNoTtX8AlKokrbZn+YFGKFg9KePW3a66eNRHNTCBubmxftcbQmtGCAIVZCpnCv/npcEujIDYy
JimqSoAAl/G09++SELPzt2bk9rgw0fg2hKKtB8AtGFGy8ZvjXwYn8bPyIg/Z5xRmBOyzvEYWeMAL
5gQbJz5Fb2E7qyquYNseuSEOwQDSpptfqLKuamr9s8/Vfbz1giAxOHMCNEoWZq9jVrJrNZVKj8k9
Vw4P9n1bHxNEIBk+2RVIGFNfZlgB1ClKoukzR/0VQUeS/hd8SGpgTHaKX5RNtjPFfFVz7/rinUX4
rksXaREIpEuz6q2UixkbACwyibtwlEl7p9ba1xmxiCh04lxEz9pBXn7z/a07krSgINIt0fZGMktS
tS66uWry6f54EzaZuFbB6nR9pwOe1MD0iA3XsKkluUN9tBARgzevaPCUIV4oAhGciTWfKwSnD/uI
+XKzjTQ0jJIp0n5dnykDLGw8PZ6Re705lLV4oeavjnz9hgq2+OT1ow0oOsUidquKFa3fWGO9wcdE
byC2wkIkeVYAiiFCt4QYH1dxQCtY4UAWpvS0/DSzs5SCwyqC/iAqG8CtzQwy25ShksQLe73ST2Xb
CZyp2/iP+xEUfGLV3jJ8rbKIdVjSSFTzAmg1Sk8YFV9kx+E4/hKe6Af/8bGqXWdjHp9268W8dQ11
+2MzNdug8wpfqqnaYkXD0RYU2pMkMjP1OY6cCtRTqtwJ4WuGhVRxt9mKY8R9muPune4renWyphFa
/0LFpwdg8fn+HMZ/QKvgnCjKrlYbTIF0ePX2RYqurdtXkahr8Fg47CtoYK/k1obMr8GQvQzOxy0x
5jalQLg3f+C96P2Z6e1+LlI42PMS2eON4YBFaFXE5xHP0tQiKqDkfe4ZaQVgI+ulJBJXQ5zmJhIw
iaYGCs9kWariTsPosR4rOLkQ5Fki9esGUkFzWbAG3LbYIuFdGC3b/SHTLYN0qhkQ8OzGgGJXA6H5
c6zC+RGWDOVNGLuIboVDQbh9AmG2WgHqfUnBqwOfUQSy8A0dTGlgLgaCNFo15uhBXjwtmdC9w9wl
99LG8jsO3AS+kEkzqPROCOk0jWuxtPyjHsFa6wqlZ6XlBBy4vwLYIpgNhtlHrlL0yXbpORx09pzX
SIMFSU8AHOUzeZASh1T3cMJ+FNxtOEeXdZAbplA44CyFFI0M+SbX9zdRthBdJ79f9+QobJUgTJUg
/hU3BsQmbUP1ueYynd8k7E80J1tieOhFjZoTfF8qSV9Hn7LxnZeIwHL0z+JJelPKg/ghxE0ih9vF
c/H9Unq0PacjGKIIle4nI6ISmUb5S85MJ1WuwfV/U6z77yGSKTV3NnkegCeDfwQcco0X2dWgQOTg
ncGnuQXLpI7DbYQWFTAMLtYkgWVdxH2WrlPnpHqSdETip9Q0H8uVZcJiaAsyb03wHp56ilk4FjPZ
7HOW06tT4ENC5XNPN1RzRM+RBClLbhEiLtojsBcVGRgjZtSvq/xE6NWeXa88WLpT6EXiflEbS5Of
6AsofaF6ROWbp24I4XYcGfNLf3nzTN8jsLXRKgecvBmZ9IFU7ddpICE5j+hzEfELMYwBYlHUhJyK
JTWwY7ixf2TadgCgJVI2DR8kyj9K3YS047Ed69kpLIK0snJi29/Bhj1Fxam+zsbS2keu0QMsvFe2
s5MgsT1DiGQZyAE1Tmng+mCqOcl/hI/TxIuMFUdgDEHQDpg5RyygabpdzLyMKZe5x99m4iigqm0i
osEaV+RAf6ST37ozNUq1/h1KRsKC54KHP6V4GN+8HRZs+pWVbsqaRYJ0u/q1CEVcpW73aB+YtP7Y
9NP9zVPsLz2YhHO2bzBpQeNKzvaZ/n+KBmZ/nTaRR0+uHFATpHiVwUG8ItQOf+MfH/Jm4VO8Htzw
FSv9zflaqyE84yOP1jJF9yCAAa5/MI4Db7nc9F4zbrai+Au53g2A4QOplh/7dPvusR3xk7s9t5t2
Ssq70usn8x7/6MrPHREJ5FDZYRSIaJjzdKLDBLyS7zzWkbUrNNrKFysgF8zDr7CgfWetueDszBev
zdwxM8K+nd4D/1Xm1nC8WoTifmTatpPxH0BMQKwpjTAWec+VGIGt6L3mR7JJFrrwa2xOgWxLtK8w
ahmdYJYtR+g3Mpo/WrBwem/rLt5XYPhvI7dS9ZZGt3BUGdGpfeMpoaH97oDEZxhzUA6McvaxzcN8
Hz+/kIH38cqlbP9bIwpxGOSBxqWUaioZwOGaKFrcHZT/58UT9oxWw1s1DpmAa83z4t2Z5xSevGTZ
lrHz/Zi06nExB8R3ALI4VcdigdESkfsR8hlWXQ2DSDCQUYAmSKCA0g/6vU/ewpbmE4+5nUyzN6oM
Fe9vPRnHHqdUnfP9bF6rtNk2GfmUfxMFFP3CKcM+3k0KLW4hUo0UltAIjHVDsN+AlmAiVhkAorzE
7+dmijSzd9ZTyQi/KLgVuH+7Q1uD3yVpOm2RrmouQbLRmybjtMPRIA1v0ulB9DzycanJ+062onkZ
M9pknVqOTUcbv/wvb+0Iue5Htvn8dZD+CaM2mwUbufU76WUskhiyVRqs7WMeVE+ZXiXQcItga42L
h4gEIK5IQ0/PKteuWjb4/QF+l/deMDglhfe/IIZf9JpXirsqPiaM7g6cMezilD1Fu1TqjsY6E80D
15JhRCF792gO3AC51im3xXs8q88uslpG/WcJr7HV0DTnAGwdmz1/RyKROyOVFQ2MTooTEeSdxIkq
XgekicgeUkKX45QFBe0SzJPvcRuDILQo4FJ5UH8NW80kaQ5/sinsA1gJtbVaqHmisHDyEmTFCV6q
qhhm70lmkS3v1nYfmRH1IotPnXC9C+RmcH2WIGO3EWtu0dTbJHVm80vETr2aQmuUNnS0bxjjwKi3
H7InpZrm2BR6hBdT6Y76bpJVIeh9NliWwA/3rrHwIxWvqcdnrit38Y0ZPVjUNwp/TGOz4zbOci6v
9jOBvS4q+A7Ws9n81aHMZCJNMUH2Xx4WJj8N90FDEXKkrK5zzMh26R9Q2A0oUbiifWPtmf/2dqoY
UR/Ilk8E2KZ5SsnD5t8k/3BlrYem5A/Ukn+wT/zJg0e6eoPRuje8mVkGEJf442QdjSqzX5sdv2sH
voZ6abM4F3qUnROEDdCroLAQ7FoUfyCtNYNIiC07mc4yBMpeY9jVk0j6vODuosBZnQ0imfwlbIKt
sdsHHfp56Qv54rPTvCstNdqlBsQ8k+TkbORlJ4zMJnvKJvKPRKEgRgEuO3yDpFxOyf8WNn23i+Ud
1dyWytbGk6+zG4YhdkYPoTiEgjn5gy2Ffvw/jEklQEMl+LtY5kwJbQ2J+FlZ63ILoDP/IBbGvspR
7+WJWbGBtvGbjdaraYjVmzwtYhJixGT0i2Tz90ulqj1jTDj+9mOjMGunIDHPdNzNXroZ31ks/XdZ
UPPvloTbrvLMu79vNVQrdG7B4jPfzHRQL/YW8DoJBIbmChb33ylVSzkDljVl2hed9gZ/IlvSOYGe
QX60L5hUFV9Fy0mSOwLuVshio1CS0YPZurF0Y04QGtqok7fMVX7vU8NiZETM2n0AR5DRmvG2on9F
n7vG7Qj6/ck2VUhYhgwPblvcudU++5OGJQeMaXlQ8TAw47WQDBz1m7/QDOyK8Uwp6aUT6G7jkdd4
5AjpRoVTePu+/ErNSQiN5uc69bOskj9vPfwybM+NSH8mPEZTutFJYEPFS7cK3PogboWujGcECycC
MmpHDF7xL7eK4/MlBgjO0lqKOf7VOgcgd/98NUP9rqzRhmdsjPqACtNACMhJ5xpW16xF0uover9P
H/RNW6vE6QjK7xmvzda3uhlmOObPG0d4DIFer5J9zlLWxhP9tyFIJ5j+2VGId4EQYZhw/nfP1wWx
7Su/8noVq0RIsAhLd2nwXbquSU9uOxwaFEoKxgdpM42XGNYYjrPU60TfggW7Z8PMPvUhGLxHZgXr
oYSu3JHxlxbp4RI5MQuGmv3zbhSyhJ3bVrlHNi+/5eYKRcWtg0/rq95OYrnOwqdRfyMYHcTyBxtG
hPceOglFpX411/cMdcaL2iFzDoH5x/C7v3y4/YCs/iQCIZ8BwYS8cNFdgAZcDLvk1rjEyyzzBF6w
Cw1o7oR9JXddxDDNHZOjUubf0NTaFD1A+mICh0XJrmYmDz6KXRLlf434QR054rLUwR3NmskQxv2a
47NKUwnxpcB9hZNn4QiE4GvB4J1syvOBC1rjjFEB2dX3dVMVCuDldMRw1OVk3r/eZkvYOlb47fXK
DkbrcVOrP8pSa9Iw1WpKA5kLpe3YGtb1/C0Fm8QvylsXg+hbFQ31BOjHpJrm3LDL/AGPz6Y5u+jd
sxQYzI4G5OTva90swaQy+E03RHdQsgiB6XwgBgm8ZG/uK/t3hdsCslRDRiw8DFi/91OzpW7cEE0f
/mYD5p//DCMdBKqsDJ/JEgEiTXXUSArVYwFxu1tPOFr1ROTEY54VdH8+6dRTyvA2aPIINLYEd4jD
LFp+NiEpDerzrJRaYAnlbRS67M4r7N4mQCDlv8Lq8TuLsecmfzGs/CtEBDa7P9k88vWToyyXRxNv
4VJUfMFfpT7KzhBlkKNZE8MPggqAIGG1pD0l06M2sYvNFVsRwCLPzjpiTRGCSVo5KLkw+CXdPbOp
RA3JlbsouuRIHTde46azewmX/zeH8DqhCLxsm0DqhBQoXJJiutitluwP9j9jR6x7rdj1c1zAKhY6
4uLiRNqpPHJOT2nrMt6DkQC58bKzfx+R6c93oEndlqangX87974W0h7iMlydYN5lMwhLBZFjgEIG
gpx2XbKyI0Ztmg5b2BlKF7jCyvT+CsxHykZxQUxZEWuKzE29vPqtlx0NVoBvAzYX5txW5znit3TD
tD4tllugI/y3vGMu9LTqbAb22gSi6Bq4zWeHG60ITSoOLp25gZ968eyxpv3jqhHCmY3KXlNNRVkN
7ihy1REFl+wh4/OmdTBHgy+tk8S/dvlzOpAr6gi+evXRlXiQ88w+pKBa2vGKtsZj6afaelyNcYJJ
+trKK9KUrPBwvsiprKlbo8ryqMhlNqlaK/b7AH713AFNSaMA7kNVwypd4UNt1DuLc6vZEPD6ukPP
D16HTa3xjkgMGswFYnUPNV4h9x+Ywr0P0Af+12uTCJwJoQx1g3iuVfZ9WNpuxHbmc8qlQwgI/Nl+
/zMYiyObQB8kTNZfXCaes8JtQciakQ+g3SC1h79RATqTWBDbxaPC1FtaY8sBoZFL0BLQeEXkSmCJ
Y5r4z3X+IKx2XL1XUZziOVRpNN4joGGIcy++mmmRjBUBQFvdaJ40KGn5hJfoKx3A5m5jdAXaNXCE
7tbKGnrG2pKD10DiK6REpvzWZtDpXCGgM+VAOBEmSIol5pk6abP5qNeTzNrp7P7Cn26tV5O7Cnkg
CQvwEvrk8yNvNYsU15vIwJbmAxwAoLqef5Lyvjtl0ulCFhRy67VQvFU+INKFTy/QJ6xJ70XdUewQ
D7zVtqI8TgX2p6O72OzNOzIJ6hKGLgHEX9e6YLe6SWXL+T3t1LdJxqxAa8Wg/ANxjdI0X60QqSm1
FdjICmQKoUYgcVoad7BPnzbO2mT2MWhS+b84t8HqEXotIGkvwj1713XfAUTfyKy9yOj3QDoMZO41
EuQNpkfslP7bcdpmWTWBC7TtLzCl4oEuEN50PY7DMRDTUlzXC4ZyVhUGFe3tIdAJlK2/Q1OoH1Z+
4NfUaZ/ZY/hHGt8jKyL2gVkriwbjYHZtu48m8Q6tfyWGypgKZvNIS7nstMBnu7UTs/Rac3iol+o9
Ej24Rs254O59kYJ+FR8zVJz3tjPpWGPS7BMsyk6os3CT/rNmOGWJwzJ25HAZXOF7uByNTibd925X
RenknkmOpPptDb3ZNBBhGSOkEdpwQlN+8NrqB1PRmTYGChhFgBRGP/Ojq3ytVGE9oIr+64l0Jw2i
Xb4uWQMGkJbst8xpHRgXGZn+Q9eApgL96i47++/y9der/DdYV5IEcWmxyDle8kWc/6dWrBOslpQa
D9wFnXbn6Kymy/yPIBjSHeshI5O6SB6STeqwP8awzB/UZs5sc6lgONtb1W23aptQ10Eu49aISJ6m
ba6OWCAYOFluSnmPPoTuBHqlGVDEL3Nhq0xhTkDOgb2t8WpqGYyJdNndZZLyZUe4Ni4RYRmcyFCR
RyfBnEBtJativMf3QjXAN0CyhOtkxJsjrHijTVRHthm98U2HPCJgJ6xvMSb9yIlRel1aLDQ8cFbg
3uuQ06kPQvn5Rj2X/l3/z2hQwop3AomwPiRRWdlm60fQX3+PQJJQsRKyiWQyHckxI5AUdCIo5HXe
kytC0aQZeKycFvqpiwAS+bgiLoJ4p8puCncxnuOH9lAvzBUGnipAP7LhBrY8l4BnyMCjtki+llcV
VrMmMCx1OennNxYoZ1U+rxX444vXeIPo/7QrdLSnuYeaCUJPV8zvdJJYZfMsZSIL0/rWHYhvH3Q3
sEhiDzGmJem/WD7uZncTFOZvzZIYEDn5aurEANealpVgbQ0Gi3uuRTdzV+sxymg+CmjDbt6MwASD
YoB1cdfShYhwDWZoIKqbw5+yAQ5B+dbYXo7pulpZFp17aW4baGdauc7SpGdqBgkfnJOzf9CGvOn+
9MkA/tgdT613BTRMKYHqs8qZra1+l+ihJVobrChuXgmq/QtmKaAlMRZ74rKymOR83THFdfKWQqC0
h41hTbTfdrKt8LYWns62dlgTIDamdg+XqA7OlGFwxKibpS9zJaZ5Sg1YVuGfNZu1iE56KPMJTb/D
adpIgyR1ac5o92ZyFyioPJZYbgw8zgtcpw1Rh5oYkswCgZKWZeyJAQlhdfU5396kINUpftd26nDC
Z9m4lwar1tdthsazQELS9RWsaer7dKb/5kva1bY/XUlV16qXWbXfJxlcdzLtsmENWaygOX2B9Hma
jbN4zyv0mWyJ/qxjw+eSvXqCXwY3g+mcrEHYvu+sPJO2vpiIOwbTJEPfQ1APNVyWMuZMgdpGUpOy
JAyqUFm7G1ifBF1rn5Jz20oZedfTlzLEQorb8Retzwd9dm0tD/5cRhhlDmRcGIdOnW5BrJ85SrYU
poJlogkSH/Th3JwlJLBkczTvUHj0NA3hTfV1gUTz254e04hPvBXcECnfJ2kddsUMEzafgbcFF9jz
FNlsqyEgwmfN/1RVX7RUYGpss4jvqBkRb146+ForfieJPLNmWOjlX/wnMEu8ynoHplhPPkRJN/X+
EMcFVmRMLY6beVHcnkeKAMamRqJ/YSwDllGu9noNNK96MciPS+d4VU1tPabxD/1XoaRBu8R6+oif
2EXo6h6MXO7UPy+r/xFMzHEcT5ybQzrV1pLciJ9It5Ak+P5JgYTlvyyamZ8LxLgnTo7sP2T3ok/l
jP83l5vMSxq+8C1Di5kN+Z6aU8F52udvgSrjiUvZ5O+N/FDdtUFMbaUgI+nvgLvOcoL3+2hHW69y
+MoS/If34dMDe26SsYwO0ahcMLU04w1umK+bXQBsLsQnYQm1TgdswyD3E9Y2sYTqHFbJ/dshCXxA
OBcqxKvdNNCKsVty4WXSY1CnWA+MWd8H4lBFeyTH/1BJV4x+QwdcLYx/pddup5jzFebvRSzwEsFl
z7/p5BVSp6FtS75pz6iL8xgpVJqZ3XFhnPaV37+3H1gHykOe+j/F76VSodvrRdAFsMh7F9iiXB+t
PumU7eBfvyMcYN+Ih3U+OlqhGzomUBgVzPuBtTG23ZrHItmH+FfmzWV/3+DOpDLwEzOPYoMsChpW
lMtlnFZLpNTZymY7dFZ1XYxU3n7ud5WQBuyOdfjutsYixE9AGJ8Vjzb0xQQOlwOzU7VxXaXtf20e
2QL2Uw8MFkQoGfWROkos+roZhBs3SUNzTfBQZvGKSFF1HasQiSniEfxRQzVdAX7OKuQSQT8ogpOf
eYxelQO+/SaqzWnp9O8Vh89TgrzF2wHUJjvz9mz8CLVNi1wjYUMs3ImyYNXzhZ7V5aLEgs+yGEt9
IY1tJ5mj85uXeTvqYttCujltL98vCdjzMyHOHQ6vJNoWQlZIBiINIQ3YcS86yrIlu2XemzK3NVHD
7MJ/YcvB9XXzgXf0vCYhP22JOhTVQbzl5L6poSeV4M9MSX3oGjZwhSJYD8+vn6qf9nDihExsxnuv
TentdSgoj8CeCYHAmXWDPeHXq7wQDHcWcQIlOvABiIj7Fq6++CYN2ViTN+sQ+ctuMn5g9+2G5ezV
ojPKSx9isu1Dm3WdN8Y1iMAwEsnRC+djLzFFqmTesptozUZy1laoNaOUdb8iPCn0gd/lj7CPe8CQ
p1iX7rZ915ATOERokMa+n4gNKGtnUjxcW6CduuyPWU0LJ/mY0uJxVT3w/rxz8WSOjuTACL7Inkoh
TU+nJd6kRfhb3QLwOvLhGNOejV/31OhTHid2HpAl46hz1hPBwD4R8SmM09zYLlY8y85Q849jZ29r
7h5HCA7mU2DmEQ99wEIfkt13aex3C+bVf7sMOUX6ralRQ/klhIJUWj5T5E4QIrxe913DSbNdV925
mBU36fscoh3DulasB9vJrEOJgnXnDO8V38PXdWwbOSilgAsl7w9ps8loSO3UM/wUJ5XpftrvN6YD
jqhqCGqP2s0TFKMjx1cKe2GHYwWcMLTQi6koHnkdbD/ZZ3z5Im6HfzIIDI4Rlky26yPtH7DFGG6l
6hIQHqLSrnRwM08NhEgBXO3iDTjL70k2Qav7VkxER1yGyeuOTFanjaCx9bLXEx/QAsoyarCB0w1H
G/0ttv4/SV7xQCh3dLG3oUk4viM0nCJLq3dnKDXBFy/c6hki25Ns1hEbQHKgmZeuNnjc/C24du9l
fUPqvlO4e9FshSQ7geJGtRrQOpwVXLb5TzmDddJk+V4ma/KJNwzUBklUVG4/c6MhdtLIziYCRYVP
OOa1DPcib+DcVCVamDklCCxjdGSUMlX8SQKv1WXDZ9Huv4sczlG9Vb/g+DQ90IvVCQYHCZ9u5v/+
wESGVZv65KMMgheO7zg5baVy/Rq2dvobMC4G2kPAMODUL4FxmruIFZ3gLE3KQdMDTvrXi5alwTmA
6h8CYABoW5311fhX0lAD0pxdoHLG9pyus77Ub+yezyY6b8BP1wnO+WSVvODWxaizh/wm2FyTOgtT
K0WzeQpPPYvAtTmB9vnjLyCTt/G4DZ39ODksiTwReM8+dlQZWEl0mn+yl+8lhjegi71/ozkM1Ia0
+HYHA/1+00b0Fl6809jqFl0HaG49VAHz6OZg+JnLUG5BseQrySxrcugHmBLtBPskG25lbrBq2T5Z
JE/2vNOLvboHZhHej2AAVn40Hu1ppK7+AAcVt4ZH6hp5QlmPhENw5s96/wjgDKXVLGF3U7/1GuGV
xb4A/gqPAxgwdejzpKgTj9cbCBMRlzJTz27tOtdeFqje7HnK7uQplHipOiiDbvbHW5jBDZIMvIHq
Vfu/o/++Jjd4tXInmNuLcReUWfr8cq4Kwgv3RsXwqtbepl86LPb0J8vuMD5bwUz+B0u3meJu3lT7
XYUie5HV3NDwk+QFBDYyReXaKZLuz8QpHq3R7z9o9TYEEOetFYBSuuqqFTrv7L/DAXK/QFh945Pg
qmklEyapp+vVSfz0VhP+jhiGiVRuvQmWFp65EVMX0DLOubPQKiF/Cr6s9oZOOwiqDqtOlQj/R2NA
od785tBs1HPWgdABaVqHgRqInPgp/WU1dTvtWOUkmvx1K1+/JUylyM69A/W+3Uuvh0YWnrjkKDSD
Wxb/RHD9o6KInxI6YyEl69YBncgpcYYbom3kVlQj28RnBEaqiUlOcAY6DkJEvJWSz8N2dEL5bE1o
34NEENmkjZUWiYn2m4mw8X9AMFh1QD2WySSeKY+SU81XZT7tSm9rLO7cHjg5fzXGrVqQbuTZ+oBC
nI03pheNSbLakHITMVHHighNhuET6/XLxnUW9KYGhjYe/kpK+Wla1KpAn3SccvZMGytcq7Gkw96v
wfEZMScVOpbUvqBoOZG5zROVFaWoqnHXJQm8O6ot7bVNvVSBCoS060TT3DYN2+v/QtAvmN7ubGdG
v5kwcdQ1AezpQ6Y5B+KGseGFkGK9sNUJxzJuBUMf7qOwCPqCfnOF/cHdq0a863RW5fVPmMS1hDjU
CIkOjH4N2x6PzIhfMensWbTaa9VR3skMJXZAk72fGD7mwno/44qmfWzBVhbSipCa7zJVl+IzC7GA
LykgsT33AScA/KDpZF6Lov+NtINncYuQQY1dX1WmHFlNrk+snshS9Jct2vQrXB1HNQkQ4hVnXDTC
xbn0y6cNVzqhYqpLjKGT4b4Lt6siOgvJiKRTDSO7dEc28rApvOFcXPirgdskEU8VtcU6IklFcw9n
QdQD7hXDo+ewE6HW2I8XjFHvGowyGCnWTG59LL/D3/dA/vW5RBubJh3dtjx/I1Lf/sRPFuhEoVcg
DbA5xq2P4s5JaUk5uH6njTDfST68PaiRXYcdv8IINyNVpif2n3GFQ4Y51Se7WLInH8Y3KgpBwlQE
FqiYvBDs26bthVeaAOyRgVvI2EQmblw9v0O0Embi3P23JK2LKE1vIbNW8ag7qCpIozy+9WLv4U0t
KL4nFp1earg+WbgO8VM+gMIzW8XE0DG9X7YQZq5gTX4M4kQo5OHZzc++5w0lepr81n/0aJt0uoiC
sFkUz7qIyxwKqC7YdWoZp7KG0HUZDrVRr/BGpCQaduQ1D6bwoYbZ/GejwbXCA/m9bywCGD+5b+2l
bEiI8rgKEBqGX93gn8zwlTgEhDcRvJISZG3YakmhGy2iIIULViMst81as7dbQTKB8RHOe01lpOe5
3tJriIlUj1DC4SpR4CiDrmSgKp2PEATFQO1tCmcR84PHhHwPfQmpnqQm9+iBPon9e1dGHXNDSHGC
cvvfITWANI6WUIBa9h/uqzCMWg1mkNWqabs8v4Eh1ldHyxI8TAG9gfu9cZzRfSiqpFTgzVRV8MhY
cufU481cOQEYETfVZZKh3bfsmlXLKQNV7K7fTH7tbQWH5GBqI2EuTmP80RiiEdsFpESJF5aHrfcz
jhZLxYpsDvRkOCqYBvVqO3/ks1HH/mGcp1JzpJblbz3CPCI1apiSMhIIUoX8OZLQmzcMI7J0kqHH
rdZOpeMvA/aDtr4J+uOikpip1SHFSLL+Lx46c34AHMU7STFxD/njq4AXovjkPd93lc/lbIMxbMpv
CuCJgIWFQ8kdt6j8VGbmtPpogdGETC8xyFNtJLnY7xPUOoSLFotcTC3hcUKcpZOZbNkQ3qN53iyO
kHPHk9d+pxKVd/c5F/OccWjiLCAcfbTkaAIeTLPkGyIuM4dv1tb3FjOLEw58onigrJzY3kvJmYmQ
AFMTK3EWVphubpu0GhaXInMfhuSy7I8luVjJPZEfYTgNQrDgdrMtt7r0GSQt/mAP0cvc1fqzy44e
dx+MBZedYnOuPu259Znwm4euAKKGCsUaVwp9zp8MyiZUa0BuW3zAnSdDKS7XzypfbqEylRID2Wlt
XsKR1uEJIlDsJOz1YiLklz/sURxP6rKUjVC3HLUH64AGG7Kw4TPn1fCQ+w6zKycWvISLnyK89D7w
q5pZ2YnXOz7nhwKjY4T7dXbe3Sni+fCqOFtxOjf2i4cnuaiBluLKJ9cOJp8iINdiCd8tjUZmn1Wy
4iDDyWgqJMO7my5mlwLO+eGF9F1qvqnwjjOkwRhbnt0Q8CFJFJfjO+m4XPWy6bB/GL3Ugw79YHER
Cl/+lk19VwQYdoD0Y9i5e5HvF7zOkAWI4Q5TFPb/KPtMylWJlhlLQXDcCQe30OWVxHDuf+n36mMD
EPk5HtM3/IP1SV2iX4N7BPpZm/hA2iIXExOK50wlIH9sFAe2dAaXMhwLH7o+n/wqYyAbP5xDzlMw
XvIm6NikMegg0FLy0xalCDuofHWa1+R97KMfUrTNZ6+qkhrHTHo4CDTX1E9s9Sq0hWHZ/QYcP6fF
yP3Xac2gOn372DnuYoS+MNtr6u9a3UvAT6nDq8REt9Z1/kdcySJSEBb5MROXFSuXQHx31AmSZiU8
BHjzbwb24cwyohs5RkXQrzn1vgcN6Os1NyPRspLO5hzvbQRN++mmS+gJV4IGSBVm7F3RIcJwrwIy
kmBcidFuT050XJYAJVzUgrlGPlzsBWIK8UvWv+n1LJAvYNRH7xz1m1ieDtyFGlgsiaW6k6H5RXcB
Xrkh6pPt9l+4JKHtRJzCoKMFUPr7W02B6eHVMSifOAKNiZ6/U4Ma2dHdvtOT7nIhz7SzDH+rhigy
y/r9Iyb/7a/1L657BcYP0zahTtMp5LSTREeZEQ9uSPMDw6VZVqXFqoBh0mqINmFyKLswIDUwqHKF
9x5vt+J5hky18rUc06/BDr+sGGc2dIUPqcR67GiGxdysyyo4BxaZi3MO7YQYv6gmzMppQXeACNL0
z/MPMtZR8tevCtZD93U/nQMKGXBZy94RTJyvnpUCi/4SL7V8FJe8xm4altslozHjsFE7eQZujz4P
LtDwVaSxitQsSH/jlUlQlUfgzOlzGGeOgdFHi5+N8C8FnePS/3OxcLWY0CP7+6treWmVhMrcq+Yq
bXr8hnHEcUgTA0j1j0nQqfnjyV+ydW6zTvSsZZTXMNYRUpR25xGggYlBpUTOyMcFfWG4N/TIvlTG
Z3/Obk1b5g8afX0Ra466Ttr0NMBUxmbkZps59O/auXdMaYJalBF2u0pTelG6ib02PD30JtihSiuF
ff5O8nlFnU36HwXPj1UHpoobfyH00iwsEPMr+Pi1/Xt29JyO3oWB7RAa21DkPepOlgWM1Q3waPWv
oXKieP4IY+IF260MssUSsx0nXrojm1kWZ1hD4o/vuxd0pcOU1Ibu/bd5fbXBKkeEXoRQ4r44TC7x
3YoRjgMIPoHgfs3I0wh0IFLOtRVec5RjfHxv7HncYpm+P3cYqQwYbv9NPHqmhILki2kamhzII+m2
xtbctVFjNeeKIM+//a/6WdTLYUDRwqRl7JR56kAadkATE1WkK2W1JcNT2yHDkO40JCMO2Bp8Z95g
bQX1y1nz9eNjzLm/gwUBPrdDnpBeB/I2PmS9f7qvN/s6WiGT2yLCUjP7tb9X/d52TtE7GRu5aBOK
5E9giMdFTwjsxEIQ9JHcDIZzlZtO4J6KTbD86uLTIZ4ZQmQXPhn7MxKoXHCDSUPRNc/Nupqg8h89
BtkC3fVKqf5Hf028oj0cY/wTxY3yPEDC3g51Wkr0FyvgSOztQBuGmgWpD3r5OYysW689Jkq4mjY+
cdLbZBHgyCm9yD+SfeKiyiTMA8NHJIP+ENO+xur3sMZyB1I98GaCkoTWR0ixGgLsMui3ms/Tly/g
5a2UqbDEJ/uOEczj9teAoznaOeuYIOWwTcFCxqlg2VXfgqdKuX476hFunjc5YqndJ+55qH7ABew9
ZpCmJ7LiSJAnt+BBZZfE3tTKiD+ArUvDnKBWVCDdMOzS3J1UHRWxgPsX34Ba7ElHP3uQ+X9eTTT4
mSrVW9AwrAQO2tTFaq5LL3b3XwVbo5MiRtQ9ogQTsdBsryfQns5Cd4E9i/m9F/UhruXf8MJ5PmQC
Bp9wt+fEGwEUQa2TQbHsdgDy/fJDTfFnyEB6Z+bfOXiq/6ctcXomHOHt9J+sq1JJ5RBgyI7ElaPD
i7I35oS4vY1WX6D3VeMWnd+xxAre4h1eERto17husv7TVAepPx/f5TxS3oCVhQtHYz9ZEQQ78VMb
zMLjsXO9LrnYOveSbHNlNnRnLtzvTrxgNRVy50tanUuPYGIz63TgGV+dD8VqB2WhvN1+09JZA3CZ
gTJpbovW+Ey57WrbUM3ZyErSIzIVR3doJ7atkbx7Oj2gbyPWG/dMOl6KTvHtSv0eeJILs6Snh/lN
Qg0H8rZz44u4SjEcx8qGcaLNpx1hmyIwQCmDr3GIIaeuWepL1GySIHca4Z7JrIyyWmFfyn+S75yU
Ps3qH/g7W/onFWPfOpYNRN/6qchnC6zhfuVL6R3B+BFTI375ukUBFagpk9AGfW8LGJM6IuR4cGto
URSk1uBFaH6MnrpV+YzG8YpzDhA56kWu2P7nGC8ts8HU3zPK0OIxLDoonHAQEhYYoPTU7dYykInl
kKsRvH9fXSksvnwKC28hCmv3xOQ74M0UCtID1pCmrIjBRfS/AhxsehajoXhp/dc3Bw/6bzOUsgiT
ufJnCUjNQctwCMz05AZkUUfUdpDozHk+xT32M4B3OSB7wESyNevsayNbWf9Edvft8dOwei4f+sc+
AMPOaZPMHJr6f0uq8YQ8KMFeanBdXSz4VYKLCL31PgoRD2CluC7jd2O7WJWqEIZ8dtrgWeKhLwAW
s39PwGUL+HVB0Jfr0bfERsfkZAPlZqRFpJmG5JRmAY6pK2MWSeL6+sxMlwEiA9VA/LUhAZMBjcJs
r43FH2jA8fArcnhWfP1OcUVVAIV8WD8WTwOffrp9YJgx07q3qGMIjhd9JE9RBsKT+FBl/r5S9YG+
5DKd3ltosTBON+yeyGjfmwh7By2miPTQxkdWJMSmgT8MWPmZttJJZ2xHUGFHgO2kExvAyjyJZ5LB
YABsSlhv17x9lyNhY66sswo3GfDagZfsgvF7RcdVMIlPj4D4bBbjlaz4Fl5/Z0ki6eF/xbRiZ2q5
dPpLoylPHwJ1hOgaNLc/A0EvrCXY/J9xBoxahPRRHfroOPfm5CBuJVuEYyBL7rkckceqiKug6S8d
BjbSvLlBo+xRIOnOZe9n3LQbQ47QBQAWTnoddDMQC1rp5HigrCim6zKJB0MqraPF+CarVD+XZa0W
fuW7pOE4YO6G/rzVHsVJAwLqRHWEShVoAkLM2ng+1kJhuYJ28wd80Ragh6pum32sWow++Yubxice
QjCvUO/7WyYZOGQbnohdndq4h2c3WZESvoJ6oRRwBp6SpDf/z2kdrmYjr++4nPAiMkJpqP5iRyW6
hvbKqNBSh28zAUCtSQmX0Tdac57XnzofOrcw3yHurLyAX8Vls3ONybSW6s3AHm8SuQzBcn6cXJpd
hiUaZTYQltCcacggZ99wZwJlLnh3se+w1DgwACJNDmFPV/hyMPgs8QX4Q4eealHtkVfu41rrWQFz
+Vf7lj1u8Up8hVLR4mc6Vl9Q68yG6NXDJiW8Kc0y2b+ymsgOU+XiU1TLkvqT50L/7+3W5V/isyOI
CmU2XWob2efO2YFkS9Uv2LuRjdQZFwxtVCwc6SXtucApe/DPSPGahE39pM7FP0bu2A+JpVuZn3k6
x5A+2nIGJYy8QL1Ne3BfUzguCeahoxxJXFmglhwcX1aGP25qZUE0wBymr+RwRszK0SHW5f295cFr
Un6LANycgCx1pu3kJRhu4tBzOSQrIWkShVrPBv8UBWhY0l8lSEGrCpJDOdDcVs/CQBb+t974H9UY
2ePXg5eddOCw01XD5FfNxWqye8uyRlJuOqCsGYbc4hnhmw/rvNbecVPadWMWKuu3AIBg0T/jWPhf
p0TH8N2bXXcdhvaxXzG0AZZzKS1TkOQwM3aeg+E4KbYYfV4iZk510CQ1Yfx2hjF3D71xS2l3ZGXd
moWiqFUh+6QwCj4gQEuNpAKRuNZ7UhftvpTyAO57EFVFXGHXGYT8aUzWuofWRptvnIp5gDDyltMs
CG+qnmwq9or8dzfr+Xc9sk+Lc6yRj7UNzre8BZy5NEdx9hVO++u2AtSOaScf4ve185aXLp8k9Tb+
vbonEJOSvnvINo8kn3bGZTGW1L6U+r+78Hklyf6M4MAZPKQJfcEGGeayYC/aievCtXnim0BCK+Nf
+FCLuavC1+A1d/f0ineIBt1pytGl+n/bG5RTplgP47KoEcOiwsuLl1bINBvimJXhFqvkTHvzy0au
LCJDqe/blTRXnp0pnWgSpi9vHLNbChXbNnx3BvoF7IWzrj3HeB43UahxQt6+DhbLjIx8pq+lrmZ3
C7diXyyBCREWMk5VUtYDB2cAI5CiMKwOmVaXabeC0HVm4g0/fPEvtTT7rxL/a181/RUJg+OGEiuy
0TOlisqFhravJvoE8LsgEIsUhvgO0xs85kOzB5LOBCdE06oMuz4UJb79KxaokFoTW0kskxeaYWOJ
YP2RI5tfmdvH4rdKFxabtAvVO6fTALp9ljvDPOIRYvOFin6pdTa/LGui/et1VlQLI9oLJzbAXxdn
9/PkshtiBaErSICXbz+504b3VKb0cFpEDaB71Y2plbVNqEe88Gl1aHTeD4Vgv3RkVKHeoo7PCWw7
UGwM/pJFJFPRB+jV2USAJy79cb8N3QTJtpfWQZSEnPyD2lhwh+8KE1FDlktbTSzAulFQtxUIaVuD
0P2Ht7AS2HW4R/I/P+m/Dqn1Nd1YbfuDkKYeuOY9xHpxrWQPX9r4lQP3Ttwt7gQVSIyCrNfEIiVl
xB83PPQ5rWTa5SwnG8dkrEFBT/9qF++IHoPpGNk//+8bnStsEmfx7tN7Xkc9wyIeZSKvWp/Zc09y
N+1jLNQU5l/+tpO55/guOHxRgJsK/EhqTIKd5fa9Oe7oszuUm7dNs++Jn7chsScN0thMQpgt2gG8
aiXwda9QBoKUw8eYRddPLKtF9JQ/tFf42MWq5cw9LsDB3jfCTWSOzDpKfLd5fIn/UR/SqDWQIQh2
QZkSqu1uxV3ZeOmPw2fbPJi11kTzPo220nM33Fsjhrm78kwe+HnhONvJgX4VM/QIKrbQT2br+dXZ
UAq0QZMcr751b7CzGYOTrgJAbfQdFf5QSOOFG06aiUk/XKAGLBwr8gLODmpK3057Bo5OZUxbHSUI
4uyaSk5Ze0JuHvvZxmjoZQLf382tD4Gwjsp+rcMORXdWmI8kbZYsO+KHSCNS39Olseas+z3YHdg+
Yy6iJvzR9OPhI9nQjboEt2KnsCwjKNrgVQeYl5Zwl5Ih+HTNrcseiyZYv7P6zGzSZ64y00Kj2FVZ
n/+P4KyHZtnNknHzX9fSm/ElOkPy3O7TGhSD0EL4jKtGGS1dfEaSIdb7es8EfOVHkd5O+4j8M4fl
jTUQIvxI96ZmzRPdykTHQP/G9onX7FOKL4GxPAGOH/IOjcGGjVmw1qVY/Qkr7p6RMKw8Q1kTzGk9
BIJunmAgR6UIRr35NLn5Sv/oZ+LDT3TFSl00omtfiYr0JYyIDroRXuNpL2AnoJzwqlqLkrFL3MUz
kgtO6oh91ML4Gv58dxvigH4axrE0E5ShpFDFz7ak5lkcno4JjvKeSWCKlTPSbhcj/i86jpU5E7pG
QRtky3HA/WTZ3n6wZZlvfHhD+hBhc80/ac9UYhC3Mz2EEhBBSkZNqtH3fDIpdJThkPYwFuV3bjPM
SW3YnrC0MGz3sjLs30zx9KSX2MaJp/lB8H3AVc62O0C5laJSFDhPuUTIkllBgasnnkNsVz0WKhlM
Qkdo4s4dgRr5oK71q8J7YR4bLc85MPVOjUC8Dt4RRqTtgF+zE/zC4GPzAnKp9VMx/rDzy5mGK3i7
efyOJ4aCb47dishIzzQtdnVh+9foI8PdhQX7G81jch6zJFcEYO2vl82dvrA46nX4SYL2GW7/odYA
JbWg7HRLezhKx6wN6MA6TE7aXyZeM5PQxmxZbYJSoGR9zQRFJzR8ujWc58E1QoQYxPIQpjRfJ/65
73veHtQjkGZTzdsSMqa1Y254JVowyVlpWgiYhuJ+oKD0bHRDjEC48Ggj89mDcNks8Q5nNXg+naSt
sK4ufOwHLMa5yG75Yrsza2CVPIBbw0UXmdRB0m/9LQp5K1FJNaZXpg+8NTzqu+1wTRyJ1FHYfPb3
Wsiex3w5ApdqTZEdqXt51lBytjQPM7I+ls6CB6u3OGkaGwklBx+QrdPYJ5FYU4xwziB6Ijlmrgvu
wIP3LgZYfugNzVEF+DP/GsW9VUTD4rO3ieXBMP/ItrL3qCAg3oouZVYEAe1X35dMdrB+lWrKa6pv
8uZcIi9oO5hAE2adP1tVBy/p6PZvOKqBeXI7bdCifptVPD4gooV9Oiw9qZpkywrDytjVO9tSRhvG
WO6RRnhkAcdiXg9LjKlD6zDJuCfCOkzlvswKOyD5ZXstVfkct+jbFyLetj5whVFEPlmfvJmY/I0G
SNkYjnwAJIMlVX9TQIorSTCB5stZ9dcQ2V6ZBndQ92PTf74Jzi2WK5+Wxn/2e8i7bvNap85vxWmM
GX7SG1F9Ml1/dSHRo6yX/qzrOWjH+udhusB3klNTnRirL2y93l0GFXGWaXsxxLDnctZ3gpT2UNsj
ecAmpKDgLXNS6s1/zsPL2O3R83qINZHTp6jr3MPFX6fk9NA4hT82pHUIV7Gs8q7QYVUScewr+ulL
UdP82kNia/bBuB6mMxwIrPWV/U//q2f1XCn1Dp/yQ+W+cvuAUKbAo8ZX0wM1WRDqrZWehYwySyTn
7wgnPuyzVw48rTtAV44dV7J1whJdT5K7GMP8M/SGpgOLS2/dQALd4vYv2d29tUtvHuQzfWtm1veL
EuRIl+6qd4FtX4SEKUuZwV02XbIfNnWD94LaGxD2QaBTm3YX5/JjpUq4HoKJwrwY1topc4cxlX8k
ux8q5GrGArUAkH0uUdGlEuPKnnfcnfuIPeyS9ensFoexAr4CAKSSwpENO2vjxFDImOApoxnj9Zhs
Q/FEHWP1HeGK9InFG9ygZvtjuWnY2hM2zRJ6ubRKRJVWRrNzgOQyCXyw4IlSd/FaH5XsByJ1L0Ki
Ki5zXuVKwYzOcxoQdh2ZL5uygns8ljiQ9MdhJWz6HKlbSNz8SU0ebHKE2ZuaKtfxRunPETQ5ktCe
Y9qXXita6S1/Ckz7K8dVZ/ppgnRMavulOutT3w5FoE7IWPvB6JjwqdmyjQZUH8PS4pNTdAC/5NNk
AGo0UZcafREHPiFsFpr3nlAboCU5hUbk8h+9LC+3cHfdmy45y9jvbfv66kHWvxhfDGr4NBKx4gaS
GGhNiU3VAdNgkEc00ILW4TGQwXq/zZ8bnJmpgLSAx7pGtb8O5L2J+wYHw2Dlj7DPNZ9QgcJ0lXBa
qzb+FHYmKM74INYcgzpO1DXQ2peM9g2TBZ8+30fyJWidCI6vMA0wZAgJnCSyblsXpau4VaW99j5d
JT6oISDoxO+pZX5RBa0D6ysiYkZVpdIEW9XBl/NWZC2j1f2xVJqp69Pd2yt3NF6o8naGmi9gFCuU
JWInRTeMx3rs/z7yKGlKQfBCmpH/ncD4YyTonFlfOTUHyHkVwapB9a6+5S2Tx+sIYIxs3Qq1GkTU
heBklY8TsrOXi3gLLj1rjbm1PiePWhMIAgtN1V8m9+3xCt99nYr66NWhDhGu3g3pgpi4LQfgV46O
kEXEeRrOZV4UQIHqXUafKB/H/KW2jvt3G6G/lnRNUQFHOd+K/ihPkZ+tUtzZVdpZHW8VxQPvlATt
lqLEAP5gQoGkOvWIqxeNxpOglgFag3gXVxgDNut7HJtjAdagAztsP7TYEOxlUWoVXejK9ppPD8Lu
llLUdOT8IM8tKTQGnU1DCKJkUETANqsvBQrUYZ1+C5P0OpdhjM+3Md2loqktEsQvBEBuB+63CnDf
GuDWyldRxFRdy8ZUXodrd584uUs3zpCV8Efh5eN3vtQ4qHKI2w7FkkZSTi+KcDqkcwnjBZC9ZgLB
lcUBI34/A9mvIoRjGuvM3vQFreEAgJtxpX0J4Yz0Ko8po27jJmdHpmghygWy5j6ADASmbhkgfaUZ
Jydou46yOhjK73qtRpsqZ0h0wKU9+agjQWniMTUo49tevix6Vukbw47yqMI76ERrZLd0nKHO31jZ
ZD+Cg3f1Jf0AX+bix0ejaIOiZpB/iyhmD9EDzx6QxPrFBWvQfvQOn6Wbl1USj2s9q+4r47jAVaRN
FhzNqEvE8mVG/hjdkHNJX8Hy6FnvRZxTHLrAY+0qrU/ThVSZjVz4/rIkNnPRsQsSGLNeSFDwEEjz
IXtHHbtfWU+Y1wpSMKgypVxvBqyWxnVTNtDShPn3/dDFqyWJRP5GTUe9DMyiQsanO3yfDBDfwVGg
U5iJAcPbYWfUlp9Mn105euNm0Yej4LBrvwrdmDdRCms23+kg7zWNak5rosEJtsUCA6DM8hsJJvq6
W9mydG+jeA+aapcW6KtjwM+fcXmmRuehebhOUBiS7vSPDcweNQ2ys2fHg7CU8EU14PhYAjgOpZDO
BIGOyIUBFULB9Ve/ADe6tPeJ7L5gGzCyDg3GUo/+Kgu9zm/NqMVz51hvxtCRd7+ZS4oCEopltukp
4SG5r6kZwqFnKY5vQzKxyQwvQEgEauXuncJ6nXlaiUTV4EcAxj+04Hrx0rJQC4Wt2SMu8r8tTzRz
/m3j6xLK7XRYxPNAIUQbI2lO45AA4UCS5clRsvY4HgKLL9uzOzX7zeRdXGowzhgoEQ480rLSqXQA
shKz2wp52znDjjs5/8qt64ZWFK2oOeWWsKNm0UqEqxNalaLVTGcGoyA7atq6bY1yWWuQLOY0lEkN
7VR8N+lsei+/nN2GySyIksBHY+34AzIHevqOlx3r8qIbzfDjC2jAzYR2fJ78RkvAYQaUOlfMjUPs
zRk2st6WsS+5R+ZZJMay7CViD099GErFmsxVnmiXSh76fIF//AMzOwuATeROkK9uSiyRyhYUQFwo
1OWlwVTTZvSvAzBeZR6e9ejNJM5sriSzJB0r7tM0eVcPegmzAiZqS4EEEe+CfKhjP3raAteUQ8Uy
aiUK7Rx0WvB7FO9OTEOjOQhs2LTjYGOw4S8eTEUkP+xr4QAkGFk6IH1Sj+sf3UcTdZN27X7lwIKe
pOLLpr5qx2S2LXe9EHwoCsa1YnPedxjnfn5CU1ZIN2CgI47oQby8VliqqaWk+NY3C+KU2Tb1KYUB
tIKRJvne4pcfj1MOYKrKuVGD2mDc6WRR004GOpQsYfDfb/wWtfHqF5qEEVMAHlK0rFfnYjixaf+l
llzGIsgblFR6WnHth5kgmJrK8T7Nf/RhQMmoW93KiqslfuVLu80ooHLUV7qSBnOdWWEnz8t2oTXM
jx7UoQ7o87IfRBHGTx+oiGw8IrplePwL9MZAalw1fHFnQnjd1cs/RhrIGZxIuP33o9lRKx2Oa+T0
LPW5gi0GDir2f4sCCVvhJMJvgWL0TM9fsl/S4IxmhxN1dIDlnFr+MFmf1uWDngPwmVagMS4ac/t2
JkTRXLzodKr+onhADlqC8i3xWDL48ZwdyflpuNBx7aN0U5P6VTpwhVZaAN6IpbgtlCrZ+bpa06sW
dD2XoCchkNzYd9GhYxJXmuRiKO3VrxLOZkr1EYmvq8O1bFn+UFEPUtKyjmwoz5UbuwceLTsEq5/c
+HkEZ7xEVrxRyROyIzlJStWtCK+Ib6TXJWwqCzi2uyQkifjA9Uuvtyy+Sk0c5jS8NwbFRhE+5ioy
nLkWIACvoLsLXcy37YnAteyJi1ACQ2Om62TuYSguD9RMk9QD7AauKgweFF3Ny7d3r0eue/x2PHqV
PiFw53vwMqvorY78Iq/yzzFhI67tLJpfv2tjFg+E96+Hg+ApCMyQiS/mXlsMvvWAGaDFGHigQuRI
BUXxbcIzSAwQxY3bCdO/hdeHx6BRARXCm8JjHBRE7Ji3ecUjho+V+wf9JlJ9QIc34RXxDAap+Gyr
UrFPEW/GBUm7v7IhHiWykUSiy61A5KQEPxyLiDrxtV9K9djybYkLMUXHITjvliAli6rke6weGe1s
SYSo+fm+2zbWHEfWffJJN7gJii4BTYIJ6cYZB5o1o8u49c65W7XlZGUCQlBAqROVKVNTBO8wuqYZ
HAr/WOHq7kJM3X2OuzK/tkYuzTI8S0y7Ic/dpI4fKzDPNZSwvVLLfYnol8T/F1Wgtc4cwJpg3l9R
po2JVY2fcxr8xMpLkN0CqvNspGMfsUgl+A3kYmbCtFNo5pvza222CvonyieKt0zNxE90IuD+CD4r
M57Xu2HvLCm7N+KxBVRKW7c86Hw2OgLlReNE2LXnCHb9ql53SYvAjHExouQYFAD3oOQ371KwPF3w
YzeXhrac7dKGixLLYLGnZiGtv+LSypz4GwVR/QM7GfT+KVrJwkcWzLQ0zb89aQBW1ZnPpha+XLQ8
2UB7cU9U0KeFcbADIpSaTqoMbm4hVP5x5nbXVw9j2lSvyfFyBtrBArX8WQ18oyQNC7RoV02qMnYV
RayFMsydv7tjrLHkEnlTm9gMmdHeHGIvPbAbx8moSZJyhccH7d3bcAIlcDLuYS32WXlxZBW12T8r
EMtE1DWjKK8f1cRZR4PXtYO1LX54C/9FvWK1nK/L7WSQXPCqOnN50ujmGRl4rWZf6xJa4Cnd5v7w
JugKiO9VhzU6Je1L9BZZJeclBWhVqEq5ByeNFXIKrNsdYzTpCfQ/ryfm0rBMszxjhnuEFHXWzDdK
GJhpoBlg4C9GrIW/sdf8tF4hRcESfy78aNwod6hwvpcdrDZuwzh8k9BcH2jZkhXYTLuPQJF4VEXY
2DMFfQDBjEELZXd4dCNcdgCRQhrKHtvXwO1mBgZXxjaYjGLELaxPibjRX/7KfU/AbwdxIC4xc/Gb
wN+YPiOcqWCGOi/ppcNazdDaoymJQRdvzwb6PgG/u8LPGiQhQpVaxbf8TuB6jO8pJkfxvy6iz7CX
R8TAHoy7R/TGlajpsIFqJz8imWLvk98WhbeN0Mber0nLWDOIM5K2FSnRm0g8/WhYIob2bIMZQ72y
mlnn+m3OZLI8025ajFuQl7IR1KrTIuB1uOBBcH0MGahGdatJnc5vKRIrZOZkxnXQ3HAjXqeKB/F1
L4gEGqAImPbLUzE0LOxIDG9Vb2RaHwHieVdvoUg1Wl+MUgktuxRdzJ5r1G1qNDqAZ7yvqI1rvmPq
3YcGKujZfRktkd4ArnRgoPQoANKLIm4dLn6X5+5VdNhW2urtpaSE3ygzkZZprHDi/v38w2IYQpJB
fEwadchpgplD9rQKQZw9ECuQy0+fLF/AoZzsobEL3kewudPhErKgw4a+97BuE8GLNpLPuHafX3WF
qqikaxgCnKx0Zol4eWHyU5Swl06KV91j4T41NrEQWoH+GJeXeKKs5dUodayKy/sXetSB3pMtziCc
qLo0fU//uJUGOxchFmCGXtQr9kVYPOwu23BwlB8XDujkJ7zph7jmM7rCG728HDz65+DZ68tfgkb0
BXcYy1yJQdu6Mm4KwMj8vYCiZMZsLQINJty5OicTn5gtC9enIk8fyUF4vjWKIXxkII+tLcSpYK1M
Kc1WxiC9Jfp+aIZxxmPzwLyIMKcZ2GpR5XNj9mmv2Hxrr+0eNtEMPmDuFaIDxzNqyB1rDd+F6rtG
/MzHmY9EtjSL0WEAkNMS/oxGDjDKu+A+8hNz0lbj0biEPthVTkf4hbykaSWbgwVyLvle2dsu2Q+m
pM/hj69angZniGYulsPsj2p7jeiS3MBiwqVH0PkizCUSBAON/r3VozlH+7xdqHJo4o6UCEWee9ld
bjmGf/EpCorq/RyAolyj/pu9Q0SmVLIBmUgSoyQsCUGFj7AS/6aum/0mYNRu5Cwy7eEEWHaxZH6Y
tygUMz7rzAxAqQTi9Hpl7IMmEs0mHtsuy/CuyxB8Wm0HHrQZeC/1DQx7J/dPoX47iblF0nRsTAmx
T8fy8c5/o6yhCof8Tid9SWH/rOzzrBzlvbQDcaevhP1AYDgNLfxKAkQr9KyMrkO5UAZbY9f+z5NE
iKXup5uTBJvLze255jZrEV40YSWQNcj3+aPUyW7pXBRJwt+Bkj1sm3HEAQ70KLmd/ldHdRwNioki
ghz8eo/PWhU/gW2m8mTST1iMUB1PpJp3W98YpyoCXp3TV05xH+2YSXhKCZmsGg5QG4RL8IC+yB+o
He+BDjy1Rxvg/ouQSrRnbAKxVZuAsXGav852YaGB8nfcuzy77LgYV6HlAHyZkB5w53R/zb6Zd4tX
vW0Z35U9ox1BLvrIbx13p3BTCAkAQ8IqbWD+PnCTLrKG53veQEfAlUOlj4q4zci1zSwpTX72Akur
s2Lren5lQHxSyXwiwXB6l6ufggeNW/F0th5dlKSmsEqtlQ1MZY9FvZRf2LpFqopmeZtDynGiR/Ql
ZhYsYRalfXSB3jTw91tiaTXQ1JCySNr8fOBt/99/kQYt8jFWAol6X4JJExlgBn0yswwUY58zxm3y
lZcsdM8M6R1vFPc7DIl/e83a1KoxTvCk/ry2jBqHzfvps6yb66FlV9ZJUquX6hP+r1ZfpzrqzSV9
PNzZtv14djLINF6sytfTPA1TJ6+fmTaCshiZ6jLgTlij/dvz+3JVj2GDV0jRRjvbuIbSIC1Uy+r8
AOyT906D5RtPlSoedrOH0W0iE5xmLw23RYFurqnOs7B9yIunC1nW1GTUUZQg8GmEhyARFj5xkEUd
ablK6uv2FGLI0/uOb2C0goj0gykGRYo0OLD0mhjkNUINfJYyPIBP653b+MHbNHgFZj7bcQTugty+
oUjDs7lomSJxjY3xQ+Sjn6l3DH9w2RFYKt6jElVR3SWQ3C6kb1w5e22X9JOhCS+TVtSAmen2wr94
Mttl35ZpZZeWJSwDaPBMOAdqQ65QWgfRkBUivXGSmBSNxf3MEq2vNIPRnVOHBGO9RgcTgRlH4hQl
1YAdNuK6J1z3JsQmui5J6oo+/J6vUw+HVe7KP0m7LOuTORtbLVQOjNWrGDM8POfgX+0RKq6tMjrD
hfL4AH5mA0L5LlGiPaF6L8/6v8jaOaRB8x38pGw1MtRxrRiT1VSax/gtsTeFZBOfftBP9UWPrhI9
9+RH8HD4kT3vIzEu2qce4mt8LBAYzi2yLlIzE49MRlnbIm1R4udFFWe6j24qBtX+RF8ApU0a2p0G
VT2tgsKmU0IUI2KHS6mB9SyVY2yAWMtsKs5O5f2BTkSk5dncoYxZ4PCwNg9wpeI7tJR6uAeMtPov
hjoDE0xZPW21LHt4o2xaRBsqiGsnpyUjuAhzwVJSZu0AxhVd3pNJaGx1eifUr19h5ZxZJhO7D9Jd
1n7NTbbWw1xXZYpw7XTn/FaOOVanb1WWkkLX0bWbkucJ3HCPOoQlGGwlgTPfICR29aap1cgkMvgD
Uo8bd08Ya2v2H5f8OgLb5hFc0f28iu96Lh9pPCj9bCAXzSgjFZOvIVmF9ZlmgVqbuakfmI50oqjS
U1+z3naR8PcELQT5GYpUjF8rlyE5Phutzw6c9f6iEUXKKhrXYzp0Q14CgXWafN/V338awaQlWMVs
ao2XDbPU7wGxqdB6DgBKSj2yV6kds/j7eZvh85WsPsKf8MrIcq0RD5X2WDmKgT4zyNGFONjAErxS
DDTaDPXaNqfJKsso/k49fMkpPgyftA5DknyAVNQ4Z2QnP0pAS54tkzSfmxukKCiMnrmQ6/DQPAan
8NG4hbS7I5isfVViOWk5rQdKSlqfD0M+BhZpKszaJjlu1EPju2lcwkBaNbtjvYtnOql9hpPkkHVh
RJ+/ieuFwwNXn91B9lLV0lg1u4lzkj9mNGVsG3O8zMaqBTaqSKQrv2cLqNFSEs6efscE3j8MsBKv
1b+10P/39yDRK2M+rYxXRMa9omYH6jkhyTWpvFHh+KdAXTHeiKX4D8a3c1Q8N87JgrsfDnTOp/pr
JYSc7AvwK3Wxl3LKG6YXUP4umZjx9u9l/7Qfgn7Q90EuwDvf/2LDNsg+oZFNRvk/X6wEmDloa7CW
9QsdELhaC9522weonZm4z/vJccPYBPZIShiGP27OICG4O6a8FGQuHWXdCaaaW98DFRYhNgW5ThxN
VAXnArp1QPzR6Y5qDQUHuIWSdt5yMJCRaXah4XYGuKeVdGM9bMzDbgXHhv/s4xNepA8VuDs6SrQO
hafOdcOe4RswWpS9Td6LyBKue3YQrSKIZ8ANk2nzomJQ51rKahWslEhNhl1RnoPdcdhatY0UOn2L
7W0B5qWxck0XjxOaMmlBEiJaj1bWbvOD/QPsl5K79gcfIiPNkucWZ+Pctf/Yb3gtJonJe2i6Sf3I
u1DaID2qefnlv4s915HXxO5yZJt6sf4kwf1A5KenjrkSjnlIiXG7oMkSuQg0g9dv1XDByZVBJ/xM
gkWEvntVvROPlJr6AYGwZYbt50tOipIHP22QxTs+rnWrmbIUfiRwVimkRtY87QuG/ShPC2SEfrcG
IVVagHsXqCFQiQb3w6LbHqfmViLOydS6rjBY7z288P+YMMhMfLNggSBzkkTxssp8QqxgZ6uiLlb1
6UhNkERDetPeXoOzlsPzmRURlyPHEL3K+kItyj20WNg/6uc43cHjeGxX2JAXO3MPvNZYsrxPcar4
Ldz5Oeb2Gv6eIGzJ30IuWoFZm8D2V4V95XsO3jlgERCZMXF06ryt4InEJuu6kYfuABr5r48fobxe
R5dKjVkRIUyWu7sxdg2bIYUUyATo40aaoLHikXcWJaNikQI98XoAa/gENgBWGMWT15Blidh0o3cL
QTIyyvVY0NaAWMDvCQvcgo/2K8AXJDf6FJbZTXJ5/1RMdg8WYcvsNbryfOMX4ga3PeLhHKTrg24+
lsCS4mIrJEn+yjL/t2fa8ja6fA87wTdZ2mfVGX4lkTqNyt5eshl6CxwyepIl+BRmbur/FteUXsiG
ICQudZR2ZQpScz58WFePC4GYJQjSGwIxM/f4Dl3A+TGv/uXpp/Dlo/N+R6/CGCQFrvXHg+jXzH7y
/Mu8O5s+Dg1RjYwQ3dU4SzI1JFCcsLY2/eye48/sMn31ybtALpLO9I3OFVJFXZBk0pOgPSy+xuYw
ytT4ioTbp0htYqCXY0wlccG8P+R8nkOATt5WrBVJ7T11Hw2Ybyuisl0BMV4oj8WWKjoXo2zwLKl7
D3+ymjFnlZfX8Vf0hBJ/7SgP4juuBAucQteGrZTtOR3bAfloziX3AhZjSOGPq7FNm5dLPvk86im9
eoYAkNfUSK9EXSLbO9Y4UP7L4hkxg77Rr14OTk9c9S5JbPld2qn0SG/Mu1m/7XLYLxreEZlaYAnY
ZYnuxnG8wDPpnfYDzobqlnWqWUmUQ2VxZ0In9ZdXw4QPnCQ8U+mhTzFmZy7eFWVwbawGidtbQBAn
uhHrtCxPvsfSJNbqxIBuRkI/otUr2agKBTiiE+cgVO56Bt/niAitbz7Un+rKLiANlvShAoN0F3Gw
1dSOu5V9lFcfYefy0xFCYU+dqCCVC8U7y3m6CHfYSBfUGQpAueR2vJgx+uayGGK6KXS5bglHNTP6
sH6swQiyfRLeUK4v/NIONeBBWwUeGbFPxtljjDRebCEJpVCaRhpeVdz2YtQgKazWkH6yMdhTxG5b
k7Vof/oWZMli1j/Xa9FS1j3vJXr0p9t7Mue3Ow58m4hMtg86BFNYXu4f6LSCZ4YxvBNb8fcZBZRU
vHIia84XyLirBLBAlu+6voxNNvSKLTVXX2xZBQszw+/8C8Ke1sSdKLgRdCluDpuXhsKF+e2mT4OP
913QHMVUSBhIlFCj60E2GU3tDX9IuAn2QMolFdMJXQxspVmTsmTxpWygE4l1gIuFhWrv7kIknDwm
BA9wmu5x4N0IKyqUjbFvb2Ykx7i6cYAkUlwNfDNoq68AJ5/KMlbwLxqq+JV102xejSEczJpvJqWd
8zLvpoiXvQG05/0245YMSgY4EdVqSBWnhA/ulByyIloyPTgx0yEos7DuviBLFlMWiLcyIqC3C7/i
zkUjGBUUF+SghAuzY5ihL9pcgTgDnBXq9LpqYi9PaQqMUGXDDgkfbh3eLU8n1LHxI5Hf8WjI78by
3Upd8JHI2KPnKgWRrKJLu9KstGsZO0OA1UdE38l2iu5C0BSqd7uQ/Or3dKiEjhyOQ2RQHCJ1gutZ
DA1kEM9fIaWR+tqSfTqau86sI0Ltbe39hHyn5WcCH5iJgkqsHw3cHIQ+KpbWO139Nv6wjsNRh4If
4YwXQsM0JGbQgZt0EnvefHTcpJXpW4qO9CDoEU6RfgXxvLGHA9GIiKBTG401SkArrwLct9JPfoEu
0ISu9KPTEzTPdRW0YYa+7fSAFtg9gPL82KCWpplw1XCowTniGgNGee0kNIiTjawFie/DgzODLiz0
xcIvBUznQOp2773ExOQUNBz+Nz0ZfGtLZjVHCqn7zaW02rHSNwR05FhUOTjIiLDH8aNV5MlaJnG0
kcNmkJq563AYo3x0XFsKay/58vgj14iJF/47Zz1GY04h6NmhpO7/VR2V+R4DEHpG0GG28NoF+Sd8
JkJjEaOKAEn13aGv86bKAppI9F+2a0s4ZXk8wN9sz7pfVncsWldUzZ/qi8HrVwiy2GlNhfcDwD8b
eiV+EseQHLfkDgnWpeJC9dv5o9/qKjZc3yVYSj7PD1zRTuefJuz6GAIV10pGiMhenuYGwZSWqS1S
NQ/tzd/ZIJOfvLw2DoMBOHRHZK2qhavnYsHbBuunE027xN+pGp+BAtwT45y5C4q3/wbCHUlzBuVW
HXMqZiGJZ/E+efC3FwUFeIqIwamKDcCRjrezMUTDAlqvfMTZYtCVWSrLYHsZBhWWQdS4cjZlr10c
Q18ID5fv0bRhBoDDvu0sbNr3wG+DA6NhE8K0TVDXcMpeydnQu2amnp2pg3ZQOLBa0zhOxy3F+gpK
2B7iCOdvxpiydHSHofKvu5/hLrw3mG+n6NUh7j2bdXTpF1l0P7mDSyA9g5qrdZqedYJTnTGkSvih
A6sZWbGkDE2HF6CGkmzc2c4ZXXQMa+Rixkdax+ZWYw3c3J4Yuq3I68vYZ+ter8hZ8tooY3pBBVpx
N/ucRwte6pZdVCnWi8ZbQVQYxKzltZxrkrBkUrHtZvBC7iX5wkOC5/O0RB4R+GItLxsqxNwRMqGd
AtfYURnpxRBy+HeZSPXt2HYJZSHzemCTNH7MzUuQznA3I1/awo1ceJ5B3V8zTTu21V6hkUz6PuBI
fRHbswXjU3sSPM+gEyN+6xvpjfZmUVS7Doglv6BK0miKlnRvJuiM9r3ufQSrBJHlWF9cruAntFTj
WoemUbtGZGyNOT0pefn4cJasXX0+Ex3RP/RDp+bJ12hBryw9u4JezDFU0tJjgv3eGRvz2lLv2J5c
P8QZivraVLm1n/hey+2t+L9UdbKR/aAqyNM9DBpdwdmEgR3Cf+eX8ph3u32bPuycF34RjoaKovIf
FSP1+XHBI5EAH9gT9Z12pVorUt21pdsoZfAazcebvjDTzyyaAyfzs6Up6RyEfm+iOsDM8YSQq7AF
ShncT9xySMgAkR1ZGgC4InuiCUPfRHKStTpU2WTKFoO0TjaTcgf71kVqjhO4feWFss8GIoW9hFtV
FVExuvwBrxW8HecaIp+nMj2ZoUuXAxABW0IvvJcfE3jUDznytx1E1FjnxXA3swycdafCZGNT306c
59lPhfaT3kwwj/peeFY5J7OAmyzXefflDKXk30ZbqskapNza/0SO6OzPHMtnCl9sDouAy+IYmKZc
lFeWPFlK9Em5md6Dm6X5aYWQ0UG8LQ63s9LAp4ccDlhmO+JJAlpJTq9ynlPnEJfhNabcUTZR+u28
YEv6nCkRePdT9i10ef0yRp2zSl207KMPM5XYVUAPX2Iy+RoHkrhojhNmrCXNKVSjjiUEmjUCPkvV
ygxh1HjQ1CCNsmYjkUEF70PD9ukK2y7Ky601uyMiiWgNI/IB25lr6YNPW0FYMCB/aEFtiA/nRuu3
e8S5mY9asA3Au8C8x5eIMzKQwqplC1EXww683XIbefVuWJ+WwIJHEcVLphuFno9jaAwWX7FRxBCg
zBgjjw08ceU2OrWL51vOUFgcYB4T87w/LQHj+a0Hu6mmBZ7ufSZ6eneHeT/zuWgs9eD0YQaNwrQm
tZOuZrJv5ntbpZ20xYfM17f3aUHht58Fm07lOZQoIp521Z0ZRvG3VOKpcfIy9yE1bqk5166mS3cm
l/s9kDpuMIcp+KsNe48PVYVo8w8hb71XL1BUNjgg5gQQkuP1QywICbd0RNY/dBHqdIpdip+hHgjq
C1uZMHM5okvrPsC1i11vaYOX0S8JES2qgI6xZiCH/zy3yPb3Qm4PZXMK7LqTtNpTf1tDJWVy2XkT
X2kaxhPMPprFkLS1HOdpjiPwOp6HJTFvp1qPN9293Mpv2hYr6xoonYIUHAii7QmKjG95rYPhMskB
PVmsYdZwuwLV/70Y0a+AjRbWAcVYCEo5HipllH0/NgyJjzyILmouTIpAv91DFtuyKqzy4SEF6b+p
nqVz40mHytYIMKxf0MxGNtrlxan64B1G3kbem0Mtv4UaVqrnn80kShSJCTf8edhz51RPazH1kwHJ
Q2cSnqyXU5N06tv+RL9bs9pIupvyW50g7RT5ALb+Y6Y/T7vmEyfB/rAB+kuFwefWYXSp+Z+vHqqR
EiZ6sFaI1FL2teeNHlYErPBcAWm///QMf8sspEiCHG8HjtCQcHFmiKmgGw56g/XTcMd3jaesQnld
9lIXBAzk5JSG79DmmYG6jlTBfZyQ2o62xDqwRssa3aqgKfn3oSJ5+RVgO5+1jmRnJ3laSjEUyX3M
vGSGObczR7nUaxZSqQDlgmqyFzG8qqxrt+ONtK2spULWDXdC29jC0JlFmAFZ7eO28jz+r52Qbc74
4TLJZrhfRKczBIh2pfou6hMMMyhQyL3ohjgSXS3Lg2FeUVp7pM9gNQxV+60ZmEg1xicdhA/nhgye
WK5Yu0obCWBntXLO5bjY0jEmqcO6nCngCJci6i6XMJKGRXHT1GVlC9d3hTD+rH9exSHR17/48pUY
U4vF1jRhHmHwLpkC90kV18sNb064Ubt7gUtWSFnyfr+ZiihtafpPGaD1Hqd8eI9SFM1p8TESCC4l
wnxUNiC8rJWQb052VAPZO6tKJg0t9FAB+A3ARfgOnZu6pUth9mpVLbrbqP3RKzKvVJfD0fkOyXBw
cjv+MbfgpZ+jHj268VQzE44cSLWjIXksMcOrcKNC7TXPT3U/zjexq4mL3M4Up81L1WZ1SxdzBlUF
pF4TsxBdG/gIAFTufFxAdWTqK01i4a3ebjtk0He1k5W3rOZbfMG3P+3QCv1pc8MC0R8gN2hbUbgf
RE343YviefQHvVtS0fhGcM04dUcL98vpPbBXYirWLhPCK7wnBtKXWLfNJ9XudBF09Nl+Nj1XV/SB
9XgQ+o9srDnqtKGZw7S2/nVhomVJzbtNBq7Ro1KSvf9QsuXnCEYYX0MbJRdJNZuVX1shpVoiJezd
rw2V68PaHpVO7xlElxY47FiGYHG1GDHcWlhTF1iLBdZ17RtNvo2RW7f0yeJaDsNfknNrcoKy8w7f
Cfgg3/Jc96CU6AemqA6nf1xNeGje2ELt0Y6wCt8cwviyTAKfIKDen4CqCVYIRIAejffScLWybKcc
9HQGXfbw/cvooeGqIQ0CAlkO6+xnGWt9w0NoBB02QIgLI8S8xoF0uptO169xDHhf/R/IjOjDzTLT
+FXzXQIz/MSdDCheauxxrt4bZg6aCJttrxVOn/yKBz6Fzsi0rHlyBbsaxKB68/DVLNldSU4eS7Xk
r4CrseeGPklSbz8KWW3gaQXeRSilheQdjBMj86G9ibmX0PLYytBD+/Whv5X/SoUJUV8xnempEM/G
J8K4FtXxrMc6JaEDtYp7AHNm9CSf5I3a2LCAdnWUKyVLSvyXXphs/WzG5caixiKQiL0Gski9l3Ut
KRJBBxzOJiILpPjsxDbiMY9oqXdKw5/09mr5jES07ktgM/A55HCXG/vRuMmq2JqwqKzA403a0E0q
hYgXzQzfoPuSdqTFPrXrxemSiCxwXA9ePxCGa9F81BQBv+X76kKAiuf8sxg1yMBhTOtswgRhmDs8
c8lyWjfbHNgjGJQfuqJQZ1w1/T+Eh6c/d+rBjiBkbsRM/sgvCD/m65uXHChRAj/T34tFUjLQEtpi
8m1DFBSsU1xg4uEmQHWNzIeYfXEWWCsMQ4f/SjcTOaq9BkP8lyNk1ouAqqIY5up6M5QrD+9/dlec
vzLFu5waJiwI5Y6B3rdKoVvyuNf5COwei+PRxgr0WAendBfyEaXHnKxQKmuxu4Lmp9YyxU7w9nSG
scmFc8DDtgmxT4AccHqj22rqPaFM392OPM+4EeiqsBHzeOBrhrENWX7uwbrltttVIuFSVDnb5+oN
FVCMhCO97rNkQ0rO1Ku/yq248F4GIUT7GUJ06Hhsz2YfYicurjp2aFcRmsxuimp1wkzE6ovHiAcO
Tz/oqbEoNcP1ZiUZkNDU0Vx75sndj+iH/LjoAkHB7a6iZm2oATcumpOTpasN9pOWzsyc25XIkwFE
cFPVOxt9yeeTLYeVP34WxYcuzfrr0Ro34s93THQOEhoXMJVd1j/ynETsQ2Wgj5SzwVZEOeF5kyre
Zh5+6wxtX/kzVp73y3lnNtTEBzre0MW2M3fGj4xr4/W/6dEjifFUp8zLkp7zRQkbNXQGDE6j6h4o
Yjl9rBKcOJCmeBeNAsegYv9JlYGlp1Rbtpl2c9pGKT9yNhZPCEQvGk/wAZOpChuhbKrDs5s03QHQ
XpsEhyU2zDm77HGQ+ga/BW4ds6bRtE5uCpzJU4Z8Nk0xadsc2qJKvPo+sOcMWrVF6YmUCvzNXaBP
IAfCvm4Hfx7XHwFtRR1AtOkSuzZe610OUloQkE8abcoxST/tTT4fm58OhGpTVGfyr4tMEhF+zUK+
1XYQw6f2U4n4E80mbmEBUMzzYTsZtPcsssKaZULhAki+qW6ED8NST0Xs8Xj4jHJMm1j7MFi2OWM0
8sPa6tjJs/+efCuvj/NYzESO0KU91TzOrtTgXvdn3mU4Y0Q6cIFyob/WVIYdmbef59MAAvqWoZd/
QW/yxgHKXXiIGXG8R+YSC71grswRrsWaJpWtg97+k6h70tQReBFj3CZeY25ULZ+sMBVaVJpWmO55
FIx8LGEz1+1zyASkcZLTK9ufJf5O2Q7NF9oNTEjMujkEh3e2kEREz8uE6ds3Oy9Er6MfPTabkAel
LInxMGOqymJFlA8hBdFrc8yTmxcH5SCxLtvvbe+Uc7MNDpKUmBU+PVWf9IX86iABsQF3e7SZ8VGJ
Og9WkqAqwR/hZjAqWgH5fhOSvoy3caPe/+l2Hzka1DLGYYK7zRfQyKViKZ12VU52jMOjtTAVnHlL
xaPjhoA8Nsy9sN2CxF3mloNJDU2lRlS069w7Mp93epBxU3Ew7ZT4LucNTmRcfEv1OWR6n1+H9ij8
clj+cILxI/KO9jVphe1SMM5yfctrhBnUJD+TKKLw4qsR8XcnE1lo71gyGmVDHzV+jHL5+yLKj5KS
nPIDEOzx5qjZ+RQyZeXHsAcnwCNGgf4SdRoz4DoB+zc4zzN6JQAKPg0LJBVJkIV/eqYjvRw81x9d
4Uxau4X82/33JnKXAZNADul2DJHvx/0gZ4cYZF6z3AGgo0fWPGmkcGj77EZ/nzernJyXvX4X2bP1
5MHeK6R/sGEOY9hRgUnSP45ABX8DzmwRE29mms42eJWIwRohkF6xOcj/X9ZrxY7XTu+K0VpFjY4N
WjADo3YIzGza7VF0qdmw8MnwDSmyXNMbbGEkxnKkKaimru+tjTsHRc/dRtbs3DiposFq6nDqvqLP
9F4i1TevfFLmlOWXEoIElkppA6FX02nvRCSlhsv8HCDuh7x+p/8dbL6Hknj3gqpVbx8V4fiZcs6G
5ny3PrKH+DMxj06HoNY9xMngdhb9RwCGllZSr04CYHQQbevEfi9x4SIjsz+VZPbL7wGP4QrnIvmM
GseqXeSoelAj1xAsrV5XLmvMVdbj3w1aM+1UhEkuMkBV9ek+sMmFxGOV5t3Tv/qUMfTf/owGnWD7
jWv11lcEtufwlhQACiNeepmlf+adaQ+K21dlc9wvRYrZ56X4y0sZWOvGhEJ/S/hofFEGIx3+mXcB
AByVLT61SSCOj62SGqQUpRzG+kq4+kdsx4ZgH6RSGS+6I+0AIhJB72TdQ/W+vrcf5Akgqzh+yBiG
LNIAnPWLa7lkRF3y4f5qgrqPBS4DMytvI1dkAvdxoFC65Tda6Oai5z9CxW8IoCVJaZ3g+1bf4Uh7
3UWt5bt5efQg4uzw++1xPyWMxK+O0V7sd6xKZrnDp5aQ/rKOFik/s9xglz/jIdqxDIzhdf/IhNgU
7aqwHHXx9+AGBgQgmO81UFLkCV6t2pN84ES7FG2PEUzfFd03qxcocnigNhnuMd/RWBpQjHlKadQT
TzizG6rzG9kIVipuxzLK6X5ZOdrfeMBNKU9u5JOVUqsfRDYwJdJsxKxUxBw+ah5E1KJnhvF3kMrq
DXwkFrNFPtqe3M0+xwHcYbB/Cjw9OQmXWFoLk7ICj8bMB36gQGn7UYa3iI5MkaJ50te271/X2XNY
xfx3v3O7T109drpyGptLe6LKsduElAYp6yTaoRWVd3Ra56U8wXdVR/VagTo+bVyL+aj20tmyVPSM
wshIOBy+lm7waxRXcbdL9dqY6UJS7z6a3RF4CUt4eGZvELFQBo9AcGD2i1AYGcA5JL2zYsSbY4I9
XDd5nw+CWFNhXkFoFZXGhH6qkC84A98yDquRoAWtlTL1HMMlIowu35fMVKXbqLwtF6uWgXYpfDoi
WOLkbwGwmrGdjDUGY5ngJ321ffztlaSq4Un0i0N40SnrOkQ0AlLAgS/Ogs/jzQYSvbqaDzKIPorW
PQW9ozlLxTPRf3m/CT4WDA6FqZhQYgd3cGT4ueCuW713pWVvOglWEkqAFQXvccQvnFvTJfJrRw/D
XApDVgr3oLu6cIncIy8lpMlTEZURleoHiDcgEGyXre2aA1qP0QfwPPD7D1zDlL8gjGtQx7Mt6DE7
k1HXiihzF4j0+RCxNgPG3svHb/xIkaej/GYTdIyr7m1oZbxDMXJwkFFysZTLC9T+HQbXyvbJW8Bv
h/hlaeHTPAz2iuQAbO6XCCj1i7N7T0mU+hpd23MkyPLMOwBj77jh4IaeG4uUqbNw/G1ohwQSF7+C
ge72Bfo9i0QWMUzvzSKerLxoQUCNHgoAH15pjv5VK2KXcsvKJTwfyfWtNN1Rw8gc9ni82PEI+FcK
luhreJEFIfdI7oUFa88TyOOLUNk9+uaMtVoIZPK6LjpMDBOcDYOdGcziiN1ntPJToCFl2KEBGyiV
D41zdBBNniis59Nvul9p1E9CFD3Ub3diuVoRu4awP31nVMAnKlcx+6nfZ2rVNeeCle9NpJzNCBhf
i2quM3DUIW5w1gA4BQ+uGwsV8nsBLdQZElo3d/GC9nHW/CDjcGDCI8xn06wM/JEkoZngRjmqsBzd
sVLWJ1keay0azHO+ugYIMHgm5DTJFkFOZW7KQpP88sjQo/jBtCARFIcbmjvZYD5GKYw7QDR9N9hN
f9/WPNGr8pJZJX0wQHIU3wFrR5bT5ndF1uz59kZO8HT89CCUdQhmQbQxWaPrVHAirWtO1/BQPkhS
CiWjKyzmddM8i26cUWpjgcHbNATSNupeuLJ8bWyZyXPwvrmFEIGyrDo6tGkyyKcxgU4g9vFRIsPw
NJWbWO9vn9Cw7Q1/DDHVI3dqYGtLnZzeQhLvCR/WUrn7Rp9Bh4AGjqNu6GRhKT+cd8s6GtDcgJg8
KgefvY5A1ax1ha/4/52Se1tCNyR93mmF2nYSpaP8xJ/67k/x2+7BltmVCjxfsXm0bg0wH02p6j2A
K+MKxXEV5uozT1fmr1mStr9KQP959B5tKq2Cvs3ROPh2xvUJOArC+3Y3wHqN7/FXrMuSi/kY/6nR
3nSOmWGITEemQDKUtwGXxEXfFhfuZyrHjLCMDOD44nI5ff9gK/vGZmRbw0EO79lFEUDI8hdeQzOs
UpT+mNKRgeZFVy1iAAB2uMWzdf+zVunuLmoVAuuw8KZItFcvn3kd26hMJI3uFjzrqzKWcEZE9l4x
NHW4yuMdKLQOw3qGt1DNO3kc+H8iqzyIyObPKnAWwzXRPfNsj+BKfZgIg51iLru+f6RFQDXwFCAt
i61nsqDNAO5IsQ/MJ8dqWXBfhFdcBJ+/Ug74NKx/EqWL5o1V0Acyec7s5uVWkO3aLo5/HdP/SuyT
8SNVD81h9SnbQN49dMeFu022+m/UskwAN0+qwhjJyIE6HDe1U2kiknwfuqtX96NXbeiuidCTvO7v
Aal7m4xWAHZ0Q+zI+hc3ZGWC1sVo4uJD1FgiO0SmUtnpsUmYC0tlBZ0B/cLiPeTv5rU/lQpt03Fg
R0G+hl1FA4JQRfGeg9M4rbuLlJPzcGa954rH9O3xh1nQgEe/uYvvvfRaozWFA0pmLyumsjeu8BQF
blNVRJ6EgIIef1i/H8maCkdJ+F5aE7WSrmhDADIqNW+sa5CJjNYafPnfXKTb7yQ9XN8LdRQ7x4Cx
8Yfn2M4wDBQHglv6hlIAOs8HRZ3vSbQcGUZQYbXvTVxthkzN8LsyNahjjpaqit2mfURiOkO4BDOe
Tm7459DD74o8vUMBk7s4wSewS4UOQ29TglB7VIiKhTnDD1yD7O01PNGN3I+mwbb+pOjRueMjAsGt
CbXFr4WQX60aEAVBHRXUGUfgGL4R549Ud9M0LOshZMDl2rPke387Yjy59EWL3kG+HyqHGkJyo2IV
wMW2LZ6XXdNpi6vcKUoormBq3JFedX+9nfD/gIlO1x1Ssi5TBeuQ2Sjm5DVRkWFqujV/c6MnlAOb
zvo4b5q0K/9BJZ/YDsHd+rfKR5/29ONsTMtcEKL+jBgOTa0UWh3uOaUGi/UznV1HMRmxchQlHl9l
zec2CyC2NLNQG9Q+M4LpwxJteItSVjbUi9YKZQ2/OEgKGz6ZXhHRUvYe4NwDG91PEfmSbKO7yJQO
nqVO9NJAGyxJvz1i0JQy63YJpN93m+kAeDSkLDUlt/okKzUNfXFePxhz3aSK8sP5hQci/RAFsRUw
pIl/aG8JRhQGvAlQs2PUJOYr99q3qlp74+dlozlZ4frHGqzanldzenRvYoRCwF47P/7FLE8Sq7oF
C/QZ/5hMJqrbMWXxcBUGbHjZHqHwl38ueXrOmg53669MHFYWRKYw1hBsPPnP3mGflGiMXxxLotCa
Qj1niSGPF2EQWS9X91jr6Wt0dwc5zTbO80nZ0d7OeHhKRKH7uKSPC6aHWgLY97alngeyKFQhjXQW
MJjw2dgtsTa9ZVAsk1GHMPuwO1EYb2S3AjPA59iEmNwMfVaAOlQaq70DymgDBt+EBxAhZs0UnCLL
YEN2KEsIvWgaObetpAw+GdnrLs2SvqQzJUDxCOn9vwViMaIJ2GzFOeW43PBwo566MNdMrpO6Nt0Q
Fq6gIPg8pFatFEd5BzDhy9xYVNB9tPRCsPRQDyYCpK+y5uScnbfTJgzTsY5V0PGIeUb5Rxvdmr1y
bfp6dAs8vjNmADglQF5bbIwOzp/X47+jJwBj8NLBqyVjbqjqy5bIJzE1uWQdw/T4f4NX0fIHcmup
zvT1uL3IfIjmhS8n9XGoizgUjxt7C4jz2JwxO79idsvHuj7ggNyFvdMI/87MRRjNESI1+gU0FPjr
gQXt7oOr+Z1RVn+KKY9GXKRbr4GkNbDq0AA8Zes0SwnoW0wXNH6/uKuTCikAwW5r6AX+bXuXdWMw
rkJNQTaL6+dKgS3mxtC752tWJMAv09Y+Y/yx8L8s2lg4L1MSnLozjDSAdpKRemexqYBo30witzQu
LJvus2dh/Azywoux7zisjui/5nLdKp2HFi4wvxOhtSRFm6POc+AGPSIyiaAhAzWPS3RIZMagWlRq
FWDU2DB1M1G9bgFOBk2hp2gW0lUE8H3DJlnxtWgz8Rde9jOvIfkJgUwOgoScGdaMfKnAOMweFA1U
BpEj904WbfNVqeyyGXouiCsmVKNW7OMWVD71FITUti1UWD6EL6Au9QLp5pTRU07JRZ9fbmp/tkTR
VImuO6BvZg/OtG4o5B8KFtOfDgPvv24SrRYLlrKyqZ22JBNZGPE/1kiPTn/Ij24jYoME9CkqWPvO
2FSVWaCiyrUvgOSrStanCC1WHYdatbt1DrdqrSKLYUMN/qkUt7f1ti7n0Ed99p94AUny8g0780MT
w8gKJaBHsweYT8BhCSMGowfFXXoWxjmA1iJskDVpIHPOw0wo8ArJwImw1PKeFkVA5DOZOLf0PEED
tFTGB9kDeA7U7FgeCZuIJS/VFLufa6VAPMNS9jBPTcZjH2q3DmriFXCfXs4jxbgRpArFm/81sjba
/fNGZiCrOWtPVe+TYj4+89jXZ9Kt3mSwtsI2W7e/J8lJtMXeXAQ+l7vDQqXg0k4iEj0YZ22hIwns
+PT+y6JQ5ojPWaGmkYc0VmPBL/yK0pGfcqJyU9B963FG8ksgwnqrtk6gK/XuvrWaruK68F7tHCXG
rnAE0BaTLyOgW04Rcmu7p/Al6hQ5JEt8LSPBGnAaJBipYuhkPHdlvweLRC4ziE8QepYHJ8lW4sYK
2xK0GwaO+7JMKADTjIoi4wmtn84kH9XeIsXshiYBCseaQstElVoIlquT03FOjlM6okgcVGfHunV8
dAFnlYBC82abIw4RbKcSOoo8QqQEK/49M838naEN3cfV/6Wm9Uya13XnomwVAmvmaFpg5yKnlXDr
jQ9cUIFGk2nYLu86fxbskfujD6iU3wR8qWuXReo/dPSWvqFCXzkBYdy/BGn53nTpJpIvMe1Hi51r
LVSlxnSAAtOtay5lN+0tWmZZMu6SSfMC8zm9eb7c91pApxCqbg5eNPeKumbCRiL4ZYCcqn9/BxtJ
cTmnJUmrRKB0vz2HxfpAJiYZKFX3OxMEqQ1woMMTGjxJIAJcirE5sFoy4/GJWjg8CIKRZeejBzJn
7NcAFj5vuIreYTyod8DefJcwkwykqkK46fSLPeyCZL8Ythn87tRzNpj/j+JjMj0MNcjeghdoGhrX
vTMm55IvKLpm6bf/ETd5MdUjoh7EzZktUjGc125lv/cAKRr6F2ts23OIEDxySse8P3pYQkCsTOQ+
GfC8aGuIYG5dCEApzbqHTx99n35wwv1NHDR/EZsBJiMRa45BeH9MuTjmt/npJKlpBwvOLl+rWqyN
ZCXJGEuezWCyFllWlYgLTG27BHopMQNzDrCGhhJW2TEgPJmvH6afAUpKWTPh6F+kFXXn8g0c39Cb
5bFCXc0O1csLqQCPHtv4RQ1KgsL4XqE5/dq5YT4cWnHS7joYCqn+yZnIpci3vuDQANkc41xLVGfy
vueM7mKJajG3c37r8VKugY+SY1/6GoWoFoBjYR/kbm/IbY9nnOVGNZDtfohDJIjN8+ipCLzjQ0Zx
GN5JqZLXP8LwW06LSD3kI9Ee11n9TM9ecd9Z58rq19rTdMgwUKtgqGS7bUec4aaYuBew6FxzqiA6
OfzWv2z/kQQuo79WotrKf5R9vX2SrcwavlssezVQGz5ekedG5Qb8odHq2xhQhyLyRAZgpek5gZ5B
VIdP7cjVxs1xM5Guv5qgiUhNAsyCmkUEJpCqTRtWnmHZWJY8iPCZucDDyZmQMPfHzSxXnr0iN+CX
/sZODLMpP6EHgjyITukhCR0lJAlT6Jhi1TbnUlGHKK5fyenNmt3CJmKovN0vI4RGkwwgeOHH03ah
6ih7uAQz5SLyY4bppoJHkQiP/oPCIdn5P0ZeSAO/A2QLc5efuVVnfq6P4VHSK3TKqY3lechI8mVM
ny89cpHXb13YggSHG7UYG+iF9oESJZij02fKa3rEK455rlTUtIB7dBdj2VRNIpzZNogAcrKnZPzT
yhIWO0IgHFKellUGibkDgXe4d/QQJvY8EyzeUyRXYaUJjowzHfSpNwT/R7cgQZmGJdC9dpVb3Bvx
WrtMsWeZnIZ7zof6ODRzNOTB0sTg3MLm/4badWb7yCFzw+5ep9aF8BmKBS1X2j/AoUSQKoMpJmu+
qnbvg3MPiEp7HLHfGsPngSv9t5Vr9ZGuoL21d9LPCwFAiN7F5W9rEnb+DjqGJT0hxdA6UGwujJ7g
iBTOvPjskFj0V+iLGmzCSRBf3ebs6+TMf1nZkWK4pNgGQMMkIH59+CSWSfFX0Aht6sw8+H00Lj88
KKHlBKXLBacbAEOhJDfZGfUCqGxEru3vXzjR0ei07B6hv60XAOubLiiYawD2HkGNaZ49ORF6QSY2
exDXjr0pdKufn/gxdTspfzCvqCUBPUnXtTwDa0Qva9i6TfMsDmXBM1bmE/6lUFA8s8K0qi/MFB71
Op2vznRzRIXMpn91kb5y/KRFUO/e42vHhCcrv7GXQO4TqKaZW8ZIP+CA5ehCyll1HY2Gtl8zDu+Q
h7QVYAlbOCTRDfkfPqCfPXlepS2aA3Pw6OmHBg94HgasHGRMBb1sUruqlKkeuE0o96eT3exQ++bX
CJFAkqXMLowWizN4VRtUodXMq/Dz6zIIoC70V40OZPz+SooDUXHgArEB5YyMucZw2/Yx3zfTnpPa
gD6ZSIo01RSwjOoJOS6B2TP3NWZpAFtQMG6/FhYbiA/Bm4cDSzcDiezqmYuz9AVDMOZiAK6QwmtE
LUcoVR6nnFipKRToIScIPpNBgDaEAv62Bne+TYq6Mm+tKnVCNgeUD93Xy4HzhlyylzP3JAYDwgSu
omaWXqKGHgtdUVvCme78Owgc4IjAHM6Q4lXzWKgzHmaeRsdS1bsJAFMENtk/1pW0wh98JLeeo62x
o+pxcckmgxu44Sk3ID46ZWE9qKGTYVaet/SDpPKjrfswqyWoYav32frlRUh6YpvtkNtqYWnj9cQV
BhlvWIjD8aMNcXCVU6f9InX+7uzyUq0AC4JjgBxj80teMskHFgJzDmIfYtyLVkO01yAH7C/7eI8j
duedjBheIFiFdM4ciM2NntE5os0hImBXI35EAERPVCai6YgIxnWZggJZm9JrBM58hqRkCgwziWhH
Hx28kNbBCwj4s3Zkz+V5ts8yd+ROFo64JAE9VLXnYI6OCcYt6YpcRQOzEu3841T6VydpPt8gdQRZ
hhHmtRgZ5OCT6+ZKSophldniKvswBttkbsyty23PaGsIU5UcTwYQI4BpPfcgRClQyWjYt86vijtZ
boKh+Hsm/Z6xF8QLgKNidDbAJ0ygYZC+VBS/hjh/JxMytcP203VMBJHFPtYfTT/cD3kaR5YmzI54
lIsC8+lcFKn1HsHoRBUr9Rbzjwg8FSBgbt2AMvqw0R8xT5KLfm9SlGoCRXo38F0EAZeyHX85BSzA
XEJuVl5zDw9czP+4g/trd5hUfkYyh0e47aMr0JTIr+6S4C6GyUjdCRAFzkZLyJPBEDKG3DVUt+lk
3bKznOIqDiVoWDdDiVTVsnYjTO7vwxl8KvKVUizCjcpdWeV7X+bUWfFyGYKm8t2rmPsDHaARVzIR
3J0jJOSxbGp8OKlaxkwlDB9U+DdAPTY5IETb7loP2JlZhr5aiN5pAxyrRNhHOM482EkEVpNCvoja
I91ZvrmNRRDVCN/IxO0WxPYxNc+onGj+43LAFJvxHartnznJws3+p/h8DQ/Wi0FO604jSG6wjiAC
m5jumNPJsIoqRQQSCesEJGwFpjvWS4Qyd6T/z2U8jKIaxwLgLTE5+WtBLmu7UEy1JuWb+BHYOm8G
C64jjj1nO+dZxzYEYfp0gQwM2h64lYRXapS4miUxz5oXqONjGpcw3DOITsq33BC+muCnzrus7p2U
mSeICM26g2kJ/Sns+rMNvdX9hS0b//OR/LNjn9NYf7N644Lf+s222L3JY1zCZZvSOXEa0gsYUnCn
hKzmjJlkeHwvCy6Vhj2ikyG9sBoVspQJeTtiI1vVYPLW+hAG04vX7SgFppPU/xeNkUOqfbokGl0+
3NqY7W1dtf1bMvUNgWni1wra5Rrbu7dFflxG8NHxQzNlSVkbDUBS3LUyNTVRsCi6KTQOo+w8I3f0
Q5HUax+3iP9tWbkECQkS/eZTn5ebnJ139LfGH5RTDEJdpPNBxJGLmtdI37p98rofouyLCjols9aT
4eX0cG6j7UA90r11rWcXvAQa1rMrVBuMzI1gq/gIWBl6CWewXMFjtYRnmUO73vCqPAcYE3bEU3oJ
NwWYzqUApULvTKvAz451A6HwBDvHqSu436I4AFqhXIDm5kofBuAx9s5o7ekj5nTO7xdGR1yVTNdx
bg709WymZuDD9MHFrppVyifa7hjOzKvOxRk1ZopATGxImCAnZYW4eyEne0cI/rxbdVTzbuOTJ/oz
f4OpfZEirI7O/42tH4vkGCb5vaCWKvzS1UcU+hcKLbdVGf0Cx1onGbtYV2tObY7KSH5pJNn07TxB
iVIy0fWQGRmrHnrEFWHOw5zX7MfL0IJIBpKQ34m/wVIQquGpuN4Al0UNg/z7Ap3nUW7LV/2c6r5K
ImBguXX0tuOxO3nDMYXr4kLJ2uV5QyQ/ODXG691L6HY6dQ5O3wgjPnG9373KbWc0S1uEvSniV3DU
WtLjp2ajfG8NnGDYMMZ2i+Sw6LDaCvSNa+LANhSlZ58nT6vdqqiCN65DgjW6edzrvrZ0KF7CcjHb
yvKhXQmSw+syZY3WykizNonkeoAgZJDdoPAs1dQ+HMITTm0JQ82Aot/TecnEMXEzPVyy26A1TEdF
iWgzvBEJoOApW3wQgc5CcbPz3pSgcN+JXrYgSwgbiNKsOUYfy2WP/V90nK8QEUQ8tjjEHFyH2N15
jwX0z6AY3/3uHCCjVYD/ZtFiUjUA5Hba2BJwOEc41Oe2Em1RF3K4Idy8QA6L2I9T1TFdy6z4j+W9
MperS/JRfDT6WbHntLaDpFBFxxF+6+NrakHgOV/nwuG5SaJzmEpzhSJ7GnVslm8r4YZGlDMAg3g+
QHtKAF9ohGHjJi1C+R/ECcezz8luKgBwmNqIWVvjp27HGIQWG6epI24YTGBkJOS5Fnn6ZKFZb6lg
coEtAABLulBnoFSTL9OF9vo4ixgN/TMUiFBpRbCSbNLTn1YQ2KgcKMTnQr8UcOkrwhyTxLjo8GeN
+xkAA2CGd2KHcFuAqiXj6/zxqLU5rJZeGve8lSXMeJH6p0xufNEl7pty2i3N7TY8S8/y7rM1EmmM
2UyLlMLsQLgumpuFkc2Lb+Lj/nRiwXFrDGg/jKhLjdxXQVU6SPnZomHpbABBEfH2RR1D/J5l2Ofd
GM1jizsRcIiqI3zPyajzxp3MpMNoXAdWl9x+d5gfgP40mjNssuEmhCpc2ivACr30BJQB/R2M8Q1Y
3CP3qpBCRkES7SLgfLhnNOrewJr9fheHtX+d1Eid44XLEcSGibV2we+DESUGcDp3BH7rJTXZauaR
GhkeFyosmV6Z+13YofL+utedFA0JGTSDigRXU8LpufNaoo8p5+mIwWv5cS3cjZFICzEIn7ZzUdUC
QqDGcbekRYlr6zlyb9j6zXWTZ2MKLY0y0Y5yCIMAQQneNwXRRcLF/GOMxDu8Los3QoHvcwlipDwN
T9syOyd2VpaDtbSUT+SZIuq4tL4NyRE4AeEyY6FPSiB/XhZuLGUVJ21NbPt8ub1Sf7QAWUJHlruZ
KP0XJDBLE1HBq2hf/ytpRSSCP3tjDipQFyjc1X7et2l07KuyFG9Th/kVh92/8v+eD+64fcDj7z0S
eJkyJjZS8dTfFUvoAohkl9GqofZhNos9uVs0LPS71JsUI9uEXv0VECp1YT2lp6+EMsnMXy9vQWhU
/tZYxnUZpVoOVbCZt+cvFv53w7r0dhJ9/kIk3PehSK2OBbFZhde2bWlfVa9ndAyFU98OxGTH+tKQ
ZWxd8baQt7wJWBfCtwfLA6y7wczuw5L5afeCc4u1UN/V5A9ZZcZLpFka8ed163GJrHDOZFoIdANj
f3P5xO6e8ZHRTt0Ljem5VF/vnatKZZtqQ8D8xfxIAJnAk++NMTpMCPpgK8L4K7qT+lWpoZPlh92x
JroXkr4MSFZuj5z42jUGw7OH3wpR5b6OS1rXuFthokP2daY83bZ1eo2uW3p7dHm5KWc8r1gLylEW
sogdwq8o78ax9qe8OVOKbldkwdFuaOJ+kkM+H5gD88Qm0B93mSMnE47Ur1Pnj68R7G8lvpEu20FM
pAPeafcFKY+y9Hjdm53C1r5coHGekZiJbluOr9cE/uyTwGUYcIKViVh1pKEclSI4dHEHjhEZJ9P4
x8Jxnod6jVs83CvuABIuCYoZzXFfxUy4SsYerzT3QzsNjB2rnN2L4MwOVswFt3vzR6doXUZJdR69
LK4rLbSjYG6c+lSwwVybWlhbaJKcd+WiAXYWSUBF3DuI1F1yCPCevwCRVGp4gd5+6ncbh6cCMMlV
BKCkOLLpCVUBX7yUQWmGmm2thTRVQX0WQOA/3NFB9R5wrfrS67zjMN9emTilJSEmTqsENL3okSIY
mVCCwZgHzQaxsRdmjnwzwJu/cPAJusvm/EQeJG9sW4IqLis3LeGglwyyh1rfFBISCtIkGVXgCwD6
v1O2V8rb8V2gc+2u8u71ufkVmp/NISNKl4qPNvMiwoWJgt9mt/net4WHK5pN1s70Nz2RBjRghvhC
5mCTnSkdn4kZmhnDrRBtHQdfp7SQ4kUnR8icpinA1Fjrr1nesZkoTF9Fa5frN9ipTUSI9YbdPMn2
TS2BASHiFWAaaqmPBP6Ki/r4krBJr8KEw8z5gqd20+QZoYG71mBIePcGjMW7dzKKzqNthQmh4Er5
gekRGJMcsOan5zYV7VK3HUZiQseErLQ+sv1mmBcU24eCnKvPNAZOt3EQmvGVHsDtRwO+eBOyyBzn
MoJH1Glkl5FvDSVYgEha5oQoq4H0rfRHLtPVoxwS0Uixw5Gkpd7y/KaE8cBmpzqXyUkEDLlIlDKe
2OaykQCAWgq5VodapOh79MvvLaKsVK8fHEwv4F2l+9WE8EP8ahzgrXQ/TXqHMeLtlYhxyHXfZsQc
vb4E+aZUiQvsOaUcP912ksUzbEyCK4q4IFGxEfQG82k1/i+OKnkobQw+gyKVaNBbzG7mfEdWM/YS
WN+iS9QQNG/lKsXfIqDSdUW64qWwEm8WK8wG8o0YIiMvNjX57gQU3gMxJlwEI/le6WYeWUt6oKqU
f3xy0qxozySfLM1dsrXfF336/2litWdS5H60e2sLjXcKYY9k70QcIKeZGdWywemgORz2KO7DzoTv
ISDZZdBPp4EzlUcZrGf7xLtYVa2Hb8jhi63oG/De0+4VzXP/Bmv50qmT9Q3/bPdynLGQsaoGK/YJ
/8N6mIfxCsx+BdexaBjU+fonlfTY3tn4f5kjlgvSVaoiKtqKNTI7T2Y4A9VG0OeZeNSIT0mcg3xJ
7yuBX2PSHWMGKI6A12ssg8sK8s5RJ8xKWQQChl3jYKDu3PN1TGnAb/KlPvGIYwcXUnJ9LIYvjK/n
WZNC4LHfyO+sJuVlCpyTRs4vIemVsai6i+ONVtEpnjyBEl9xaDhorkQj3YiqipmvTA3J/RM7yajr
7FRli+o3Uk6r8G4vyci3rUq0wb4W4mxTshH9Cu937UwweH8vHZeP45laAjrIFXtqRiPfc0EkoFnk
na27oBj13OAD2T76S6nlxOg+sf7qh88u6TE5pqVFBCqBOd5+bLybLNNEwaK7LoaKj7gcPom7CZpz
1D6ySSKqkMtXoWS71I3Mgiz7kfak7Ph5QfxSP0UiXUlkqfHjfGXlgs2a0aiPIuYkOg2I80QCn5oM
xEudaoclRUfWiSjnTpPEzWco2CR6vW+NgTB/3rCpYQSEll9bGOkK1LZ3qh8mU7Dbz48Kiz6CAlY9
GYtg2GINWFVKaKpzrHrOAuw/ru1pxA1M6WV1iWlBNPvkbm4jSLV17DlNtGNcr6YscwFLOuLK7xsF
CN4YGhqZSKEg3F0Iq1ejJqHgvCCBkQdrr7WN5PuAmxOAVIQr8dw++91uObYa3YdOVCNnUMViWtZY
cDT5eeOiAvjap+VxzbbP8w/b46BBJu9x1srLMYh8hQlqMZB4hTzdkgkxZVlQxvuxdnd1mAA0W4Up
5mgnK7fM/7TxYTX8e5gei2Py4v8SCGO7oE6NtQ7Dl1j6CUBZO0L0sB95z0AgNZvbFX2UUoOxL1tG
GYudE31ricKTXMMEP3BxmkPyPWXl42dcwoMn40o+uFi4vPRk9m3dinW3DAGmjtof/IQmimU+VGM4
lJ5+c3B4SR8WRKXQetUZ5M28ja6XMz6XhknOlJbRmzpLe6Evkq6OJYQbYO7vcqRrOyTOBmeZANkv
4xnJQ5ziCnt2TFF0LOPD8D34fSo5VkEiHsnu7+Nz/8FhO8FnSJrZq0RRDx4078tb4vllioeq4hcz
gYeUmuWTUx1IECuhrYfgltxb5qM40weLzA+LMVM/IRbif2fOBNIIPjTo//64RS8SG0l7Q+P5//Tq
kg5GgIpQA7QfZgu6cn4bzETb+98ZCSHs4OITuSrHdXGOxDL2OBlmZsEKauvtR0GcbqmtPXYQbzoN
ltJRCef5PNppN4nppCmLKWJ9PQBj0ZLUcOgBZ3wg6cqMrO4PvfgEjQ766alUtW2/ArfeiRpnVww5
amXaFtEJUC3KXfWWNgyn76n3KxNMnmsQG/Uauxx329AQX8xfNnWT/gSQKigJbHD2aqCJ3YcbzJ8/
aJDt4exHNSYu4HLybEf+LcYlt5ompXUgfSVYOrOPsF/C6F08iN8xgwU3l5EfvCXrcAPcemRRV0fE
nTAgz7tCVA8nr9QtPwMNKe+hvt2kRl3a7lOC5/tnhlIRgiH4FY5fRrwTvbITdH862bVyCyyUD44X
KDOaA4Qz8v7gecp56JHC04xYcE2XZynQ4LYUXQqTCDhrUtgMc7N8Nf/t83LlU6CGmbrm3kxgXWCC
p3GfOUqa6klaRSmjkw6TOTYIlbBlnQ+QmED0km9oOgfPcEerGhxb0C2YLxP63m72kv2XQ5+Xe4Bh
p1c2j6DoyzhPIooycIxnExYnrxjJD1GnWNLyzYn3zLx1Vocu3W3DkUcOFUB0VA9rBjud8LKdp9ym
+IbSrwkaLz6WWwWwAi84rrQgjM8FlzPl2G4zUhrsGypQZN3it6CHm63Mhzs5TgwC1KHg0IXXKx3Z
u0JzNWvHPY9X5p5kVPGDcV0KgpMOq6k6u/4Tmj3UZKN3QsRM8qrrVA/EieGh0uPGBgx5q4dJrPyy
vVs/aFI4adrtLOSq7St/XdqqLFFnNKwDpnjmewtfgVOzjE42CwGZCj3W+cZq7lwA4TRSusMcy1eg
NRkI9Ek6mub8Y+NgdZNJm8JvZOkDOYDwlb5tBAA5DNAEBDznjECpx6mRAnJiE+luNtSdIMsfrp7M
C+K9L+B3t7R6ZyQ06wxe0Zi7eOGMLaCcyBcOlc6gC9LggKUM3mw4JwiaGoTlW4HRUOCgiV9G4J66
mGsOrgH03Hg3L9GUfMeNJe5BRMEuDCRaVvd1OSJ3uzR4uZ9JS85MaHMByMd7s35k3Tmz+Tg3QCMz
4KiCetqZ3oMVfi3RPIgVaPgja+RRJBrUoytmLv/ovzUCozPWwJOTuDWuSgGQQaIWY28O/2NTWHBE
4p/o2Tj4BEj9GIeyx2G8nZUGCPIc80r2vBKskP+wqj50E8yM4n4gyavyVlRYDGo8to8WCm6aC6Rr
FSASubyMunvsmC+cYfX1m0ko4L8hGp/pXwO/XFbl0lxIFx3KxRGCzwqsTHQ22RRzEIjV6YnmfnQx
j3DEtNDru6KQop1/Wi6SBw61oSJ4pDd0MFqeUt2VCFpk1l6Tk96jM9qcA9qaIm9jD35Aqq/kLRlI
hMTBmevVXJG7PpVJ/Nk7n+tDhRME/EgPfL8ne+4o/PF8YWx+pi/qvIA8B5SMxgjzb49li2SuI6jY
+XvJVNB93gJ0YuGduGeimyWyhjTK+Ua5hCg+lwcOHybShW4qe0W749gzlPf+eUkAMq2d1hox2pfH
jjQlDhtmmuEvPGLAOWNhHEyP3uZNNp1EdJfYACGflbz61LrTglW+O52dhtZrM7oU696WJXTKkLwU
B2WSdfI2fhfFSLO3c4XQPzHz9FqQglHQzSZwXWQ0R385u+JxJ6DdjRzgoBs6T5eHA7ULWuREdh97
rp6AURu43L+u+tbCYEv+uTrOK2BZ1iySc10jWw+2CkWu2hlJF4SkIOkVmkmPY21201ZSytwWEb/O
5xZOjpmVYeciuj3vFGd+Z0glfHb23Zv4uVsrOHF1uhYFBTQQXKErS4ComqoLs0+83e11x8lFAfxM
VcSb5fumTzalt3QCqJPns/oercTlnaCo10l+bh1cb9OWqC1aWMLPx6hAC8KI3PkqX/53GDoRtgo7
UId4ESKc0CEzm7O2lZguhxe5SGVRVKV/Eyc1GKqCqBhUT3jhYe1XTBklc+tBsDXOX1qFk5xIsbhQ
eRdVT7Pg/lMpXBP4GRMMNX4zr1qcSel1FjrA/XwbDvHmkP4vpa5H8VSfyrLxlgPtT3YNRuYoKeAk
D4wjN53DgTh+x9KMjGUZ+90EPL0VDZkJyhLcDlT/CBEK5SaeWqpsf5T4NPuW3MG+mjkpprn3omwR
ADrEiicvlqg6K4Gxsyr2ZILxUbyXPOzCVBVjuI7i+4OiTC4a1hfB/RY3gSbc1UQY9hD7xX5dAUOE
qnJsJvfybu7r2aXRm81psD4SpN1KSTi2yKIZRsdd9iMKvkaxfSoFYwJ/DKAdsYO58a7orJ3KOFcn
Ic5RWnqrKtkYFvU474OdR8WDWykQM0CtUTUOvKN8WrbFsUWhx2qPQ8dI7ZCQ2ERxo/HFw3c//JXw
28RYbOuaZ8PObE7ZSdfHpQ/AUhNvb8pygQvYJOKxjIDDpvP0PiBNzwc29AyQscoYJ1WXUPd8khM2
E6+jTw+PhqhBX+SdDRG9flhp9nVCNjspqxv/fek06EHKkHuq6ss7NWs8sui7WuM1djw5tEfP+Le/
/gh/v3fEHEpv52AlFGJhG2LLVeGYdd0APGsZYbgjBIq1ehuWkRz4yCrL/s5spCYre8xtCIeCECiA
TDyRIUGh7SIwj9kEGdON+qcRKBgcHW+yBHplZ88dggJrPUByiWQCZkDKTmdY2UVfxx0ArPrhMzxi
BcqE//jP1xbVV8YXBJ87+PI2wYiD9BuwPKe+gkzm4vgZPcnAz/X7YK20ADGmsH4HKjNI9FZPu63o
C6a+HWYuUbVq3d4WcAhVo/pFPwIq4Rok1zqLnONzdthOhvGCy73Y3uI1J0sYvW7jXhUK7zItxCEz
4j3AN/xf5zQ81jloNlY561gODvqCxNQ9HJfSDZqer70QiKob0uDljSWKaXwc+/VQHSJ571ctXIVH
WSCNFnUcHd510J/Trk+fBlqH4GQ+lPFvYoPWDBmQVxFJf34TlB3QAAnsLdGrRaoTFX4Xp4ygEn/F
9NJZbCSXfRWS+XotB2W1LQy8gEOSpdnCd/uz8N4rX/ecco16i91D7amRets1Z57DDObg9S6dJU7p
P/2YdiG1ErfhLAIYsX1qI8IAdxgDo299Gtk4CEj+lBh5RZAgKppB2pQFFHn1HXZ+Ts10+BiPL3OS
t3VT3jIePF2fO3lJyf6EPO1vI9il/oLqHwGiDzTYYqpF80qjlDjRaBBf0l1/RpKsCGa9PdXqmFhA
+SbsT2WHcciuH5xvCb5Csm8rB6fBA97eV5se/Ob4zGo49xha+DGwdrSD3raz2OWFTkzNi35Fq3oo
ewwhSQbZKz7oRqxMHb0OgnKqQicCTnT6ecJXU0OTWZkuE3dMDFfYWj8MzxBH6zwopkms00kAc2l5
BLoQme1mgHflOWX3Kgwh9U1inSRnJsKXyk9BuwHSRGVroiw1raWxxakhNX2iZq+IdFMIkRJl7kkW
QUTtlqmQsRWrklQ9w5F4g5j2WzOwVzIXq51UCSjuTP+hknKliW6OVXNRjpQvrNxHei12OnD+zO1k
CR9dAukFUiq8VoyNz9Y9hPJOFeXZsG0216I+01F68ZLolsNiwGugk2+PNAHsGmcSpugubKL0i7BT
HNK/k+qVTIAzuhK7F0LToXmRhqtCPQG8dRjBb5ASwZmfwJtm237PcpVk5VySD5y9SvU7zrduji3/
cODk4/pUPD4PtO8GO6xw2Y6BoXHtUamml2wU/XwBn2l8CkcgLL9xpoplybxa31nns3sY08v5jJIj
8ATBpcgfScc+Kgqf8Lou3A76DDJhslqUftMuvskuCBmOSgsGU8ft3AEQACUEpVtgT+JrbY5PixHA
APxORI8xJiYZI8UkUTxpvgcbG7JSqtJh4IRbpK9WaWmCMZ9fGHWeOrlQwaBgkpVsQoqZJxLLzFG/
PR/D/IZyPC4xcjWXxNVrGLqTdgNgWowYKNKaKu/GRtIo/yQW8cWlu3CAuUnTqMnnhJ720x3nZXTQ
xX8PZ/6L84PEwoVBwA7YMbxDMYCOYoSXP34SDLX/lKFDwdA7d0aBV/t+qedpaKqxCTzXpWet0fpf
a24hsV2m4vDRAuOd7eqR/2UZ2WQ2LCwPBa8kKCAnzFTi/TXpAzyY9rwgc/E1etHxwik8lwE98hEu
MF3tAwaoVoAq+Mef8BOIqrjLOGxS8mjfkUsnNy/Ujh4soR4lST4iyCdcZjZf7w2fzdKW6VGqXSY2
oB6yY6N7gciFmqDJnVTkVdiqG3/njhUkf73vDUWzUY4fpgNANr/pxz/9G3kR5RkDbujbD4XsivVx
OSeR9UhUKZiXjJzh6nAEhKa+dai61iLAap6n6cG2lK85K/Mee+HBUjx+nYMWfBhGkDK3KWXdAxaH
SoRpmNJd4osvz0Zjr+kRE+WILbs/ZSg9NzzrNrt6n8ndDu3cFTgakUEFclBDjVtgcHj7qInV2Wmy
kuInJ/tl6Qjy4pVRR3aUJiTYSqB/AS8ehIzMNjIOcXmPvj2uL/OuLox5hukVLU+1tA3rrTU6gKJ5
VomwedrbNoPX1j85qBguh8duNQjgf+HrL4CIk1zCotonXoi6r1ub99m0el/FpQouC9MRQiqnb/DA
y+QpsDHNQJAc7n/wtJOCjXcgU2CB9nuuxj/JzFOXIicqLVL1eQANtq6CN7uVNRnrfrwgxEC9hv3G
DdyEfqor9lkYoZCo/bvIjJrRgXPw+uW0jpRnujbdOBXHX7X6gP5Ll1PDehDVJU5/3AUuCkTb5E2x
3mInyliHIZEnSBuGKTIATyIWxpDS6fvq07zXjylcZmJGtAIW6+bf/JCqWGUFEYZn5xggSFURD+Oh
MnwF+g/Ww6Kkdsw+pm0g15nQsN7FlQsWy72btHoFknjkKnoK41+t8VO3hCVcR/T5FNNaApvweTmm
TKyaj5gjmTsHEsN4HQJHMI95cIMlUO+fLV0X0wjJNoUJazfsTh90jOaRBqCJBNex1vwSFnLEV8Em
rnAafNAPIhymxlQ1Xhp4eJuqN7CKdEOUMyHqPVDQZrPwOsU1/b1lWGRkKCdtyhZhSyUC84GsHd+G
1YI+dFAlrrVLytZV4mAaUzGmnhItdwUrtZt3nB95xFWe8IBoa8S4ZS2+2W6fYChzbKmg1+XkN0dd
Jlt2NjylNneA2NBsO60+DXOmHIftES0OiLiqKuubrbR3U4BfN4GEBf9EsRPE6PO6AI56REFvMBPs
r0vKWKcXCZxxKOSF7aBJZWAI1yVKjmlT/W/ZU1OuOYX/mKBEXfZ2/uHitMzC0TdXLK3k203WUN4p
zTzoGNbay08e5yp1HbNkLkQW1TIzXc2ewsYo0T22h5xpotZsR0ZpjC5X8BZ3/fYsu9/K64OeKONy
k07L9yaZ4pcBiqVQD5shZk905mX9Vg8QJP0Y5P0oGKgloqWsLecrMz+X4dGU2qVA4N6GDwj2L9pJ
NQH3aCzoz31TIRFqIUVzE9StBqkyiS0KsVaj23x7SIopnTFWsNq1Tgns7ewf84c9O5oZR1zUdpV9
YXNrFe5sOhTR/VbaOohqUfKL3HIU0Cl49QzT2R3pdll2a9ML9qH46kezmZRHffD7FkIQ8JZe+6sC
e8Fnqbq76JsWpNXPhCEhf0mj6Z9y2+aLhQv1hENF3uTxxZJLiS9oyWm3jOIibkv+GwRQEfFjnm0y
k+9e1A4cfLDqonLUIphcYLND0LRQiDPPMkMejMTsl27kmexemjBykU3daxa9S5UWIDk0+Kwwd/q9
Q/8+t6IE9EXhCQmXVRviv8Qie68GKDKy2VQemqhlDD9aIQiBAPzlx1sFZm6ijzlgma4OKV5Z0gPx
4sfqsLr+PdK5n84dBdv31S6HdiQBIMxqDAwUc7/L0VL2RuVie8V2JzXaQCfQGoAEKRDfed6N/i5P
M1peNYhOYLBiO4LI1Tu7i3TqwtNeC1ZuYtqXWCigtlrS9T/pay5C8HA+RD2kirjjgki6gLmkEZUm
ueOxC3oYlF7NcwEnSNbNsqmpiR+R1na2yClTAQnX4vRYJyEx1HhgY5d6L9olhTVU0wz/nRbYNTbc
Ac3hOI/9ZAiF11UMnTQ+cvaI4HOKV7p7KBUtMwqqMLhaxVVmAGhRJsixlRTn/5lTZmf4orr7Gt6s
fdfMBJ7W5RbPiwV+1xIE2/NRJmAVb7nqAsjQb1cOR9ZiNGmr+E0gNQLK0b+FW2iWtDu1akmc4TOW
UHet5PqRw8f//GNbTRH9pGjhHjIsrhFYU3tQw82gf2SP9rrEuWexO24V43YpYFtraLH55Lf0Xvbb
yNOsxqSPhMEqgD74CI5Ha6F0E00AdHMxeccGvtRZ9gMACStO5Mt0ouLyVCIgRPjnjHC++SBHZie8
+mXdrLzzrIw7XRfxWfqIJi4fG35uY+0/7zfIhs6eYKi1w293pA7EqAHj3v2g0oJHFyhnAKzOko1x
WbB8VMbRyc/kckJ8zMmzMH70bvYKz5s/iW9spK8flHwIH39JZpODQML87LMji7uHtySzQNVdNtkv
XrwjkkBUjmrcVVEvj0IHtsQaEzdxQcjhpEutgDjGs2NabOqs4Fmr+c2r0nq9seaiDVqU69507F7Y
gv/DXHmvDeKAtbA571qIh144tFQBRQsYybiZltcIonpFMXw/SdFE4LJrh6iGhsIpnryqHILeLHiW
TURl2VZ8JbIvqM3nXJ/702MR2S3OkmVterbxF/oF/lQ8LL4SvVzN7DaU2a+YHIpsX+8xAlUoLMta
rL+qCXO1S5B/7+1VLrQTefeqwpPKVMs6LqUR/dwmaV+9zLinpspy3MOqai9B1pxtrbUPsoczAWjW
hJ0kEAy9aZZnf1G3FoMq99pIIH8mzh0OrFQggvYS6O+d83bBpW6ZFwNBt1bPMbzmfs2AR82LiLn5
4xGrGcIx+COEUCPuGSVO+qJmQdoWdqagGa0I7KAfELErYn9wTB9gMitiO0RI5OZcEuYSL3MrrMOl
XwYP/AvjLgMnKbpf+TIva6InfU2mZ2Ygds+R4Jt/OW1ShSA/NlQQnXpWsxfb1duFN11UCNCAjMuo
K82yfHw6ChmFNKRZElGF1AT6sCe0qusQ8EQfQUrgLJWqKDRnHYkuE7CgJgsdW3e8wosXUb25Oury
EbHOIZhYIM/lJ1FhTLlRtdTt2UfNW4S1xJ7l08+68p83CPXCuS6h+a7benxu7DP6U5D00trOBwf6
Zc54WiF/Yvzk9zF0BYdB2nZ/SS1sadJjMkqISMDVxZFhBWmzGplIkv6EI5JAfmDPOMps/VxZ9xLP
EgoWiflQRowHShhBS1Udy3YbVtfCkD37UAF0n9aq5qdbgJ7F7KsCFbq8h0Z/gkDZDoR3xA+kaqze
O2m75S90Xom9TuRuCc5j3nJx4KZvwJKv1BF0Ah2Kmq6UlPOsAJJpb63mKY2lVMJOFCmCsr+0871f
TStOn7PhW4wtNB18FnuYooTFitX/RdzfEdy1gwCuOqlvHgACZHH7jkRSU7GGuTgogbR1O5hGz6Ax
lbJBXocwcNhPbnD925N4f2adFOmq3Ky3I9dLQJjiogQdw0ZvvNS5S2SbP6gqg1Wq8RB49ULT8Y23
g4sVOSq0oYyyY4Asl7E3VKY+Yjeg2N3gUWr4L2HS3/BIsyOyzk3SBwqscCjiwjbpEZCWrf1FO/JF
/78cRocqMwiW7iuUuMnUhkbNyBNfxbVMPYMU/+Z9idhXhLzJ6HhPptkdGRsj4W/mFXnb+0X3MRQb
D6ehdyexTKLAHxKBoe/pfXTciU8qlUY8mWXIR8ZhzGspeXT0JcgCjcGp1YaD6PwbGqHo6fRTUEx7
tH8Je9JggW2C4dSkVNJGrUH2AVw+C3rSwkQ8qQ7PCdzBBmk8AB/RQHNSxFKiV10oxHrmmoUNEik+
m7oBy6/f8oRsGeubZ75TCCT9eEyWGcXj+/mT+DBIVBQ2MRbxK6668u+RhtzYRaRl98UsK+QvSuXu
tyvLO1Mm1pSIFcRF2jsq+nrTGyMeZcnW55njQFYd4Ns3bYdIs2c0HF8IV/oGzw/SBLVThLnYfmIG
kQ8PaV3loNDvNqHNue24YCWhi3xUFotUI29LIYjFC6ziJYqRTNbEpR5XVlnFl3eoXBuBntZ+Llr7
QHlyQx843orgRRdSmnPtvdgnzDfejz5bLWjiu0kQVvq7WFi36y5m6wWi3+LAjadhYvwQhTkZ9TtN
b4h9TbZpgYY/jiQBfz6EpOH1x9hk/YJT4cK85bWaXpeNFhXTnmDuZIGqq65Huug6cS9wtpqJjXJ1
PGDT4DN/tKaW/ZyUZCYnGVIAI/i/+1sSxmbVShLIU3RU3GtuW+W5LERp2jm71a6DduQf4VpVwL1v
oO3+3vmh4aV6nfhC6mFj6DBCH0KeZwPDEXkHKf8GCnOv3SixYiI/Bs7IUYouemMTHiBMbLRDxC+p
fCMVUHLKCveK96mCBrPg4EdVLvND7k4N6EQ0/uDwmJkJnvN0IocLPAMtbQ5ixBsFGyskTa0Q3S28
YYvXQFkU1CwtNM2CxzekEkRfwRQVkLUtv9E0CD94usp/9Ql551bQxUXemQWaiT/XELrv1iyNpVNL
FlXkAewytP4F0tvJlbgGAxuqEcnqVFb1CvK5UV3Y+qrlr/5F6i3xLEj6S9j1gW6vZTPrXCXWbxHw
HOJONKIdOC7ArgQsqOFg/izn8SjQ7bikoPbPWxa7hdPtXWMWNA4kG9XK8GYdu4e5rVbogrbdWrF+
FZDL+mFi5s0lSUOtIz2MkQQ1cx8Jbu/NZGDMIRfzPmJY4B5A0YOEwdnaPvsfpx7NJNl17QAX/Np/
iB2vclMjfG28vJ5O1XKlmVyFCfPE2e49lNswPy9nmi8YFIxCLmx83LAmmQHEEDRRngU0D4h19X66
5RyUH8Oe+MyUBOI2iQamPT8PFtmEfJf2EGdH8nq/RUJb3xxkJU5ld2qvpBNvlvNVYtcU/qzXPrMg
m1OmzXcOO8DM1kbepkvp94jlgJPAucEiYf44E3GnFNKfaOZkBYv4ISReyKZHNzoIMlVTCi2yTAaw
7NUw9jm5IFWlxUW3J1f+yPfMdEhuunhpewe2nBzJzJahCzGFx64DVIx3rfmJPQuA5vh6nufO4PPK
5G+BJvZRBScNa2a+ZtfaewF5FePuf/ROZEOjLlsQXSo6OmGiPwxQsC/3Jn9Vz/3UUfKUonF9IMZz
B6cKmPUuBoBxrSG6CpcvCvcG72HavIzfIKOBMMT1Y2huzPiHYhVZKiQi4r856YNKDZaCiAX6jMLm
8moHW0skWf0ukOabo+gQHNMQaznW2Tck0KhkZsyBkriWcZzW9RQMbZ2poTk4sMIaqvNGlLn4VutJ
abXE81r18cuwdhNQ9DQ5blkdBDq/wxNC2y6L/NtNkcUSWPoKeVLtqgF35vkGX+GkYbWkacg3hCvL
eKXnIkgOuxu5F7nIGbLIdkQUDdFO9LO7EEGIpcAhJ/qjtfd+8gcpeAj7Qrv8vDeTkOs5ci/LysgE
joGCsprU510eX6mowmaDBlsV1sTSBZKTppEd2OQPL7aStARBprHisugEWqdEGSCiLZr9KfPeK0yv
tpFDahSejDazNPaAOk67mtob6fXrRcXSTZ0ZRp85ALTbF7qAFDBdbBIKcL72V6kcMobyIinODsyU
bCeAyJQkrgGo9woCcc+zrOniUyJ/nSbRIhtQEfZlxYT3ui0QR+lnImowecSMs2b4kFKh1Tu30q6n
/ppXMdL+/8QO0OmCHQo67rW993nR6VIpMviDe+8PWbSO3u3jQIbNNbn7TLrdPPiuUEhiQWfgMAcF
CC0ZAgNZYPgXzr2YtNLPSmaL0ob5vRriJc4TG17XbYLmN0DsRvHndUbxRWNrYom+DACFz7rhisoL
3OHK99orTG4PPztNM7TbSiD4bKi0e9aElalPZU8VSNCSnJOmS2uj47fIQptYCRMfJPkhn62geRC1
lksAZD2H0AySE1GfNNgJ1JGeWZmyrw8OOkaPnv23OFO49KOXtXvj5U0WDeiWXxFCFW6Qnc/gMmHo
DteW6vh8btFrcyCyStf2cx8aMKJ3pA9Fef7vj6BNLqZkcjslHLARXT83jpRqP91s+K4SzC0YOEok
FTgiYxfh9WLsFR76RGNpMPoR1syW/e3jAkFK1iJEQJZDSyx3Z8jM8ZKlAsfjBxQV43HVnD7yzDYz
n2NJEDA12Rd7dwmcew3/VFLhfac26gHHmdgBKtzBdbTlkmPLrAHzIrUGLovLEEe8MC9OGw6icHXp
q4otLImJOZ2iL1ZM0njVu5QUOJY1yozJFJ8XMkhYN0iD1AFEsp9LwxKMbJUZmGD3YfllgH9kV1Wt
eHm4cwj9zIsubTV3TPSANyyMabfelm7tg4wgl2fOxJumGfyUjsyv3+kZygmRhRt4Yai2cp9WfOJX
RXK4OLMc5KJ91a5kZ6GcGSR+VUIYM7AHFQ33h4brcc/Z0Mjp2gknNV4Jx2M+2gGzlGTnjELVzj69
agQreUoO5nyxZ+ZEPiYJ9Ey55A1y6BUbpcCtDI2SVPK7/+aBng+lP8yvTWPpy1yv7cdrm1Vr/KQ6
rSMFA5BiEQxGXKAUNcxO4bvRGmoi5zdo7hjhljw+OWqTD78f5txGwn5mIOPwfJTLF+TH5N6dGzqu
nBHcrIAGh9Ua7LI4npRKL9p3BHm513kMi9TXvxcSZ5UBrEQPsMPKdYGqaXPz8koWQtrgg4I1r6je
EdZ7BarOMXqoRXsfauqcaungUF9rDAnQsANHepMPPzQFLRb3a4oHuTolDf6a1Ql6Zz3EQwjGernN
F5gatnXC9i/vZa6ftpNmutoTG6yrD5cnGEHEBF7GOcriD3nRGN8THmrV1wR9u534DUAJByN69sjO
KIyTD9Vn0VN8RP4o8VwhHsITCqYbmTJ6ND/OWoENdAxSAI65vONYg8ucQo68cPdAr05PufyR/Bq/
YCm0LZxeZRXR0rJ10nz5lCJZxMZRk/fOFz2UVi48Iyv99YWO3dcTzwh9TLtJwYzyKu5fqhpOXIlD
f0llhxm0/k831Mh8UmpWGqapICnvIlXsFat/MNufsNuCbRmlEYPtz6nHOSMXvsNPT1TtGHwFeVLl
pvRl+/jj2B9fPDnwfKtrA6/1U4sD95OI8gULnIYEsgky7I7q65kFA3F+ujkGats9YDyZt4lXLTjj
0V0NlUcND8HUxoFGiyiILWyhnZFQsLzek9EVqLMPub0AM0LSqAMr+upUU6+IHQvwzub7HL3HbMTX
jnRBqgvEuCfeiLeqtrQIfm7JPTvEMrjMv0Ts/lcxblx53+kWzyaiIUc7/OTy9LGRysgxq+ZS4IW2
H2HacJJVjj4u63mjDCMJGfF0O/3sLzYo6+cc/WfQAuDWDR2ak4Pawf3c5IEN54yT4+uyRKY8VDZw
ALEhjKwwTQ3xdyIVfdgjfA2R3gCq0c19lsIkxZrkEHm3XHFllHn3Rjw2P9dl0/ccP2qBViqXQvsg
frB+r1I9E872gAM8d+em0PIGkkgtnQ7gUa+/2GuacjbSV60SWQwcGuY3OXZdLmOVLuBKHa0PLjCH
etJwz4QaDcVkSu5KPQX01o0ulAJwO4L+oP1qB1vM/BJ9MkO226l849aPRSNkkSKDYwPqwd8BexJp
SoUUA9mqUWpeMLLEkkoR10mL1mQrIYzCivhVOkhbFmkO16ltATwYSPL08NGuUqfssolVqF5AXv51
o/VQDG/1bRUl/rVyTB4RUU3DZop7qDfNqrl0GFz24yZsoOodcjIISggsmuq40X+Xv7b8KfhSF4bN
jZX+fo+X66oT74vA3/SI/5Nrt3n+0moe5Z0tmNSy8x4BdIs+Eeyas60IxuizZZCfvJG7WQTzrzh4
XhJWq5LNymtuOsEkyK/t9gHG5nHgBVrpw3ryTUEH7B4yUNY9FecugovyRSa32GxQJFk1LKphTJag
wZGAvkDVNMDaMHqsqsEsgHDCll009Q3DxBeOhcTFz5vijZuxToy7IgEq+8ZGsCtRdvZLk6+1wTc6
H9/TEryl2yxTy80uQrzBwprlAIuZhYNABePjNAg6TwI29FLpYVTqPhwsH6HwaH4321Jk4vCrcRu5
7VDBk9T1wxiwukMCd8JyRNTJ9vWicJqftqQEHSA3INdvG+ylteWxs0F9wNPFhlIwmH1mqv0lg8pj
N+imxyCtG9Zl9xrHEUCcHGaomdVXa3uh6858j573kyUdoL4cIhUdKtsLDyg2suhIfNxUkA2VTQ3y
fOafvy5RWeYEj5nHmfJxh6NftS/xvP0L1HzY+C+pjgLmdbgDMO7IDj2hN2XsUg05H5itqwhpIa6I
FfHhdfWyYEnd17O61X5s4kPPD3TVzcWoIDbHI/qxaTvaGbAzQAIf//1oSAb0hvh1K1m/rJx8q7dV
pT8drXrv3aY28rKRDDmCha4Ynt444A2b9sGcmeCt+0URs8oHLnZZkl1woc3QBAC0YOAjwDn1vgyF
2LGI+SIUJji9ks/MQ3bQSqK4Woxr3E0FSVfckHMBXobEIrd5PmJ0V8iRxTDKUsvtqteNDAedQinQ
nGyozTU83mFu64TfIZpDPASU6QqQceTBoY892+TwO0/Xrc86VMAXl4N6vTEpcjDp8zjp2qpCtg5+
yIiFtcdkXMyKInQh48Cujmb5/XKUc+UlqSnhDaG7nkbT/kulRAkLIK3Gyg803FU6h5HckFfv1Unw
NRD6o38GsCdrx5JhzEG3wgvTI0JOFku7NtJOZ6CvhvRdESpLuQPG/h1ri9n/oOpYPaBapZ8AFyhe
BoCuC5NcDi7JK1/hu0Ard/CSR2Fwey2yJ0Bz3v9Sxkj0zJKbaZGAYlI6f3dszcWxaR+4S5uwEu5I
w4+K3P0J/B8dGJyyLWwL6hD1HEJASy+r6ddQmOe/Wq/X+sVkz8d7WlcfRMWVJzotw37ZkOcR3xmy
XXfNSGpooDZqVp0fR6oKERbfEXQ7P/w9Ap7D3lHZ4SM1s1hmsz6gDM9IPqfmWHEWna5MNWFZecVi
kGM3tUmO2trFO/nCqx0r67vk/za6QJcbgROItwm7VZQSLVTfqANlhdYihYcF6t8ih28Ljs0j6xe3
kqv3GRNTVe6yBsEx/jQDbfee80AmzVRfb8TKX9jnDazacoBX/TI81VQBk7NkoqN4EfqSly00WIa8
toOAc31xxgrGC22iWdWsNU1TVHO71YiI0lAf5fFaJhDarQJKmJHvbRJhgRm5Wxub5fgiNarruxns
XmQpJ5FTy28wDw9SkMKuNI8iTgmFKBS+vk5HDynxx0sA0o7PmubSMyZ0h7BZDZhAhXDZuySeh2zd
+EHV6nyg4hl9XU9o1ef+zbpptVOfzN0bAJ3+6w+vcgRm5QRiSRx6rI/wVZu79i8MWcnpYmrxfwnS
QGD/BotBFNmVhoF+KHsO5uSj0LttqsepK7Tz3bs5GgeziRfQ3skz56Bh1x8X6+2Eg5HLAEje3J5H
8yGtoGPHHPOlUNNfLaKR0yr0jb+2aOD8tWsdfDwQWzd3niWRXJX650/YgEWhL4KFq108UF6iHybm
SsWmmBGD0JtpVQJQWqHs7fk8o4d1ZH+oeEblKGNc5b8EW5xO2d+gRBtqFT0G8yWLve96I6WVhhHs
1gKzi4HBWFALF6ys1OGTjLax6BC7F9Orz0WjKiGTssNC23rbS8/zSnscuGPChwBxumGv1jXYFj70
BKI3HdrpqZikfwxSZ3yBkPeGaa3fBfTzi8E306CIERpMnU8Oo8IpqSVyqF5gfnt7pVIg7aQXeOke
I8Nl1e62pwszWWdFn7wxZrwMLWdWwY50RxuIaJejZGO93AgUlkk4WrGBJ1xELoO+kUh4yQluCzWM
/C2e0o9SwSPingQuOlAtCuWb1LJD4q2cHdYY7outNqSRbYJgY9qvHQCYoUi9RiGkuJjcgHVbag3q
C/PK6NedJReFizsRSXfDeP2SDhNcXaF0APG9pVz+3To8jVkpc44IlIymNFwJAEmL2lmLbgd443NF
tIrYzU18xAtvHK3GjlpopB6xY0NBTLonY8bAJBC+BdRFBPMynkdht3RHu9oRRD0I94E8vLKXVFuF
MpCIFAh8xwXgyZfij+SKZwUy+ot0kFNLFleCZcyhv2w3VR5TxZVsn9eCQu0gi7CPJdqHl733cSof
CVcE7IEKTHxEmCJyWuOfrDKpxCBGFgUHSzWTKXtMwisQr99Qz8+U44s3gMu92bIcPaSo/Re+nv/E
oOt4YKJ9zsItLpsJbnFN1fol3uNp8NoH3B6XS1bEzQMOX358LOPZpQ8Wl0cAsB8Fxfmg6VioMsr5
J5gv3sUEZOPnmP2MyiWtRXetBqm6vARZfaHnvl8HLvYNECOW2BIIPHsa/xxTMT/CufhxJTfFe7Oz
knF9jbFP4sjbn2UNXObm8qrMxsgLgWShsoJ+9ZaT1FsETZ8CnfE1q9Qa9VFOk8T1fWHRVIzVfsb8
/2OF7zhR7rVrIpy4Gw4E6Ncg58MlVsvXKnmPB2+gLKS+KiiQ03JyVh/MRcByMHkTDTEykQd6WzmQ
0xY98bCKsV5so4yzmxFiTv4uzJuzhDp0mSI16GYUvXh+PPIyM6B5s8T6ayWwGtRdPSwMgHWgDh6e
gr34sN4UhSpP2v8pYSNVXR3jGLOhdn0tvWABc4SAJSuXOKSl31l3q2qWXWNEKuewXjjt2pMMQ6VD
+WMLaIxlsfq/RqFJbCqSwwfwmmnB8+0KVF7uBKo+c3YYnFLRRFtb5ds5J3qD0Imh43tE33AFXNGO
PXDvRMJ/gd8JQ6GtoBWCd+kdbOprSXOw5q/mE/f8FOf0Tn9nki7f5HVRMfOS5NQjaLCTO3ePpxAs
+AEzQ31WwCGtZ+0p4d5833ilx5JyM627N5wxKoNNZNrPER9nLVSQL59jdVuV9DAuVaFwXX0Hm4oy
L8CvhkFVruZ1FaEleQn19QztwXC/VMDqStnAaBHM238FlxK88R3XNvrdNTsoKlNELGKY9uCaTMj5
cr6mEtCF21cnFLnYefWwJ03X8XuO495IH+2/p7xwhNpc0eytJTMc19cT5SsgwN6lwpbuX42v9hc/
26wAUfKP/LLHDz/v8nUGB0FwJ8YXny8q7udPB9nO9+M3e9V3dKHX2cUCEpy8jdLKhDNZT+iwo87D
yc+nZ7s5N8d8r5y8GPafOhmDIy/p7AwkanrPgB/lkOJKqGL4ZuGdU22vkREDk6vCHmYfNLrMw6uT
rEHrXwLYVf1Z8M54MqAMAmIAvGQWv59dQIqG3326V5mUuKVRQEYopA29rC65mToK2ZWO4Fwfyy27
oYgd3M46goaXn+XeuK71VTOefZPPx5u+32YBG25fkc215rFwd9XOXT0ahCjjsSJzOA93xlOq909/
zWTKEXlaUx0uONfq2JsT0IVcXNibreefrX2F0n0W2mxQC7NdvHGnngvyHU+W3E7V0WXUQYHJDKW/
LAIxnqt07T2UUUuudchJRGUHZufV9953734Bd5CU5GQRsDR4Hc411w2o+0Y7wHN9JLct9m1RRVzB
RQwFACRFMMQKongabhN+GtqF5xoJZoYutWi8C6N5NKuPZba0BrCxmrnpP6Q50aKjQOy6zcnBAlUU
Yn8bf9VgDXpxt6KB36hBqCkdtm423c20N1u5pF2OMoHKmW5y86Q5JFwqWbw798uRz4XpFI5/6dnm
JVL3gGNib1s0t8xMrQUUOiNDaPIm8FXyO5+pTl4iiggbdMEXdbmaImxxETZX8NzFskqN/ZM8Ucdx
DdCgQVIRD077OpH+DubJMKdLSoIJAde0jo7z4V+XDfaLYILA8hOUV54Mvn60PHv4CXoEv8O1vCU9
/KVjJGa4N3c9dO/52xIqKcWYxi3EbzojauzIuAHlRc5E29D4TtcddPNh+Sqe0AJQDuLbnYCXLLn3
GbnDRuiSZdvhtDxsRCPF/IHbcpr+5fP30230DhrHtn6DlBDXSAHPdKMxSeMPhvL06cv2o5PK/ZHe
hryJTI2WhRWr3fpNV4oiY3gFBBi8vxRp2qd7UJMxl0ZqryG4h2bqgTLpFFABIjUEqRW0sOsWqQAn
fU+xcWCL5oMKLMs9kFHZ+0URwJGwCmvWBM7v8ZNMUDi5BHyb7tEP3JnjsH/w+2t7wudId5gIA0Xq
kVUGjjleAiaCADk084X0yJaJPGyy8IDa/p1VYR2xTzKXnVq/R5Xg9abOIWQpaQN/wT9liiF14vwm
2FkWKEG7eQ+PdxaXHdLlTLh+VBSeegA2meCDY0uoE/o3aGVen8pTDbyG8qRVLVB7i4GlKNZFVVKk
VvTgzfz4JYuUSONzrgwgAIdOuQWGEbzKVxPKrEuj/tGs0JWb+gq9MRRkhUWPYqOurfeJedN7gE+P
NgT/Vzr2QrdE+Bdx+mSjX0pDs+vlcR43dUzn0et48pGrMDm8t08T4Q8X7r+83jZw03EQk6KiINcg
fjveo9e+tALnPMLDWYgGZNjvHFVb/bYFbIj+UVlkZMoHZzGwQ7Bfz/k4JSaItjj5gNEHYc4fIf3z
x9PVylG233up+4pMyupAr8qxu2e9ghR+xdWriKLIo1E0Vy9Bp+vxvhQuobx7CiS6BHNR1tmhyL9o
qa1kR+tlO9t3k5f+5WlNPaBVUJYoM88tPFS51x95o0lJcaXBZFpP17PqGbowx+eYY/4vz9o/Q7fl
gBDUBar6cxiv6xZkWvyOyfvSLwM4qF/mPbuPMcmeVBKDXOa5xHadn36HHyyfB5FvoafNFFOU+/Ud
uRE8CsDi7nqd550gELmSlbultayYRFV0YTGkrnPqXf4vL3weyuB22fZ3uzY/lhOVngYE3eDQ33Ga
y+xKicJyBDSw36FjtGoXW0Uf8JY/Ra1PijittpwCJEsBVEljM2u1owSwVzqv7TnthHJvKH6YhBwn
a6wov4ejLBHpgrvaCI5/B+tKaKblOCJ9fD08Am98xizDF7tq/iqWwmcb3fuu+hrbUYKS9KvzRW3K
HopsJ4SgoqjvMAGNBW2ucg322d1CT/P5weUIT2tmSLOYFr/xUMY9fo/mi8TEaPJgt/n9yj1DY+cN
Cu+OGaf5fHnMV5Nh6PgrbrNoWRFuqGbzmX4TDEih7q31783dr9Qr3Ezl3UlWR3ptnBw7Z713hQAx
KmP0C5rRXCP07FeReHRAUIAOgQwaOsp33e5luPtQU1OOR8JQRauWtk/k++KhHlYOpGdXXoclloJj
+EQu0fWiSFTrSFlVguENFy+rgj+RFT+0W8Q4Q5wvJSYFoGesaaanEXc8IhrGsIrVx4TjBZg3+7hr
JLtrmxu7jqFFq6XIez3vGyN7/Klt6JYzzy21xP86DsNDToyz+v8QQRusYR9AQA8ttgLCpHBNC9wM
MmLrS6prbHDdPIOteD9KzghFNsfq3lqAcppdfYqC/8AWSWlp4tvoohdCi74Psi4f+Umvlj7v4loP
LeNo/8a5XoWVQj2NHqxtfzs00bv/eVYPrU6xbY1RlwMrUUbuUYm/mvI2NhegVMrhlQH4NagG8FI7
lKyfsaJgxF/qNYInul9YxNuSljVW2vIrXwbGQ5t3aGnMUSutnbEVBHs6bYa5FyxJ4+auXgb6yp2M
bHVWojj9DgchXCsQAcZdwlDoS9RSNqbx8TFNR6JkjGQVkKSfkBOJ3h+Vav4BqYAoCRXRqrda2lBN
EtkxRvYp1ep6kTS3ss783oVrEGl9pLJ+0GGB+KK7volEAw9fuOnbhaVhTcmCuZ9QxzMIyvUX0nnl
ARnV0cIHpIKaya1iQEnnU4vxXBJEy09V2dkCk34c40pRS/bPXGPtcbgfiQKBR00HbvxGQo/khxSs
dcANoC4dglrVDXG0AuLyo4h0H2iuTOOxKQbvlkZxp+dl58cqoN/tyGv8Fizs5VyL0EWIbZpz7zJc
QqmFcki/X5ATSumPsNQ5Xd+UZw7poLtDi72sDTnxUzZ6A0/FPk/Aszvwyiaj4gkGXZkcYbiFbiX+
GTYLoN1Bs8DzUF6vcofoE75dvI+ALPVHzTPOBTrku26+9Xf1WmIcCKGirEhKDB3oce8iGlp2TLG4
ETJ/dOD6Iow289sUGQefWD/WMF16Jmlmjj8jqlVLuVLWPnS70TW3Ds/FeAqIhacF/joZBloMSLwC
NK0tFlun+WCgsou8gCMA9mypJIRjMmnNwujphk7YwPov5pKVzex/Ri37eRW+AOZvYfbmsyhQmC4s
/8NrXjZFaIUzysoPnvIOq0oP6o00lI/R+ae/ESlIFWXbKC4OMMqoIEktJ2opxFrZjLGFiK711Kv0
A6ugSMqe4X188J6AWTy2n0kjEgSlQ2nuE32NGQ4Z+vbt2lwcOTLbUum6wXf5e6xgiQDbrzx+eL6v
PmF1hBJQcGu7FD2p0xpTA6TR6/8Z48H7BgEPVyLodiHB8kp0rDGoDyqpWMFy9wp7wPtCTXyx1eC6
pfE3i1Wbjk3Hqgintlo1ejlvqo5MNi9fcY0sFI7LO9UCy4wgDRY7ozhA4ZCpS6zB9bPS/o++IUnK
ScVxS4+smFWTapgauIxTsQ6qU2/gpTbtAQ1e5SVhaSpF/6RaBJUQzlDE/pDQgpQj2e4ybuE8ddAi
3JoE7FVI9cL3f1aepZAqOsOCwiKqOFlKrS2OtfGmokXsJzeNimtoH5yE1uMIVTCeygmV/QiiUDzF
x0nCIPptt3J+CI/5oPy1bHxIVHkV1TBa1CGLkSBXqY/ut0plvpcP4n1VsWJiOQ2WBBWEuNaL8Tqu
H3y/TGG5KyfVeJw+3GzcaJjF/7MsWWUO/vX1XQX2mPAk3wGjubbcrRme7Ubd+ltgE+dvGt6WRqq0
l9t7WBshBAPUuilKkDF+ZJRb1LXhOeEkQjMa59pBRVMrE/jNRxynOJ37OZg631zV8UsBgpLuvD2+
DM1vlSuzycI+YYLnM4fkG4Ahd6Yfau1G6lNU72B7VbdOSb7hDq8WYE8byEbMb52N/3w2J1+pz3GD
t1d7Na6YDdC3hdlCxZU9cyC4j+ze4IgRDRGoUPlZqRLCsdRfW/36+h2FGC66hSob9JS7CHZZgGIi
HN6HfmDYBJzjirmw3pm0mJqK5yVXP6qq7R98DMF8B8hEe2QD/ZvPFJblH6uN44p3Gx0rrubWl5YS
rzDUesGCB+4Bu2zJay0+plZQaeI76mEVAJJuCSvmHZIJjuRezFzrBZHtAoHYDSzIUwYsVRg/ShrS
/Puw8z8RU9YYG4VY8TMvo0XXSjZolFLCchXF4FbXn+lj00lqQ6vgglQXtgozGTiBwTtephKdwOgZ
21Qc8X5x75/xr9KwXbgI7aBaC+PbKXZd83cuT9RX0MwNRnnuh0b9DAgLvBA1EH036ADSTBMx3OHm
teojCBQEPUV7w2OuHB5TVhw/Aqng3ouUXNuFsebMLUwOGlmSfZRXKT9jrnLAfKQBWwTMNFD8R+Sn
xEVMMFSWvJqsauyd3CAXPSSXnXUhmiJrGvO0KYRtt8M3dSk/oH34LvzMV4uvsOtwIYCq6M8l0hhP
iQod47va5HmQxSZ1TROT8SzaaKbIoP0zDJEslnFucO0uqQCKr9kSLgaagiqVZfW/TCRT/LxSrqbJ
Iwl4i/6+HVzv7j8+MuL9DfjmAuq4tD1ApBvgndFcJWUUleDnpb+c1IVmF8Wia4mpHLz3Xvlighh2
MrkNoLbMRU9wPYjlVsRmnirGPNyMi1NIxqVXZTnXtjoj9LfB100sClZzZWgvdhGAbyUQybdUIoAc
xo+1TyIvMcXi6TANhxas0MRyXJQHil7PvxjyZKaQ3NtboBiv5SWgL+271p2MH44ZZGqbNnwVDaBj
2MP8NoNq5iElCHdk2z1/WHfjyN6i5R3SR1hMMXWJU9sjNuXrw8191kdwd3E27tFU1iUphqUOqT6C
PNak2OCf8eiL5D8ULhAb+j0DpflWU4F2IA/kJkdEfdxRzgOl+DXxHihJNrY2+1zGf7tP+S9xAmz1
mAR8uXcPC8Px61W+rIoTM5LG2Y8NXHCkrhhDdJJlsw+LSmz67XvjxYvJlaqaKaphO8kLDWX9avnh
klq1Cra+5Hfys3xf2ETrMOB/U/Hec449aGlvaYNd/TM+TMZ9R4IxJPcclsJL6Y4EuAucZZTpYjcV
fapkJEIVuKIhMNuUzh2PuH/xTZJy6IcFkCS6ir9gxQMYUnPeCuzTmikSrwz/tmNC0FmtnneZ7Tbq
FPVSNBrP+Eq9fhPIVVuMi8Y1cfYL1M7PclHkM78CtHqy5helhsgottDXdmfyzn7EeEDq33AP2+zr
IPQzkXt1c1DePGWhkGobNFXsTISKBIPv8KgOX4o9CDi8y2LUIyvXVRBDgt/6T08NUWjRd87ioAXU
Hg2Wk68JUtw8TOU2o0tp0iJr3ssHGCOBAMdp7uKKkYxBCZZQtSELt+r9kCIeFh3aVCLhzfUBdcyO
ZE864o/tWlY+MUSkM3XI8CUnXlJ0zJVB7MsnZijzbBCiuHCTvpcyVW8nAClpANfEjFGJHiJ/7laI
LXQRkXkP1lU23qKjGibcDSlmeRcGdfzQXq/4Bf1CRsqhQ0+h6jqTgH+p27Vz8ME8bIaE8NtJEJUj
sxSYfhPuuEbTZ85cRWNelztsGmfD/QtYwgqvsR1xW9ljdIyWeYUB5IFz1MRBGsboUSXZ/oouS4s/
Z5TPPQBSwNNUe5KL2iGRSeAT2pbZexe8zJ02c393vcr8zEG3IE7LeRuVOViEPKoUc2QryCrstDz+
dIHlx1Chm67U8AQYtDyQ9/GZoM6U38X4tWVeWuT0Zf+iCIhjzd3emB6GwD74+dFaTfqAY0WI/v6g
LcrrWU2TmYwcCRiswGHH3UM49hIKJpB2Jy1nBU1SGLqiRjqGJm7xrXPfO9EmvC3vC1ETaBAFcn9Q
n/YRx+qvl36ISMnCt8UHzvn2LuyM7LicwEtenDJdIaLZrANGTKoshXEDSjAeUCRD8fz2TGXSw6UD
Yh1ohobVWyLHJ2Hs17jN/efQQrJ9WNWZH7ov39Es1gXVpC5hcPq11okeZDf05YE9/TJe/Br4kT3g
0YvTSu5WcQlQFT6Vh6DZzJ0U72gM2KZJHAR0RiGz/FkhhfAGEpr4+7gR5nIUiaCUs+RFPCG91z1W
9NFAPmHCyme9lsmDRRV/06HxZgUQSOaLwtEU3x9+EUlGFpQ6MacKANGMZF6g5Eirjxmp3iQnhPv6
eekDOh5Gvsu+DprEIqFoMVnDL1d/18AYkEvj3cEex20fl8V7T4/t3J5YFLOsDOSTbvamEQVs7Tdc
2ll2fpMz/cTwfYtCFVfQ4BdWfTcBZ4dkhFoefUvzzPdxQB76XzrY0N9dxHjiHOsb5YQkt2fDD+gs
LvKKpyrXQPR0EK/cSq2NU+oxlGGuN7REbkA2k/Mu1a3G3VJf0QaLgA2z9LnqJiudnrjBKBwby0R2
uD1IejXfVumibQDWvwklF/EGjzqeX4koDujf65c9i/5rkr2lP5BejmTcOYzoODAKGqU0VHuIHFf5
i0bzYik4/wbCVnHuEb/oBasZo7iu565t1t76VC3BHpQu51n9/TGd2BEkAo+A9zNr3VCGuic84HqW
eivvpiAxDmAeO+sRj4oJcIF4nyn8xZ/GoIYkuGrudff6i38Zx/G9olWz/lKGnxo0ETbXMdkdoTE5
CobSybcu/AtD0qxUAsVpiAvYOAip8tDSkn4utEP+nWyeT3nM+jD/eApUwiLbupFFG9HunIVzKofR
dFVO4u+SeAASj0WGeldqKxZZ1ynwhJrmlRX8u4kStPao1QkA1jKlDJB2JDOAa9ddUl8v18dhdhpP
Fy5h8cpLnZOZPQBLmhlM8yoqREpVTGXuoc02uv7Hag3MTbqVD0pr7iC0drJWqsCWp6kOHe14rb8b
ZE0kVOVZCspImKo+rUjtsuTjwgxBKFCP6+xZd+0kMKeWfhIMhgtfdNCh7ACRRSXPJ2sckq3fFxuw
dSc2gqUvg4JfytvBBpLCEgN3sy82Cv/70/2uiapY9yQEaGrunIa6M1V79LTpMhpIpQseKf4rTcz5
y9P3YXhGearTsqdImBhzCrcDAf/FK+Mm/RHi7VJSqshw3HReBtIDRPpTdvFgM+ESEAXciJRWzNxk
dWF9T659zp7osIqk35dNWFILhGQJBPZ77n2Bm8Q0ef2Uc8kBk6kJoTQWY8j5QpqpRn93g15uzBfP
CoZNzKdhTi+32mNku4eF8WdlhWDihzhOf6opqITgb+yqPhkZ/Bm8GZawf+xmPgaVsqxz1uyZx6RH
+FHJLhNJVjwXTLB0Ncb35E/xDiXa3MmVWjYPw52FC5mzT1GypROgaGQrpsFr8gCG6Na/D1fB99aX
Y+IkMiCA80RcpdwKIlde7ea6ec0XulQzSAbYrz5SdXRFLsUUkgjd66ubZHrkpXVAJ9c+Rnszbpi6
UuCoojKgP7vjim/kgbryEbMvoXHF1GBfFjfTVsV+d4q4WjJKgWXFsNuRdUvgRie6iSPSN6/ISZAW
c79hnk5de7HA+l2BNTFiIQQ8iN4m/AdGXRoXcMYxpIqWFs0C0nWGIh3Q1uqWpgHg9/cmGQE8t0ls
6WC4XnbLz9N0XM1Zz/E/EUWHrbFGEpu++ZuzQrBUihq08Kbqwh45VNp48UB3UezH3M8Oo/uMVVzO
oXwUwcHxK+t9yfFprlUshMNbHbYur1sAv6gl1znUKRM9k8iG58o0gVmOx1uio/+PwhMLOsuA5It5
UOrcUvYdvXl6uDaJWM0QzO4S6StcZH0cFHspFDmfymqbst1Kfp2PFoJAS4TClvHjHzRvqh6DmoQW
UJ79a6d3fUl/Sq+k8fQinh6XYbQ0YZkNDIiZkIC8w5mwWRabcHAsGYPWx0YcxSaGhFl5eQNuKHgK
I0xXNBB0RRzrLqwe2GF46jfhdL+rYo1L9x2n0Ez2doUl7jOPbFOs7gu+SqFcwFT7Jod/RVvvahAq
v/cXBoRBS9EAMs/6co0U+usQesHWOQvVljCdCcERbni8KPB6IlfRr0+WK5NNTFuHlWAAN3mXKfIa
ewvezeVKhKFOMgAeefWKkPl4S/THlNWe6NOXeq5NUHBjcc/mVjslkI96N5tqdBh+IclVm8HoIFfg
4V9nt2p93s4EcntF8imozGxeWBvOT8bDlSFCfwG2FZwJQvjNvQJLnOjhIJhOChtp+B8HbXKHucA7
hfLjd0HjtHHFl2p2dnd08Rx3JSe03sunTVpkFzx3GTbUpHJt9+dKa50r0Ix+nNnRdeuPemqcJB4a
9Gpr0QM29UVaex8WyxFijhVjhwR8/wdKMrhKVViQVnNEeC9s+nNIUd3Cs0o38r1A5PQ/iKpP941v
zH923xNrwW91PGbVhN+n+xZTj+hqDoO9g98h0ZsvDR1/D4TDOqc/INzn+PyJ4mecIOWc4wQKwrBY
l1QS78OzadjD8vBcy40XbTykOEIMKP3Q1I2jR05u4nNrhQHhE8FmpMsQbg6MEwA35haRsUvnkdTf
2MvmAlM4jGDzanzhBxza9/eFxl2P50QWEe7pDYjy1h9FO0P/wnE8RPCaq4U6dsIWCl2/qPigaHwv
aTJw1bkjj/a9XT1KFzJJVDap0l5Rr7OrhvjlLqHUmWvuISuJBevoNGKtbmHqS3YLnj0SlFBdfm0z
gHzpvc3h71hGTbN2bDAee0ZrkEcoeZUfSf2wPp3gEXj/XboeciKYzsl+6iDVTVkNcLfvQAEdwo5j
/4VQ6TfTAHXWaL97ZcoFnLJfNfvpkmTm0B+tkdNFRkEpEnKJdX10zTI7X8U9Z4td9Vq/+udsDWUx
CL0hyZLTVKgYXR6pymyf6f0w0GRAYE3fCjD401OjDzjaab1lSuZ4c/eDf9fGnT4zxcgf17O7OpS6
cqlfTz8EoBcBHGwYlOaojCVJuN4skUCoAMhvFqPsfz0kU+a1dlglKvFRit0xTvSWM+W5Tf+B9dN6
3DR6TXWKGU4dT2qRTFA25XFWLEhNZcIhlO9Nl0GTSJ/3gLtBLQu793VyfkxpBPeaRBJuW4y2t47B
ZBCdsY6w0oNmQktuAdIyR+ZDct6MuuxN6hmxVSrFjKzevmbNbnrFHG0MI3dgBJh6vuEJZljmpoYI
MQwpB475PbPZX+dn1icbqMbe63g2rz+Reo3k2Hd6BEieqf5KNBf7nrkMZpN06mX80N/P+vyQvK+K
a1xdrklwX96nCJtsLph6fvQfOqQoI7iW1yCFLuG88fxbjg9rBR2DGVP04zqmOkKQbVz9bIMjgiH1
s+iPegpkYIr2lDdFHJJUgJiU8CcvN64yDzckM5cTznbS1UPbtdtj0ggD12ilrHJoorYZLdALcu6J
nnFIKBAJmj1SNND2i10l+vkgS7NwqGezgxZNiVvHgyw+D3rUUE8kko3SCBbkOudrWgwBByEKdnnR
R8BbQO8N+8BZxZpapnMbHlckpi9o0W6flekx8WWCCJ9h9v5MPnO+m4vwMNlgkQEXtD26+WCWd90/
eJXA5qX9QT0cU1J2Sl58IdmT38m6ZXWdwCgZbLH330UNcC9UStwmCm/Ya+hQxRqItADHulnIprJ8
Mqz/JW4aaUmsOOSl3E19nO8L2ryJ8hRqHbt26Kk2d6AbVidUxJMmyzsFxb4wJuZGSsA/Q1ZxHteR
bwHw1oMhh9LPaZog9/3D8MDMPRzsmANfRawQsGPAQjbOsS5KP0ijtZk9mm+EuVtWEpgNdBEWhuDc
xipstDPkPUhwaWkK2J6hqjA6wo/Fi4zQkvrg2Lahi+a7X90Ax3i2MT4r5Oxte4Kb5JC/rjckTsLC
9JDVOlST3auZNCCNS40vm3t3UD1wZyiN6OpO+L+vzIa2aZKLIxMt1pm1iXO+6h/RF0j3RQjeCinQ
UgtLA3hIGvpxyhFwgj83QDkWfh8OtEQ6PYZjnmjbyd2I84S2oxeA7vjwyzWLS5gdzQvTIY3oU8p4
BG72diGwHhljzm1Z06PeVUzsxrbXdWRl3jY7o+ds5FMf9nMzZP1ty2vTDHw9FS7zG092KGPUMBU/
W0PL4Nxsfsiv5mqKUCnEI4qrNvoNd4uFzHMO9ARLWvRMwXwnVOiomjE2ZSoiLGYvU9ntdgo/v8Is
oQnE4RFiT7ptOxzsWbHKx69qeaUPFofZoyx5Himm90wbgun15z9zCV6qRrp4fChlbg7lCOentMSz
+AJeKkk1c0qR8upU3IxnIh1u2GgEak48Px8pCohqnLVAx0cC4aOpKgOZ6Gy6qwn93jwIczAtrY2p
TmTXLi6Nbyz49aKJ4+IlwOAptAi5wvAT0ycTp6I19Gsg1Q3w6UR7LbyL1QAuoeuUtvhZAce80k9g
cHqwqeGR5wURg1+rnaHALCEkThaoo1Yrejb89oDiGVNVt7aW/52I3A1Y99K4Rg9YJhLPMoULNTIK
AlY4d/D97kURG+t3oViH1DGpADtXz/r42raSopWczyVkM496++Xv5TH+zyW2FNyw5As+k1QD7jom
tkkdsrGuC7ZRZ+HucbVzjBx4oz283EEYK1/+8wutTev4uFA9nnFq7EBef20LYVU6qK9gPZBF7bld
fRm6HAfG5Tgmv9/NJ5gsHARUWym14j6n3fjpHFc8EauXFOHKHkuJlpfY19/sABqKEMwUab7rw0Xr
1RsMOUlcId+4JM6raXM+VHrnwNjJ7L7IAfA6ohWT56zGuhgjDNgA0UHtFg7U8+0c4dgoz8S1rfQY
dGE5kEZJUBwE4Ui/6suMX4Irohxge3/TC9PGxLaBv/3GqadGljC/OSpiQUknAkQZpvv3UotS7juC
mySOp9N8CprGlubiVP4jJ176cfp5qobYUwJEa8woi8GqFh7uGAZA25L1eIdWG9l+j+DAJ+ju2wCH
PFrldbn3GDgVjCPFbs/Wh11u6e4VKU7qMRBL1wpjQUz7WOkD/NjLc9EZlZm8y/z40Fe2jCdnMR+S
EAV+ImKNbjff0aWMIYfvJ0NqeYzk6YLK0V7dzQ/M57YTJzrfkBcwyI09ZG17EVYaTwvzZsHhpuQv
CHiMWFfZl8BBrrVH4AW4+l/6ZqRBzt95v2QzAb6pFnrJfcYRhoanP3zcSUE8bZL3X6FXwb21J8ME
SyljeF8dquVh1Wvyf6rDiU2uUZCRuYqrrJWNZLDj90CgwbxE754Hok3QcX98B1acJu9Wy8qv+GMS
6oKFNEBnd79BwHkADrLodMi6AXK/9/W+N+jAgvsdAmqT95HlotwSdRzt1bu7Kw7WUSsJC5thY0br
7ZSLSEDbfl+eBrS9x6vaKJlU31zY0V8L05s6k5AWkAoMt1qafXa8UDqB/yE8XtNhSJUbk8LZl9fx
IS98vpJlnf++9kL9FAjtTtbWsu8XdVQqWuf/x13Q7G/gVL60MNr12Z+rhpMUcplnzXZHohgjJnUL
OHOtcnNpyEwFfGQR9ogw0btdTGx9suo1Uc5nyb7lYsT5z4lzGcqAb3+bDP9mY/yf25Mw1WA5LC1U
0qeazG6uR1O2lTA238hI1pMRoauG9mlm04e4VTqVmgXZW0ZhiIJ8ykPKMLMDhpa2YUZRmAIpvB3E
goI7r5CUgB8JWhtDb4bcbDUxrjTwtga0zmhsp4VPI8N3ToD1r0znOKgZ/ZX6tX22xaIorDeuHvV5
4tqYyt+k91slqG8OnAPrqNNS4EJ34km+qhva1HZCWyO5WBQ0//yFtJzWeo8kXQ3NatBDa/6ozxDw
CBIZNnc3LlSUGmUH7CNOJ9vFTJAodbEOzC6gm5FtShmTQT05C0ItAVCUeKX+ePfbb7EIBXGvTeXu
RgIsL/NE6uB/IyhUIoLU1xfS2pg9tC0s9DKqo/p310PpIj03h+1GEFeklFMrT9g29Mwy1WOeG7mL
q9nD4WmJEynf4ETPgDgLPKTqLfWt0QkQG67mLS9SJUESX/2F1deZ8mRQRVYWqQTgZD12pz2z+W7M
C83/Agb+Bn5uIEUwAss07EXs8n+iwXzkHPQuk3Ft1ug8cat5tQS1I3NmLyxMvvv8r7bJWM5kyUp7
yeS1mnwpj82DXIPEY8DrHbjZfwXG6Gx8a6Hc4CwvaP/sWAuq3LjbAzRUjr/JEbcCk32gEdNuc0Ws
TUm7ILxVyMKreEfaoNC9kQ6l24j+4TzUravVojCtoJTH2EggE+MuhNZu3BLlCfedDDqcIvNnkJ9j
hA9MkZANVnjBb0lU5Wvt2G/sjD4zzibXVfnaExuzY1Zq1ktWblW8HMRlPi9FDF4t7cio8ovQ8JQB
wdAzTuDPO2mdIfOu2mVy0Yo5BCZaLMjJhBr6ogkERnXxZ+tmx/AEfAtERkQ2roJ0ycD7sehVpi65
9aEEqe5Y0bI66WFxyVei1cpkjgNXbpDUG7YJP0TdFlQMGmMlnDGilSToOcx6wvCpj7K3X07i2qwJ
voRjinz7PUueRdCllb/2zAxg4IBxILN6ZbLY/OrajpJ2Zs84xaa6fphMEmFqec3VPg06qzrD1USE
WIesta4FcvwIVWB1EcFNe1Leop5+0yG91mEQQYFPnBVAxIdwhVkgc/9Ol941MOOCawHwTcG9ExKU
9U1l9Daw9MpTN/4Gbu4teNDAMPll/K6pxn95vEhNbqXOpd0NlblGITl6xcRyenwY/gWtlkVdHflx
a22NtILX+H5SWaz5+56FIHBNic6lDvaKXHuuELj4UtFZrNP2KFpSyvXQQjqIUwIxNsyEC0uBMk9z
4EOTSoLfocNahrIPrvGMTVOnLoUAFLrvI0JFpMrKHBfiU5y5IwOBrkN39s+QwXYFSzhrIzuxOp9c
h5wohEAdSDB6w3sarfYPjzj/5cYpvGC3ja59tzv8yJ0IT66B9cian5kiasxPsMUBzhsIaV6rtUAy
+POZbq5V5RU98OMEHaD5za949scokhG3D1P+gtjY9s2FIAUMbM9TUCJlxo4ADMGlw380WaTfMuVJ
LBx86wSCK9OuhAxb1P/sI3gUkGqjTAE8DxDEj/5dpkAeVdVDGvjWmQoWhdU/IPE4BwXY+5jzca8+
9cHpCXFkFk8uoEzC/VNxOMVHpRZ9/bv5Q4fCRpBemDvSV9cedwtj1Cayup7wjnpeM5faGlD6SFEA
YI1RigQii0GYpYUJ1DI/Xfh3uLxziwOfYfjKh1qguGurVVO1+8K5tqBM8LWVrJA5DFqYOFE5VRy/
UHVsXNILcsmSVdEzSJDu2ItpP/5uI+b0RRJ9NTU8fOqm8BDWv2ebBjeOAdpwZbqm82lJKflRQD3R
SYLmLM1KjnvyAJC0o3FJd2Yag3T3vV5eLWn01088z+RxO7zarQgFAIGyAfLIXi07RlbBf3q/DdYX
QaLs0Os6jXA9ZWiXh0VwF5GSBXf7SGskI0MCUrsvdvLoGWUnPSjhj/JtESvSm0mate9j+AfypeQ7
w2pnQwlcEVaeLU+5AGw8GgeidGlzNaMv1mKc/3i89YNKMpmBhK5aGh8l7oB8BraCI0XXV+ZfozY9
H89lzbRZNZBjMV1axV961/5ddTMuwwmtDYYRAVgh+ZKafAnSKQ2Yf2plA2/yEB0p5aNlvEeBcRjR
D7YLn6HNljjZdhqqIz9jZ2WPDZuSoAWtdnY7iKSlUL8hdbABfkc7GLbGTwpnAbe2qWYb204mO30V
CBI+QG4HdFAz7Dmhl1ocbvQIt+RMhy8XnLHilz8XumdEVz2XLEphU9vV0NnOnQV7iRKxy1rtmMqr
Rxi1Nw8NNOHew6FXM5/rl+wX2P02YY4PyzUa+YVAAqqqWTHy72nHnXTvpguGoqexu0ep2k9VSloR
VEfD8LfU+LqubxoAJXw/BBVpLwyMGHQXUV21VWQWgd66b4nd9WoqimM0hu7dvEeHuLc5I2CNyDyp
wod6R6mHnH+htliiM7zZ2ogkXHk9Xh439qWaVXk9D0ehR24aqZe6a3OlEQ3Dd7wiBLGwK5fi4KPe
h7MEC4Ch9fSXUqLjEyfAGLx03Vjof5Fed/DE3CJM2UKQgZZsM5eGS71qBCo6HofVees7remqCTzN
Y9wc2/HUtjU9QJnv4Vij1EiTahfNHLxu4ZjsU+6lKaiEXmXXsmiEEpO4jOseQv5V2igmFX/cx/o+
rKCFOvQS+kb5aml7QkId9sXF46ak1Fq0y6+sGlELM6bLsMyAewZsFlai5Er8HaYo4RhWhoQ25uha
8fnwCLHCyPZ8HrXVp77pDDjfzGQkEupiYe1PkP6HKQ0yGOK97VD9fF9Glbk5D95VnVygtEMgE/1z
3V8Z7JjOMkH80SWrZ5iYjFHHzSvbWrzxskLAiiWJM5bijW7MoNv0+NF8BrNmYZZ3Jc49MTdlDZlG
HByj6322Jsex8wTSbpvjHSpahe7NI6/eBBwvXDTnxsRe4Y7/IeSfJ+ydeb5nKaSmzWDbpkfcLZ0D
qS0/2uVI7fWz/XMFX1HwTtC/KlUPFhcyzVmIpzqiHaJoaS8LMmz24+HRHhIDRgrgb9StV4DzTU9Y
G0ffu5rnIrMM12U+Azu8QTgSOrue5iqZNKSwiaBu4QFxZDl1cVfZWf3wXN8QFRBKAu5W9hy6+XuR
/t4rFdjeLjK05T2rEtEGvK3ae9V8t4UEDFz2Qv1L5uvOVNfdqJWVrkPzrZGmPOafqaT4LyTy/rRs
VCFJZCDBohuUfKN5YbNmuXHCcVwysntUkdgL7E0m7gq8uYkKxiPwv2cTt+rezC+oVHEKd8HD82eY
k4Tp12tjHk/YnYqW5wsEeGQPpUqXbSmq11ImnjWUmMmW3a/Hea7ZDKMb8Sswz1sCEOLsRJ5DmQgx
Gole0D3xPfByVUcYkaKRkMyk/DT28u+GHtOV0GUGcj98WdRKRlpjLivjDrBAXBCkksTvJHF4KGbp
3BKK9dRrEAGw3RLyi6Jj21LpHlj2ExITFCBguHwBKbXURZY0Xrwd4Sihbo/m83aqd7WJuXTh3Ubi
rKvsp4AreZbiTc0yuX3muSdaGphUicAvlm5u3UBT+Mt2mGqegDKJkX35aQRaSX/ljobqNDLPdqWy
KhpF1nGdk9xkvPE2ET5ZDBVp2xGi5RYXGHjNo172HZ1dcoPHe6iiBjAabyEpl3LOl50PJN26XHIW
0HZFpVqMP647eHZCsElHV+UL8MVgs2SmTlNl+xXtb7vVyFz9XVXsBhVt7aKSJ9ayJl1eaBHFZxSk
l9QVuU8ZERzekbIn7r/ah8o5RmGh3kQIjWGR6sspq8WjooKJH6jAZUDk+znKHu/l2ebuDomuUQQb
p0YLLOfWL9kb/CYydm/oAII6wnHdBl9U4FYlFfDWukKKVpM9VlgsOxi1nqMjrZ3fgPJiRnifZ3sd
OBin/+gr0C743XCbLWb7vN1lWEjhryzBZoQbQqgvg/9ZPilEPS2ErHfZ59DokpzDNgMEl3wprbkV
nb0I067j72L8SvHl/1kP2WBuUdeyKT5QlVWBK/OaRnB8e1KjE1qGm0Hg32SWlCoyC/jG/CdcRLWe
aUOSkbLJ6hAn+O7YH+lcPQxvCU3iBeWnVyPhcmUdr2fEsM7r4Uf/gwLC4oSebeFQQAgaCUuAcJUZ
pRG4ocnomqGb9kWHkL7DiESbg2aD55n8/1dV6B3DzFSjWUpUsC2rZ/Mwn9fSOxXUK5KBrcboEj3a
ZukyL9lu+T+iC7oNZrinWJm5wjazdEJonCtmNSPDMNFbeIot3m0bPW9nOkxj3h8MGpQ7UFAkgWXf
65EE6ea3oj257cGmF/E3O8FTYuz8eHZCoOrqk1D/TrwegdyVYNiqlq/XGXDbUVzdUpjaT3b6Cdou
YYv9AiWE+CrDHknR0SfDERJRk7mYLgW/CMsSxQ9QDVrsvbkSZDPBP6rXKZ7Y7eSKpviGml1gdQuR
ojApjgaLn+aeXfBhJ3Zzu07QkEmL11IYRAoXuRho7OKjYFOBoHkxJm3dAciv1wzLNhUBP3Tryiw9
ikF6ipOTO2QiPb1kQR625eepsfvs3j3nE+p8tbBYqsAc2c7Rsl4iTXJ9AeeyYdzRAm+XzjySfhBJ
PPWwLsJ5zW51Mq06ZjzR76ZgjNfbZHVnFyjOBjwBG+WwO0E4JgavpD+fuvE2OhS7Zm0kJaG5BMWx
PXbpcpN8BN4yRaIqPXWgCenP2Va+8yeWRki9na3w3/QwzHyLqOWAuSxZINxMQP7ETefd4B2s3mKx
YRpvfDgJrmapLw3lVOPLvHEPUeBaeclYzPEi2WX3Ev3dZZ+2EorQc5j/kshHv40vBJoCbXJKrn2B
Ar7UcUjjB3evDTiddyJNnTM4UMTUgr51l+T5tEo0NUuyHmVioRdjgrX0nOrJK46CvaWpKpCUt2TZ
9taOOQltY2wJEG7uZQ7l5j6Rkq5PPf/yu7nY0bSpk/MhI4mmLRjhzmSVzNhTT7bJhIU0EE/IchEh
kVSPmRPaHzpNx+U9oeX1xuns1PWGcBJDQBPSbR/YBd2/UQL9exO5sr/h1IZnAEFdoPWarl8Pv6Yn
7z/Djbho63zUsYg2YtxGNptzA2JgkMmTz2FH2xgwcyisvHb19+H/60wXGYorAIt9Hvkm7GyLcdyO
3UI6jXO2Ymk35ZX1iUcKOtqEvBJE7fubRfhK9jB/eOifSkd1xhQnHyrS2eQcDCK5nFv381NOWGAH
jLE//nfm4RyHgfCicD15874vVdJDQsGft8QepN5WYahzl2C8CGdUFR4komJ3k94SmIashoRgJz1Y
vq8ydXa0Jx/Ru9s1H2JRhAZs+Mf37cGKrTmqTVBXyelfQWTnBPFUEW5srhOMCZsARX7Y1ifCR1WF
kMBICjpaW76gZXYnNrnGmBT7gPjVHmvFcjg3pf1inJbCdlnuYU/WzPt+he7mkvCKofsr1IGewjiV
KXqmF45tEXoC+RJKHQn1Z4R4Qqc1FVmQ4dCMeeORm+W2sZ6eYf4rfJwmaqQfkgRDbM9M6mX9a2Pp
kaQnkWXDJffGYlhy4dQk5s5kXY2h2WqkUkHR6YZdbfFHqh6ycoJO6P+n9lG09oWsHAtlyLJqL03B
MB8sUXXbefdqoy28CP8Ts14kFdt/1uyQ08JWhqkQgjyCOKFt3XRiQSkMi4doIOYuALmfmOY9xM7A
UbzNRc0LcI2a6jhPyRTD5eBFw0+6Ikwk9xotFh3naAo6cu/Kgo475mQjpn2Ebq+jGNdvyip1a2Yy
t8cQWKQ4JrLOCBHc6HpgZXDLpkF1kI0qvEVs7iRZUD8uqwKI3dxbKzUSuYd2aMQT7rkr+FFgaJ1J
sjNo7jj2y/YKWEvhbELY5j8EyyFfGhmLO1WL7BTVYbnmfBVAULdHw/ey19v8ZTkm7gGu8DqhHUQu
jzXAHB01JI7hH0DX0uOCqgOXulZwwFpMe+Ay92+Ao6F/B86O1PjkV92Mz/5CSxnTyx/1VP+NM1+F
cYtq+9gx8bptxVn660rahM5rR8EWzdj5DLQsXQ66RpwayTZVJyodule3DiF0BWBk/W9qG7hsVZk8
/Qw+jC8mSiytbDm/JpDFiCXe/VE7BOI5YDVAE9nj/RZMPgvhp40GDV0OkOBkeXI+5fpXRNG7vUD/
fLAGyzSNuuX0dgY0MXCgHAHNxf6U4r9hidFDfYgBGyzMBwp5IFnZKP6Kd3BdsnuBetSX5PaHWmue
cNX9U32jzg6wJiYEXaH14CdQuytJpeK+8f9sUaaBNW3tga59lKixyc3hLUuM+XjMxDUyCXdQH39Q
UvNvfuEyxwbxXvSNRVOa+1VuPY249XOwrAU4KthfUGiB7z2rEwPt1R1DbKeTZWw8HU2cbLzQVZyL
TWG11dN13LAHfk/QApQgI+UFKxLC9sOVtNydhbWYySrReIuzQ2Lv/ZScVGAwG5a6UKEZWzSgsc3J
QRBB3kQDCFC695wIJev/n5/eLd4+C+IxjY4/OZ1a7JUo63+7Ap1IKJ/Pu3PaZUwixkB8r+s9aHQO
dkY51tfHccPMwX+9iiu1pxgtN4PdgINZxkg7majMuBRb49oFpkCsMKhNbxMluYrfWw5xHySZkS0d
ZUBPsiG+pz+PtmnzfI1Ouu1mRpz093G+RmzsNh6+KtBQNzYhMr4J1BGHrfjOD3arzggE1KRLKzev
7lvu6N4jlC3njpVj43xCEP9/XXoCHTHTvE1mwBA2BVDVflMEvaOGJmDaValLJ1smHzjzJ5J/qkmD
XBCRDgMUgiQsQkkifyXmkfaE6M1P8QLIB4wmgHi5YBWQwELridBdwh4Q0VqnyZWRTOUejvznnPW2
qQymbCe7TyZOfBhZNQ05ZDQxvtI1i/UmE8fGvUfmuuGzXwkDZtX0tySkEuziDc9IiZBvtJcH/a01
U2N4ekGCrQNnSaASieI+SN3SgK7QasGlOWCf3q3o8ZwZUd8sKQwY6v66Nof/ifGUkoH6sn6Ry3OW
1HvsPP53lZxxdtCA6lDtu5yphI0xYS8O2rbfR+oZiUfKh8WUmO934zP/gXiOiY0iNW5NSHgzGl7m
5w8ITo+o6S+UIA2ig9BCa9k/ULHsS4Pa66t/vQH8//XfEtqoh6HGD2Re0K5M6GyxsjhEaGSGcUsh
rC/x6oDv5H6vyoy9Itg9MLDeMYBUFwJYKg0C06fsUMdllc0vtUhjFYkciKWnKB/q7jt2iC2r+OB5
BBoKpb/G7oQ6Xqmmfp+FUib1HidU4/kRrZmZHBblKoHFggy4aMNC0SfUDTTfDaslAUPnJJvtpcJG
d3bv+n5/ZpewcwZphXpmuLGEoqx1z2e2VXoPhUytIKOYALw9h2eAOUP+qA1vxJ2zsxj2i2oAC4zD
8pkW3A3lWt6kLqX/LOvrWCmfI2XYpx0ncl1IXoq7fzCL126wQ4aKqLAFY/q/a4wZVfk2GlSr+qFP
WCCuifJw/3nQL6UccLfI1LdpR5GXrEzYt2NoHub0cCZ+cnh6lxMSYK8H7n2yIl2fxDK0TVE/nBwc
qAXanbyU4domhYnnDjveCVsmZ+ImO6Zp+vZ7z0RG69BJXiDx8Elm6sdhkkPHfUiHBmUae5uTp0p7
72NR0xMGf81ihr/AxczfpQA++U/6eIo1DVS4XGrHjvsx9CwrdIsHDnO9H5DDx8NW2RD1UrHKXZ8p
f7aMtoCXrf3CU9pJKS90JotJQxQI8Ro2ZHHi9gyL1SNMwpralOQ3EN8lT7Oid7QIgovTl+g+z9C9
qze0nAjDF8w5481HBtu6G62CDdKN1i+weLxFBoSjD2HeazypkKbyWZoL2+/t6L6faqXD3Br9JfyH
L2NE/g77IYln6Q1H89Hf6LIFtPFqFfSVsDYoD3H3u1/VWNxLC2QdGJzu5pVI4Wz8nwMagrDjhgpJ
g4/hwytYv8V1HK4AFb1wEkyRBn6LPJG5ZIA4XD7uXHZWWFR2rhwJAcilVFAO4AMxG97tB4OkQWGP
2x3YDhsVuRfRXuKzYWGLBZipv7FxViQj/iIWPn6atXdncDgwOMepcxJcrXS95+e/x/Khc63A26Rn
G8IO1B/PK1k0Uk1lID4DJZgGmuIEPzDXFCUJIxobu4t4vzEnqRmLF3U9UsH6S9glKpwqmiXFwsh/
mVzp2ga1Fc/EEMqyVDK3/p5DfpdT9jThYunOGIfa5uaEYXV9ap2Oq+eWfUQ4x2jVegRJoHFHqoFj
4zXJNbT5l73Idg0tnx5RAsxMEVczdZGocOglj71tFqHWmtm1YxNWVBGDzXKCvPJX2oupLi7/ImDv
2y/02HZfrSX5mDMDmOoph3ZdXOAYn/N1+JW7IuFOqpTe5sKavYnn5SurgRuSU6cDrHExFg9W9oNO
Qs8D0vWNlU0fAzN0c//EsMzk4u+4Ee2R8KOtjfOMj6/2ZGmXy367Q+4tFLZvzc1YeHVTmoIf9UzD
NrNoJtJTcOGYtxrMQrxe2Kp/HhNSj8Q3YfXd9lScjJnFuwTJoN+ow4gEhEuf3/A/2ywJood4SqUW
5/V8I+FkRTKOEQPdaplBneOJgKi9Sud9t6sZRYv1gMPIIwZPyKqN3U/A/wL8hUTsr+6sLWWcJxcM
3Ze/5vvMjwzneBmfZHENpb6xxEyYP2cJqhYme1KCypZSOL6o2deL8tvjwBsyZaBUVmneiRvUa9t3
Csh27aSY57J0zwlKtJdTnVj7M6fJGSFXo+wL3vy/kuWBRlOuaVfjzIHXX8pGcjUYD5ivpiprs1gg
PsqL0IxHKZuOdKQ/1dZAF3/867DVg/4V8sgcsk7d8rX13r/SuYRSg/pXjoGP0U/xOKv+7EggHeih
lvx0PPpOaSvGGd2r2z5TB0nyWtW3irlZM2f8jICgQTvyhflIHbQkZJrOdSZzHQTdnR2aVbce+FUg
Tdxg0zLg8+4IlXvcE/l0+clmvwsQ/Znxilr0lLXlRWL05fJdKFriQyHQX7GMFOp5BdjeLHbKi/ub
eO9PmPUUAxjUOKMgBTEJZDIVLxcV4NKSl9Ul8VlM9ELwSt9cvrd5QH0Q7q/UZWHg/ShHrq8MloDe
vctoczwykkHd6y0nb3/afbOD7299zeePr04rpNI7R3LK5snRxKk0t4PRlYo1ulhM1lQ/Rfsulki3
/3M/jiXxGcswZDRoV4FgvUB4/ZIJzeDIfot1N/PhnOw5ijKV77RzCWtlpL1ZR14l2EdDTwR49MFr
0KEEshI1uttEP105fQTgBAjxIAAlfvpnKEl4ar6nuH0YuPB5gNHbxPIYamVFx9xBVKWkm9P1eabl
xtJrkGvp9oZVKb7i1p5bkwjBE9cu1Uxlf9J3uiwSUN8KzI0Fm6vtRjA2mgZYEpNC03LQzuYT023b
boU4teRPwkEiDGQD0NMAn1kBOv0d+FAKCIVsKNecxiMjMG1EE24MOJ9D00kVZ4q15qu6EGC5LSmC
7TPNxdiNSJ+1N62F07x5deYzazsKmGTAmMGlUQodfp8Gx46w40dC90bfKgTvV7eIGOcfpNyCSdJr
mQ+0WPhpB2CHC3dQR0GcLVM9aAT4j5WpPmdpLytA/P8c6h1wRo1XWFzeUh1hKgh02TIBtHZJ0s2b
fNIWYnPHOzNojb8svFnCHoat/i+NChV52E5wbeUr9aQ42cuOqBAhRkvman8Cs0C2XzH6ynhKn/D/
7sYlx2VpRSzbcNJYTnOvNKL94mmZEiRIB0gI/213mzQ2Y0TNuM4RC1GTKaWxyAunJF/E5xDtcehk
3WEaAjgyiSSaxx3g72OMw6GcHQQsxsCWYcNNJmL+bBpiOrPn5t16cjqXaPj0tuhQ0V8ZPVePB3bL
yXU0+ggnEORldFEnKrsKmqp8xNkQbKZRqtWclcI7KnC7xsu78Q7Vaw30x6GynFst305y+f5vXg+v
ktFCK8EIVs0WwYTsCdwSFHR5ImqCTaFkHn3itNQYt+WTpm9lTdrPD1lPFEkl5GfbJbACYoQYARIa
IL7Uf6I+oKGvA+w0qbwzyYNF0Yqi9geLlqjF2j1+WK+h9mOwVGaYjr47k96bf8RNiKk4HIpsrkSL
Pb0gOF3q/rb5zzuQOrEzsdq8aGTmftgokNUvTFVAN4DiSwyas5PN/+O7cojatpyTG5Wvbks+v6+q
YJvRI83AhItsbz8N1rM+sx2GAzJT1BrE8yJpoAftF2LXlqINmHNDL3IKAXrLLyrPRoAFAZZafIdY
YkiO1oRykbksQmATjpFVcYYZWf0hwut8wveGQlQqBhIre4uAxTmjoUbVu0S0xBbZIDOml+IGOuuz
Gl5kg0jjVxmwAY2T1vlnMGE/poaV5px/rGx3BaeeHIdMr0Iq0eW/AXqo0nNl2GB0IOtT4t7cB31E
GEdTk+EWOLAvXB7Oj3X4xjg34DXXWPK4D7zzKmrM9h+7ry6MvJE/HxgxMgc4U70nQU+pgPWoBJqx
T1zMXVOpIAKcOg4lVTRyjQCrYzoh60emftpMfi3cgWet7PDNyoHPhsJUEraEIHdQJVafwD1LYpF7
OZDqOvn4tDFohHVQzijJ/hU5zgfKeT3cANWm2zK2nFl3SYLhLfUWctJowzHWaBky9L+vE21nxAWL
Z6z6sAAkN7UnEQlm7SPL0wcbskdGvt1U+aNBDHcSUA7OG2Dtbqkttt5wECLm6C6+X1JKBhULhYUh
wP+6NUVZDrwhE5wSYfHVnUlMQ+8Ssa0iiw48EqyEHPXW3BpwEy6wEUB/QRcJEBxkl9op5mg0ewwQ
qgjuBkPFNMvAc3Vxx5hOxxC3rzAfloajC2SrjNSQGhusnMIQk+i+yN/KU1aoheKi48f8exnObK+y
tPobL5H6xEVtFeQv/ogS37L+/eXut8A+3nLASco1uFDutrndO93KDkgI3E72W9edk7wwV+k4udGA
ub/wnAR377nGFyAwy7BAO6+E3PZbBTuQnng3nxagzlLDiFvL/8CnI8VIlFEfhuv1ZfhxiwN7EFCo
15l6XP9pF+oD2PB+/0gwzeLV1pDr/I5psARExurfi7uSgkSIunkHyY9nqWMPAqRBimu67OtbX3BK
iblJKy5umARJ4KpWVb8ic0bEEbm4LAO4V8ysZ+gFPnvqMG7nCDchcWqPFbzb8OxFY17VzVRXnqzA
l/zZkwoX1cK9lPLyWHU7MVPy8NJ0xKVsDeiFy8M8XXv1UhABrAg562h5zjVZtnf7bRsTK2oZO9Bw
RCwyqle6wUOhFzpUzrJsJ8q7eClH7gZcjX3ofirvl9wCM6qhtL2HLxsXoRIISaPqcnb5g4nKIVl6
t1qUp34v7b47btKSGcp3ps1KXwF22F8v0vclJebAwG8Fot+wV6KA/9iFlvVV7/NWdOWlu7gAMG1+
Q3Qr1eOkWrYRd/fGj8U4IhnlNsTCLLmK2I0TMY+qQmurQRI3nQvkZIgfoE8FXSrqd6P3D6Dhh/2r
7zckYlN8FdB5NBt/yauZyhYyU3foC9RGiKS6n+jqp+31+U/rHfwKZ5s4rBlCYIPx6ZgGLpqNPy5w
enr8/jWSldDlpD1MoiTd5GPCf+Pxsz+EZTChs3WoqbvWKY9KfLTR56DDKg0b0e4+hEO9vvLM+fp5
olcpAndnjHt5iCX/bCQA5C9LQ7Baex8Nh+RDnwgGHHXueiggsR/lt1gCkHZpvQ47ywXQyakPfRPj
Nn66/o+9LzVdo7gf3//M95Es18O0+hhEU1w052c7Jt3WqlNwwtNfTs9XolmgEXxG1pOXQYsIGDSu
QIYHxG4ku0CoPrKADfhNagQOjkRfWe5bLeoe1jFCcthdgOAlNxWDCT7r1KhCBO4lV58wukIOwpVF
U3/tUBjdKTklvlDRIQUVfoiFSfW/XmFk7U8aEMsc8UEbioXfSYPd/0ZIdl++1BXkcIzN7mZ1XYZI
mBbru/5EjwtyGYtndDJtRtwy5b5mPLAfZLxYwJ2Y35eqDpcxg7BO4es/cNjbGXWNAfb1AZ6VAEf5
TY+ZIT+Fa2McTRB7tXDpHz5fXLe4lHcCsZIY+kmxWEFwxKSVn55q1FlIf/Uc5x7qEA2W3jAmTLda
tQbJJLawdZgxlxApky6Ac0/4ddgQsXF0mEZ9opc6B0BgSI/7uwb+cVJw03dw5e+cMfH79yQynx+G
GcOid4o7nxbh+rHn8Puk+FttpT+3v+gLxnQ9sB+5rGb4KnPS7IE+s5sW6QKFH0cq7Vtj8zSbO2/W
SSrKw43TUXxhtV0Lk4RdFgTyOOvFiUVozj/SbXDSMAejPu/eLwtazuNqt3rsA8soHaWVrzaj6mER
sqBGkHb+702IFhcN06KfOkS1zAVxntXRQ0yXXKGxjMPJVFMaq+9BQQBdJlc0jOg6W9cRO6Vug6+e
7BsqP2HXXsXMcaULLYm8N78YOYq47mDRsZPjx+dgRQIVe27GP7/cYGDEekq5OpiCPq5SUTzP0mT9
ToZYmh9ebHo+gDjUR3uXzK/fzwDEexX60MStJ6EhskdR4Gp/mllDqrd7USJmBx+c5htHzjyZhPDI
O1LVjVJyRD8RtcGdZ7eZGj0pEXXXTqjjBJqzk5c/U5ToJWHQcFo79536861xlJApYY9zip19rneh
PdTQJlMrregrDRJ9AfRCGEQpfK91jsScC6DBiuYHXEGyUFQOOsL51dpD0kGqrFrskdIQZtwuL60X
UAAbew9aoeDz496cPCbM0xtrDJu2X95rUIFtWS9IV5DpI74Fsi8rH4L+8aec9iZRI3sNUlgytUFp
Cl2qW/CbbwWoEg6r5fMCrkgKo7ai906uLRMB4cjohhOt9QKIhIg7Sq9eEIs55Pe8eLpCkEWox5+G
l1p/9Xn1d4+bEgXgfIvZrr0A4YFDjUQQynzXHqC4hunXZ4rhn3KCG17GvU1kZpkLW8+Ca8kukPcV
aPwdNFzOzRLirPP02PSHZJ5mBCQQcsQp1n+6vCKCP30VSAQBhvH41OKohVOnn5AT8Bk0a7m3uPvT
prrFW5oiSqJx4d5g5JqyaA50ED3mHwDEhTJ8kkJ9+QfI8ibJjBl4YMoc+yT4ofABpjm6SJdArLQu
yJvQNDgzWK/oIWQOKoET3VfP+2ChmccuSn+D5Uj+7NxP46vA8+cFb9mBtIaWSeGsw4E/lOymNZLK
KpaJhzcCIf38fTgkX40hwN8X5d3qruxvFMS7njIli9LBE0NRL+fEb8QdapsYI78Gfvbch7xYGNQm
m9PS2mWnYujPdZdinUWpabSb2E6Zgi6ivO7kKCM93ygkcK9z7TOjjNsiPUOEM/ky3ulbFURABtiG
jD0FStUpiySKrdTXLILJRWFLqJi4Vwq+J7K4nxR7wFGmQCa+cV2hRlijzTy3oXNSKb54zmG/GdeC
coeSdNKC92b4gYb/EAHGygeSWfwdluS2CEemBSfx+tTbfdXw8JYYS/syoIfnJbLrO+ctbHJk/9J3
KsivSLBpGqvfu2D/89d11Ndw7tmPEFETau7EwlTiY7MEcjdz5MC/PE3eWwZlk+UNEhewOwI5d8LM
9u61FdsSeK5unRphpsbozTdZUtuBD5ILcve9yBO2z2/kFS3uLZxEYkV2skb2hhFgNbPlct3cfpx5
1In8lJA5fEhPMj86f/kzMZhlaYxxT11+EZq3jC/i8g55fenKKUOgrH4HfohwQ/DWYaHkc7d4JMkc
tEAkHsfu5X8G0OD6h4sxQQVkczACIXg38tWRPzjsBBqSM1FZ/WrEkznYRWeAUIHGVNQ32qxXP5q7
sSL6kmj0lllUi14QAmcjGIgsgvCrzu23DtBAXWl6ChzPb/V7a171DdF+xbVii6jho4BPkdCD3WvA
kTFf4av/PCYbXWBcN3mqX8dECyRgwTYjCRnejzGulQbqYIrgbFWJlNxU0I5oWd7bIH67b9E+lkNM
+jkp7b963MAhiJ+JO0FEi3zOBn+TvFaN6BXRHqidgWKVOz7t4ctG3AGoPej/+KvuH15FTF2WBn4D
kf9VRwePxMBU6+77W+u9rf24/zyST6B0exrdGhTnTjiDKRWt5Q5oLdN0y8vM+O0iv4ewMPoPnX7d
BSEAei/BN+qbILcTcXd3IAN4xlkGCCOmOGaAAttc+2nsSUTZ8hLSoRtzgf5PQFw4IQcpkbwF2pGu
jKbIN8T/eJRzHUCgLerj3GBcvdyeTyHytkTfBVR/68n6xCBV20mV0zc2KCvNM0u94gs/HZCU5800
YzM7KmKbZcWGKn3fZQF1DSJSEo+ntK2U+1KKxUNS+0EAGydTq2Fv/SQgHKYNU5uUKw5Mf5xBxb6O
4/HaHMjYAdcwwx6ssBWgmJrGpvU0r4utFfpwPbHpZ5uPY+piiMLA/bZ0JDxT+HB++JQvO6vfAfWa
OjCSP149QAvQB4LT8R32xfVDeat8RAtOAwLJjsTUT9jjWq+hC2w8E3AavB2tQyV6LOtwibLRJS+s
tHEh1M+TfaXXAIXuAW0prSWIHecnRJMMq0MgJpzM9jy+5ppYHZU/NGTRIkFjnPnNBhGZQeJ4fsdP
mz7glEIq2dxKEqq1iK8X3mltxsl/L1C0fTzzM4uTjy+qFihltKBwG+USv3462yCH5etu5iDdvDEr
K21zV5p2R+2636xWzXEk1vQunJFtgTqHa7h/gGDVYkzyUsOiWycbmmqw9SdTEwa3F7Hf4goD/fQF
PQba0MIo++d7IjcjfQi+EBGrehiV2ZzUeV+/KTxdd2TtxlZPAfnm2o8pbCTmiki1ZDsWCRxtjzNX
3Si4Q/mUqDc9Si9C4FH5+h9LwQsqeNh+tAWs9YciXV4OMnNaSfddckZqZJczQiDpsbTbOaJp01qF
4uXNhXY06PojjMV4/m5owZM8I51mDLFa7Vr8za07CiVSqLKkY5DbfHXSwSOh4NUGByNWOVcPgRcq
HmCT0qP5o4Sv1doALtKcLCbUekFsvrXRh9T4e/YAg7BI73iLvSLsg5FFzoDmCvjeRwguJCaSBjxa
C4Yscxhi3FA2cafN/rfttlu8oJS1f+b4dXgoPcynQHczVNEddFIuQ5ZNy1td0wedZYswaFSxf4hc
naOJkK9G8VKQjo8jqLUBR5zDLIoAp315sgxNDXP/rNilk7Phw/1wPonyX9h2KkoIW/f2/wNjGjTS
p5c5c+RdoCKyqbkZpT3jOOsaQ34k6FzIpUImnDOlGpy3RxXVWeIoUAdk707c4/e5TVhxCaGj3Fz2
Yq2GZvhFb1KoBxnydTN9MFSYWR4YyL26semDwRBJpTjEaXVBU1QU66DHV6+zFb+5CP9JqA2OKfVW
FW9WscUrgZh0oQHkI04GiHe6PxWM4zbnBoSpExZUUM5LmfGH0N/zgb17tTeXDWLmFIP7rQ2bkKE3
jHkRqTvgGHfopwlJPc6/mSDjNVWAWB8KcDxkC+kFpxJwllxbwa8gv1Tggf5NfrFC8e0LOD+FjUUw
Ra0HIgGA7+/VPDFX+8i/HhJHzXITlzVRKhVM45Jv5TY2NPgsMqCfVZZI3LSaxdk/7f6hkfmADRkc
z+KqQb9sxUnqG4Fcdarc41y7j6I3+2R9Wsgi96dDAxa3GhF6ThRK1TvxtHj75MB+9Ei61Zvq5hfh
f+2McDkjK6gURFJ1EnCF9sSSRl7cVA/adFEHqtTYJR9lEogHJoaBpKXHSw8TUw/+iypMOJ9xPZ+7
XFMwh6KUvBX+hDRXSUyUY/Dwq8n628N63IH0xW4upsj+ojI+fwFFaDvCVCzslMfEmLsTAaJa7ZOR
Ne6yYt+WqOazGVYAe5Woepeqm+/V0ZbCeVOafOg4GqJhBeKIeCxMlXtiH3dc1Mzhe9BrFSjZ2wW6
Gt5LucRITduhNtFe3xlf6tVsyYFevgwnXhJyM1MFU++UITl86hE9oyBvyS6J0mc/YcLl/kCTjgDr
QNxup6FswYoZ5Vn0cpyD+AYvKw9UQPgrpscTqlpgiwfs5h5ArcVxv/NSMtry8dmGktuSdC1zNAFC
cEe+TrpI+2a0WpgKD4VBAZGxVNnCBXprsRM0jIa+7RIS+iWiAmeFDoQ6OQiR1mBfCOufm2K6/QnV
c1g6JQMkM5O7VNmG+Gb/syYkPXfE9blaJobXEhUXLIlKJ6IKLbD36JQM0QEByj0Th/27py5cUCsp
qHkLrDD2cRlAYrWxq/cE2BuiuzcZWpjvIfYhMoysUQIG2ParH8+aWwuG8QUdhrYAanG4CLHMctPe
CNfMOZ+mb3xKaMDC9+Ea3Z2kjFEvo2y5oe1LiYSPe/iCCUD3GRopXWbUiZ3p9FCIljDVf0F7GjAg
+k1mLdJLvQCmM/2jSwGCCZn68971lYMA42yPLRHo5MCv815FcBYLwgm/Hi1P1DxlG95jfeQUNiBd
AtUoqXMESJhvLj0KvfIWyS6vdkFXt9PBpUx0j1vtwJZy9Q8NuzdcP32EXvHBGpC6cPnBbIonSOLq
XsYRQYFK0CNG373XPqGT+Jt7QhP8tFGoWlzAtGz5fgGLqv5rxlI14zx2bS4nTjB4cc5xYbkJ1hEa
ufLoeX7DnnFvRSMQasxI2JO03LRfjIRzwmnDx2hUDS72JV8iHvqHFjGM/6vsjEqT/4KHOvUD/Jo2
ir+dKcnvSk+Y095FsC/6g6mua+BvXc1edO0mcwyHKO+zg79jv3pFgBw98Ne+tTXVBoR03hSULjNP
4E0QZsnU+0qjoipmtmASRE9DqXy/C9bRGx8iRt5tan3aqqCZfniduFkM3EvQ+tF45QgIw12qOKB2
a3UpSr/CegGJ5YPU+AedqzoBRrVjt9j8T+NH/CoWBvnT69PxBqQPyLYun6RkSG1KvGXnWCITvujo
Oh8G84dW74AU8yaJRMbD2co/+dWQCVbPigMBwA2wPzkn5tZJ7BYBwyVdBv1rin63CnE8YRFb/7Qd
OgUZfgALOGlIXqvjhvRiCgo1kqNDbR4uE+PHGwDnO5bHRwwbg5dsHRERiim67kbiNOThQNK3V3Ka
uKMkDhQrNVX15zgUvrXVrckFI0W38zslEwD1F7V4sskBwFPSKqMGoXNk6G5p1qYBJGr2BA5Ieopy
x1dodmPx6c9hsa0MQM+6F6bFi2d8/1G4hBK3cqoqnx58dpoPZPRY6qjYZhLFpkNJC7LA2qeUnUtS
n6uGeNVrD+ybMpCymuUuYhTWKQddo4hDbdMrJnVk1bwKNAnByQUfCo7RzDQFD0laqUo0TFNcj4+T
+7LvZt8aPx88ju46F43o20JChPExFRz46NM5Q3MjHVp1szouUP6UNJbl4jyJiCW/IDVLKaLN4voC
NBr90W/EvrPsv1nIEM1xLmzqW2pVijfcEuCAPeC2MoJM2rG6iMxCYVPmkKP+vG6aE22xYc4p62ZH
BSIodQVpvg/xPpeFOPgmEaRnA11cVKGzamG4CYXk0fATvc6lCwnbFTQySiYeoFhS/iVI1E2y/zv1
xs4IXEs9FCbXDxy3TDCG86NBvL3Wsd4obfI/tsDMjELSCATqsUhPmqY4BKACLFsJHjTCxSvblWcU
Y+n9QlfDA0RHZx+DXi35CI3guqGLJm2sHU+dy6ZjqQ5E6KoefpZNMcEAKMPgeJBGs653WfbvAt7N
F236b+pP8D424TttBe7cs96XxBcjFQES4DaqvjEcTfV0acIB/QFWH2rgpgasLzRrgfmI9FvIJZf7
ECM6gSbapheVT5psye5or65DIwYWRExYOJduf/SR6IQlGuwuifFl0ccmFzdsvHkOO7SsZJV3pu+C
GsFOVaFgqjAEcDzHYpLb0E6KcHmlDVTgOwdKYZL5Qo/aIUyxMy/nGUMptAVPM7V4n8h69L4HDb+4
fsSzmA5cNvYnJsq03hCNk9fyt/jJHr4lZO+xLbiyoo1vtTPvvZl6HOKVPdrao+c/hYBC0zl+CJnn
WUGpC6KBCGlGZMwmX+R9py03PL/q7Y9YDqnSLdC6yCxeeimzi2avWE+caoQ6WnckQ68mVNweE6wC
EYfK9SPEdwPM1owpIU0W5/HzWBCESLIa+OsTXSwIVwFlMM5TIZ1v86pSn69W8rgSg0MtUzYcNj+8
Hmrq5Nja3GLfcSzsLhNtl6amJIdRWSrZ/ivTEBR7n47Y3hsVBPXEzYJtMy0ITQ/3kgNXmMsnTGio
GbjbvFMdRPeijIQtBawAsLps4WfE+GzfEIpvKXL38I0kFw5wVh+IcKca1dYB35RwTYTGbQ+XJtYz
SNNGjRwKT+jErsOI+ZwWRmuFUUHrOQLtuwdYUNsLwM86dGrsnN3ZqOdiWSbqBhNIwi7jLlZAxBgB
E2bisQPgKIh0HqFFkxJcWireFdD1j2/lW/pFnFOJeP55Yf8xKZTOs/vgCUNv3ZZHoO9UqwAibDSX
aS27WQas5LB62o+RvR7TLbTaV2RrBXVpRR7rhcgLxGfjXognEoRpkrIgE9sJPcmlc61MH3BF97gl
FQew9wEuLG6+CAessp6C5xZWeD7aqgJs4jtJuER67hKMXMnPGp2XIeQ51KTUYSHW4xUq3YWqaah8
vN2DkHXtK/ZRgOmeZ/hOVraSSLMxKfkWVjehX52ESyKqL5OCjtvEDKi9+yW9woeifthT4sHQWzMG
2JSKGGgptJKkB5zCtrc0t1UrqsICDd6W3I197epAMRlzQgxf/cjMag6zohv3evdxImN34A/U/uCn
UvmlW9pMxVcsZ+XZPiKuvx0fUcb4NC+Yei4dQdXR0FM5rbBZMoxfDGSPjTkv85OygHSMUlVJXvu0
0tBGeyktZDT/b/VBmEl9Tj2Q80+sG5h4v6qaF4gXLwae4lOTL6xyz80UR7aS5yS2sGRk+DrAEtML
11xO4AgytmTiNqhiQMoKECBrHlc83HAkTI/KaNXN2EfdU4z81+0tmAm9wSOwHKUOSBgPnFtbcu4h
VfwvAkd9NEJtTjMW57+6nAMhnuPYuvyJojVG6CQEhGXRXc0YOw9k0LMLVQwLPwAOB7pkcXBuqYgb
gNzMD66RHXutBUs+tODnxVsbkCdf3ZtzK9D/xUtu5jfH36LtlZ0cjY10Wg0kHWoA/uZefYT1zD+i
bi47k45W9njfjUR2Eq/N2emx/Xrm/RsUX2VNZvmfXWJbXa/qaGEYQ7TfsafKpBMlQ5ijAG5Cgzzl
4DnUje8Yafu61XAD/9RojXIOdDF5cTh9gxOmO+4mmnxuRVw3vivO3eKM7MxftNeBkiN5L9Jjb/UH
rjuRaEr7lluzBPQi0q7eyNSO0vKBWUw6Y+fNKEa8ZIo7FkohMbNAe5iVF4jclzVM/0ij0lHpablH
inXxl220UHMxZyyW65AHQKbQWgGTKrPPElTGg0QUwTmJFyrfbdF3DtBVLjeswYjo+YUYYgTfhQNf
hteRVQAxwuFUW046tXJQe1+pqordfIfc/jiOmBfuTujyQrmVu+XV3cXs1L3im5duY9Qbe7iRFq+C
9VI7YCL8Ua000O+yG/CurZKwnMzGhVKiQHLwapKHDo9yqDWpzRn+A4MCHOpZ3SjbXzN9wvWA92l3
R5Pbthdpj5tEjTsonGJiKD1GoTFo6ZMNm1yASjg78szvABe0hSVCfFf6OuSc8oYNAuFhA86VhpkS
QYliFIXja2a38udCpMEHqz/11ojK3kFlKB8ykO/s211CmiyTo9AXvuo7KT1SwYjfPoxw0BzUXAzK
lGzMIhuFOij0ctlEVI4wLtsMmIkUgwQgUJQio7YkxltiOPigBfkGjnKLmPgFGJz7wMHszdZI9z49
FTN7ekxGcCTBRGzbLtMvnDGatXoRuTZhLvrgWINsrhynP3P+uy6r+rtbd3zYjdysLjal8qOs8aVU
Zh2Dn+JsmV/jlW7965Y1y5D5iDzQWIfzBrb0E3tKbB04elN3mqB+vbgrEbSVJ6Xquq9t2ZekRPgH
xMQ5baNa7niEcxEjxLwAZxsH7jstIKrDsdd+t68jX4D2AmVajEuWmvEsxGOx1/eRryeRLAoa9WQN
NNB9TdT5P+KBsIojvMlJaZtA+VLPR//UbhbnbdZfFaX2hYM6YwtpxtDFGPNoVHvuJ7TTGbdNLaC3
jZCXjvT7JiZ+LZeZ7/ucYXWu0YiQZk+3VkrChFrm+8tLaFSTHeyWj5FZy3db+PTIdmE5coeEME5g
adnkt5PS8ttHjr3F0dVgEPMt54e91Zlpf5NFrkiJB0vspVnQ8WWrl+FbUQOU0u3CQdQFcOkapuD8
5lpwkJtcMoNxFkdgYHB5tHdM0IXjaeLmgEA6ef5n9KHhkTQ4AkdqxroAEZvKI31DxJBYG8beTQrF
CGuo/gS9Ch1fdsNc3VwY3YADd96yVvvpG7sA56ABMO4agUkYyLLFH0xO3KwEdiRxJe59eR9XWtuz
w6U8RnLLHftOen6FbqfyaFIkeZ4Y9jhwtpX/hZGbL8h2J5pcfxRDR4h6w1bft9rGdtVtnj6nYLEM
cpxTr+tgNYxCfuLZeZVHNz8pL2QfjilEnzvyLDgUkMAk3N0L2hfo+hdiUv98V55rEoVeciJx2ED4
abMUpjfpb1yyFemq8iMTrDmoj0VCsime2yjtlDdYTU2fUQFUKC1IcpygpZ0r+shvRdUQqzK23rQ/
c6iC4eY0pM8hR1Y0i3FhuuLPPcPcPb2KPtHKTMXhdg0aYTA+GT2JXgUjxTCCDpFxJUNRnKU6DfUz
i/WX+y6pi3FJ6C0IlAqMVj0AZgluCribVru4abWIAR/dTR07cSh3eeJiuW3ESve58EEHjZjT9el1
5IqQR79Zo5Z6TRvPsWbUhTHZLnBalCUtgPQaDQvUT2iyLHa1E6NnP80z6d025NFNkyCyQXzdZNRx
jRiqJ0lLx4QEig7io2D/qwcfYTA0NTuv4/e/w0bBBJInl9yJylCOYOg77aWwfIpSWsklfnYPpf10
239fF4qogeH7mx7rSWKlWGpNEuy0cmG7EaUq3/F0CVNFNg+0NxuHKRyOsWUNBTrXEiRFJukIglEe
x1qw6XloOU+y7kJdhLjtNfDacfbwr9s2iqkX09B8GgnPhx/yaIDizkUlFlHA5+nUtcokqQilNnmL
Fhrf5pK3vdGNY+sIJfIUmLXsKO6OyGTJURX5DO2zWqjsthGJRMzpN7aqhfzjPbr9VocZEtIKXfve
8AM36jqcbOM3br9s2cC2JVaebdJHwJD+j7dOdpl4uOqKK3leV8JWdrI7CFl+b/2wJ4pF7whGeg9u
DBwodRMSkA/1ZiOc2M5G7tcg+FBIeGltaQRPOIcDQ/xCeyui4C6/zlSDCdVG21CvHnDpgFHi1omX
j1u43mG4+Zhc8RlNIqFc0SdH4/IeqY/zyaZ4fa4oN8F6dVANk4Y25ETvrKw/aa0sbUWCO6urNZ3d
m8KES3jg21moR9aEBAgDxCWd8IiZ1WVOjVS5TvbHLpYziXJgjDVCgUZUgiaH2hdhLY9+nBJzMUtZ
P1pRafm02DoPJEruP/rYMH8LHr/y893RCzIy8ChRPmSQgUhiYbAHTHuTVGb75JSwed//zM8rFA6I
aO08KMgUewmzP4cg2T9fDFALah0Jg+PzDDT1t7wkHToVmTYZWH5+1i7aKMpUQHSnLbQ7KCXpgfGx
DdSiM2L1UknhTtGMH/mFq03Jp5bt4LeC1z3KchXh1tSF6MAMWav38Ej0mXdAGh8gBJhSWag0zEHR
/MFp2jxpIQgQhu2vrTajZ5YiMSwb47imkWGT9jt/Af/GF7L723uuU3fVvxZtvuDa/6BkX6Xyh/K0
Ty1MxN8ebOk9AoGGKLrh1LkeSO+r3/KKEoAUHbCqPFhvkdmADUU4HTPs9fr7L+37pKc9nPsYtLHq
RTPaXIn3TQZzr5MVqkoEEDC6BQ1oXeYKdcTIYlgJ8b7yZ8rXSTUHMAx6SNucf2RNDK857YW3iDoH
79KEuRpvkfquc6yhUeeMAbw0E7TtC3n+UrO+b4HngEuEpsasocSSTdzYRPs020uIAZjznL7boWRv
iaNpNSYXLvDSzwTsy1iY9OXkvXq2e/Fg5r6m4ECsf8ZqQ6NeiiicW57djoKo9AUuUgV+pxjuBZkt
kw3vD/L4ReVkHtxVW45jxhrm73zk+oZ/gt3EHtTBFfJ5WlBmO67ljSUbBh2aKXOnY7o+QM+OuB6L
5DfsfYLl3kF9vSvSXUdVkSlpa7MjlLptpsJf7DaS/4Ygq9hgr6eEZlDMEH9PbAnFAh3d6ics1S8F
q5B2n9fyTleh0/M48cv6wdlSMzjkeJK/h17slrhpdmpkNYasYTHkaf663CJABb9fQ6E3tjWFJfCe
zMmwmnC1MIgE/oLecRzJLyPAWNdVQ1QD2WhmCNdIOy43AcQF3g5kom8/oDJ8W8ieOvv1wmbEi7Lz
h85KhBzE2quFBtKPgoIPUD8qDk588Q/sLYsVAztSOSzMMG9u8ywePJpayTaLG3D96Y9ImuqiHBrv
3v4piU7G6Nx2zq5WagRJ4ZBXZoV+d3dZpPl/OwHuH3dqI3GHGz84pEs+8ENNB018tNFuwi7MjILu
+fmS+xsXF0xmXasz++m0y6BflOxEQ6Pl0HuoeBQU2Yn0xTIeVsTDkblj9Z7+dZIgElB6XEovcc6H
H2fSEmuvzIHtAyDBD2/Sn68fZrA0ttthymYfqqPpAX8XLFaFB+iaEF/RgSgRVTxqQNbw3f1OquB0
/dv0gzFlU6uMrBElwBWTmtpdnkGMTfzHsa2bFdr8fVx2+YYi+BpafQOKh06IMSxyH97VlOWN0W77
lL00ADkWHzIYHyFgE5+wOOHjfmqoQfSANTqr3xQeJRSLeNjxTOByOrOI+hwZiISrOYSdWaAuQM9Z
3yzjl3y2o+OBBDoTkabXRKmr9IHyIiTphEPgDzySwVD3/nrs/nMcnwhs/S1Q+MQpkDH0PTakS/Eo
hHygesjyoNoSJJOnrKI0lqx+3VkC2NSiBEGiG6l3aTHhyPX9lL6gC06dy5t7RuXKiRZgr2eZLe3Z
6N/DehDKOezF/MkYnRWZooojwWWVS/pCIa0s87obdiB8ul0Ky355UbvBoVZ85921OZluX5z7mgXF
FrTioRscHTZvIcidEOQIHIyMHO1n7+07M0q98hTmcU38YOsXoqt11jfNXq8vluuCLsDJpiyFYULl
AYIjQFCCf3UKOmFRuHR+iQLllhC+Pkdvaae0ML+nYfc/LPupkvgIjeXfztHbJsheivjv5sqYH4Yv
E9msSe/RlZREdFhOh3xyEZX9zVNg0j8jVMIQfqgCLkV4yxFPeWzPFYGMgYLE33AfL4ErXRaXAGd3
npr9fZY0r/6a6mtbO5bmwHSWSvrGc7KQMSlpt2pwZVMakkSiXvwcvK7zTFUosXIp7lp9TVUieK+b
pxue10n+4BdhdERwok6C2Cr2X1e6nibhE3AnBJO38NWqp+B3uA8f8yQAkdFgd3KQ9Xkw3YUJaOo4
Yjyw2b39F5MXEYGMxPTX4qhPwKlH3BixTVt7gekPw+whWff/0kqhzdIMsBCM7zr+moZddBoip5n9
u5DyVuBavh2TmL88lidxzyTiV8UFiJA82z24SpA7MBCXR5xhAzsxGQ1QLoZqAMF8j7p6mgsg+EWF
x+A6cIjTWr7DO5fXn8crAybppzn2Pl1KXpT+EChtxOIONCoJfNb+j90x5vzxuApSOM4iU4sWxx9q
1gfJX5iAZBHrExjENlSl0RgAkKplqyTazsE+0gg98geO7v9ZA2H7a2dbna3chpldKdNkgW1yoZlU
/o8Qvw2UN+xlwOshyMO2cR37gMP9OEghe7xzEvv5msd83D9K5IY3ErcHtnzLVZjm4/yeK5D9Pfa4
hWlcNY2YeieVgMzTCQNwWHRtLK3xQKrR1PMi7Sq87BFd4iR7RdtXE8MW6gY8az3kmQVw7zPGSa88
eKRw/hlgB42ssJKQde9eaKesWtFdNg5IZTY/u4xPIAlkh7edP8gsLFHiJQHDXqrRMXWhQsK6g6i4
Ka2dXXhJzmemvX/I2rg1EcdfZEh/RTkU3KLZ7lwPrRf8leLLfrvglc92A55QSXN37oq/tXd57Xx7
83mDiWcg2Jk8S7u3V7Aa5AgdeV3mzxJ1BqDpKe6cIiJ03mdUHl//o0oI2cr1LK0eF+H+1XA6HBOh
tmMDBubo8hd6et6ZkX5hHxnTA1kjS9/pKxlL+paXJHaIcO9Pfj9Fm67s0AbIGCLfeWRElxarz/EO
bUXRdqpt9Yh+MUPvf+F36T1CENA9BszyPSEZ84fNcIVqlys5o2aSgC8zCrBz3BD+NrKnSaLnC/vs
+ivauw0T3+HjkQDVn58M7JIudqy8cns0Ss3SLvt+o88pkyrKRRRUJd9Bj1U8Knv9nZ0I5+bj2kNp
fpEwdwwYKyLpgzp6iTaqjEXFgscKHbvXSNoTjW9dmVeIrUjTaMwakyg0R11ON/1/oLI7DKPRatOL
iUGtcbSWHXvTVA09y++jQaS+MragvUfTohxCzOfvwo734DVdU3eQILBmNVicqamIm/BggEUY+C0J
Lwx5GYSuw2VWUFuhEbHfgxaVUc01qprC25WG1mM0mTedXy7jV8A9kGsl68zqPg602SwaxPKh0Isn
o9awkhC0o4iEZBq6n23SwCx7KBaiaf59buK2fCVFoHy4ovB+xwIyJV6WEIdzMKBfvSOFGkePBY6F
Wkk/vHBIfftPf0v4Jm09GKz/HZojFZvdWNKzynltA20GuNsW2ZDMrpXr3brWT6w7H8zFg7LChQXc
okH+k64ziT0VWdP6U5mJowDlSbiy90L9+ztcE19mu2k++XVUMalCy0QpytY3W9eRFcznpc5VTi6S
ppheGMQ4yVICD1ioJTUACk8Tkp8mkBmKJU67NZ19mH0S0xS6PRNS3pbISECOYeaQd3DC2lrLLZKX
91Gv4y1K6dmkiI/zraHG/faoQbafVgd+F1NaZVSJ7+3mHpADl8RGcUn/SC0JnlbxCJof6WW63ffX
LBNz8iX+ETIu3QSp/MskhBm4JpOHgJFwAR0+EXcyRkDXlPX7VLuPxqAtYXvHQ7gmAGu3vEEMO5Cr
k+5UOK8MEFT0L1u36y3IW9jafS4FdSkCOrE7jxOYbf2H55LjQM6PuENHNgI/o66JJcDcFfiC2yCA
qAu63Y9KPnhq0q0bEP1gf7he0jUyaN0x0reyi9k1iFufZyAwM3m0rG1kPT9m+mB9Vgbcrss7jwUN
xbjYJu1TkXhLrmKoIf5Q5c4p4lbzDIlPZaeEy3ttN+Qw/6KsnKeRwydGLW2GHfhV7laNOkS5tDAG
wlzsfakFF1jH2tNGY6x82cJOMWc/bdiopVmCFHBYuveJ+YMFzai08Uj3Z7gaYRlIPLOJoT63AE54
RPHEVgqgY3BaYhSbyvOdFIb7uugv5pEQjL02TVCITqaeP3b65520IEe1z96cWonIcc0XKECdLh1D
tN/V6Fy6YtsPXI9eC1QyK8RKJWBrgfYbOunfkBDDE3LmwaSz1p8kzC993gqIWJa36p2Jw7qM/aCi
EsYrhzU6eLO0JUt93QqR9OKOvyseWbqaLjaJMvANI03YRUrSTo1CRS5darFAD/QfcAGmmeaCQbr8
nrD/fy3XypsU+1/XORdr3Ay9ZgHJfqtROz6JCzaOxDzpicpi+UceIkSuh5XNmT0M+vZa63T40mvc
dYx24xgQ09mT1M10iWuoY3CWTZsn2KO96z1WMarq99MpLjq+VBvULH40zNBdNAqDMKOVC8MEqHlD
IEHEr95waKb98/JstJ8umsPEa6a+mr29PZ2dG7AaZNdtiiVIE5+n6MffoLNtbG8m+nktJOpaCMcn
L8c9ZGDdFu2S54TxPpRSPK8e3kPa7LzBbUf6A7P9fia2EZxuY4/VfJJxxlKboyjmfvfdx0Q2Ejsb
1TYgnY8pLZv3Iu29zhAOlfQ0YXGnAiZYKjptkwfA8o3Kwr8svSme0AWwencTHRioiCrdytdnblmo
VjaYhMeC6IKm8YBCZ8fQE6johzHAsAfMo1Ve+FNR6YLroqeyVW26ZB5OYt9Qr0Qq8AAAiMyFxhEV
0gPcrxxVzf1g4vatu2Pod1Mz5/VZmSdfirKefqujiMukKh1GXPK8JT/O8MPqwDbFXUAd129ULoXL
M43V8NF4v0VemkEcJv+NFzMs7E6zs6m1T1cfmTFiOR+Wyw9hXExxEITyZlmtopnnAMW9FVIA+MnU
mNGCMqZzSjnz8NLQj7qqUpOCECHZvp7+3tESYU+n3LPG8qmUaeJEQzfYc15Arw5FP3Jm80mDGc4J
aS9UYC0/X98Kvwlve9g4JiBIDM6oOEIikg6zhnO4g5Yv/bBGyYamz7HR6VUgMZ9Q8Id1VIr9zT70
AiEW/ppnjdbt0R1CLn84naH5r/atmaImyejtxt2DDCChgk+stoSpTtbLc9deD9lZz5nWPf/pKvTf
q3uAHX3cjH1qiu0PlOGfB/+gsBNN7beyq+6i+q9M4nnDsOECskityukTQIQXTQMcxohUDfAIAYH5
06e8lnG1umnioc04NivT440M9Dp5vUPHgjlfuYMfQL9nIHsmjNbX0CXre7fIH2ptvDYRzdALnPGI
9HWin1ENPk9jYma2SlpinyIsrgUK/Soo+/y1LXE2vWXUkDsnKJYbJgXKI5jsYGGGxqId180UupmT
tP9Fl0E+fSzz9PeTBTvYKK8lMrQ6bx1/wPxc+y+KPWO7bEGpqgXm0wcsq83EfUP75OQt5nz4db+U
w+yypoz7nNtnIib6EmIBCngWWaRnZYz7Dkj/TThDUxR59QDxlKKzrtwKsU4t8GxKROC9J4iYHMyN
q8mCYsDMY1ommDNo7Vp/bdxryOaJT3hBnj+JxPFqyziN1QM8s76xFcW9La7UQkZIoJmBqMJ+PZAQ
ve8VLSuWilnC5Gj9QStpwgSgwDEMvjz//zSF8NqtW/8QyCsAJnNXEKa3ISNybhEQAhOZGnAhSkwx
kGZzDaLhezFYyMi/1UnSYntbgAyGCt/6q9WGvsXKUq5JGRhm7o0A6b529hQprf3YAO2OJJMuuQ2J
FWFhuMs0Yg9UwbSs1m3SL4W5cdzLQUL5TyPwbZS619xBN3a20TsfZtHleeOBUq/5OXeQsLgjvGSG
/UgcIxzD4ucJDAyLajia3nacBPHUpuNvOPjW/TWZVeEOdaf30MguKv7xkuYYjneZCSeMEdDHRO6w
r7OBao9RL0SwGenZikmeDy8iXX1YroP1Kqug/QPAARgwsYpDJz085g+V2nXWQEDuWglnZ9zW/3oG
emKpucbU7sCaP7NT8T8ugv1Hz3r1T6h2uoEBcXVv2jze8bLHo5ieelbB6abjeIJpcb4cB4z6BQJK
KtkG2UoB3qBVC9fT8ik695FkQtcmVvb2Dq4FG44Y9HieDeuo0K8Lde5IhaL2klQ8LR70ad4PKCIC
cU2FrdL0/bnbVIPv+y7n6nYgdfP4ghd66gU+tmraLT/SjW+s3q/3W0hRBa7niKqM0lEk7voP0RJr
GgUCdbpIwdRqyp542T+VTdvMsFxpGwqBcJBngboUg0MS3s0hz2qaIQ47/KSongMX4QUaoKbbxaPQ
/7Jjto4G6b/TjMRKH8nq4URl1lmfXGu88nkXIDuM0WUS2OPEKvQRkCBFKBb8XTjaMpRYyirtWPGi
vN9A0gRz/nVLXsNxE8wqpnMgTg7CnW6loqUdnkEZO001R54jY0TOayQeudmyq0tHJvD+mtOIGmSv
zkMdDlp18ZZm8wsqS7R5fxyeL9EseFb4jcnD4ZHTGZaOm4VXjg2V3U+B6uSjhXzZrN12BMqyZczt
rNQ4MedeWAklojUviWUHhtj/Uq6xE9f735LkHgZca96YjazhZQdPpIUGgMyaqiPXxdlVpv4WFcUk
3DEbgXhdqOJOg3Uyh9XFazQu9XppGU9FvtTcfVIzzv0HnhIyMAnO64RGAsqEddlSMMYAm5OLQhYQ
6nI7QxEGWL/SkSihviWEaNV4PmnDypQJ6YxPEDY+aTEPYsqNTOXe7i23GJK7jnNvFRyMwoqe3BnA
nfgb0ParaxBKathycogdVNJizbswKU9akdHRNZGRICMZHj+3mK1rH7AM/RLjvYC4oaSr9E6/eVtJ
HiBhIkuhNrxCTGIoCijWv7BdLvGCct2PMZc3EL7gHZxic5kC0XyC04Pj93tDb7/6HQvwDGzbZzOT
hgJR1q6hegbE7kztAN2YiBS/ru0WiPjuhMaSbAF6Sa6gMkWbT64MxNaz3tyCajDQsqEF4Ec0n1SQ
dTzvx78P1LSwBntMYC0vp8Gcn43rURWgjjYrdO2Cv7Spmu2NQoSn7fQheKLV70HV40onIt1wUK/3
52SS66K4iPaZtQNHGE3b5jQHQeRkbtskekaHTXjDxz1ScFVn5CmgXcNNXMv/vuf8fdYHz9rdbO+y
8ZexlJK73JpKG7sSo4wPk3p3vZp/KHx6oQb5449Me7fFstp/NMCD+0dAl16DnasaaIRChXn9HeU2
8O/aocnPVLAb5mT7wnIBavbn7TfObw/erPsBh9uuC8Bn8mt3WOjnywK2VqKhB0pHeYXH0BOP5BeW
qmBL4gPAFrLxRyo5VuYotjz05obudK2fB6YR5073yQvxbyeoRdALjk7FWHrXpkMrz4nKPTeN+o+o
hqg71Cgmcy1izyO3p5SgqFcfRrqf/aZmXArzJdC9O4rrKlkqLBxV/uHspRGrxRRxk8qenySj49v3
3sqlW1g8bWuAcdk6UxNQu8i5DLoEmXcwr4GoNG+5MSgqu1D3ru3fLGSGBNGEWExCyz2iBxf3wRxM
opKPyjF/guqFjJDj+7kD6IWVrdun37fZ7j82oqFdatn2KnFVxsqP+XHYQaaOGuRdcrBZPQ+hdRhE
Mej6XJIsBo2URD7z1IjALoM3h11vKx/JMbZUI08/kbxYrvzvsoXfPsBlc0XODms0Na0EmwHCozMh
f0ErVGL4C7Wi0YIeH7KuV2lu7xVXMG3lV+5X5Fk55eb1ha460jxDDz9al0au1mtwL2A1SkIhfLaA
9w4LbJcmkcnHE0Co7pw6lHR9wdmDhKTHs20dIcUamaLVHo+5hJEHLflUYX1+L6B1TuBHEvRr5brU
MtAPb74OVE3XYE1bjU2Szjb4j/Iu9tlNTiPabJSpK4Fqnj9qzisQK1Gn7y87Q+0tEYAfHxRB6K8U
PdnaiApWBWV1m1fN7Tnhw5yVkCz0owjqymA/9hqnYkq9vJjL5PUsGCfPitNe+xuFkm9YWZcV0hvT
PrRTXlCM11o2plJ4Bev68OFcCmx+WqBs64JYwPruGWwcFv/ndDcVCu2blaf5hdwkxdtNNekR3e3Z
5aDC14794wCXggo623DuHwZWBZzWtlBDXf6RI1yDhG7TwfUip4seRnnUXaUFXDYfl1o205jSkQhw
AjdFcRpVJzeEkKXbAf9gwuPEa921eRZVY4+iDJF53MIiSuCcTs3va2XarQAui7O4qEVyKFiIEvM2
R/N3wF+oC4e3MwTkwgAc9O8PVibbX6wSG+qDhqPrPAJ3w9XzoomqJpg8FpEKjkI/djqUJkgDXnY0
eddF45Q4fqDnb8ZK335MnBSC8BN1S7jr5RVnuelJLG4aTJ0cKUmkyXjOwIP6lTPESEt2mjw37f/g
agUVW5DjwMSqjcoV+eFw0fX9cskoeqHSOWNolBw1t8nTegHty4e2QO04AC5h/4pM83GOoJN6JWO3
q7QuoBGOl1hEhLV2YUDmjl7sQYA5SpglTIdzc3Fjv/qKvH1pH2XfdBiqPh4QmPEe6AVPyg2mGJ6J
7c7mfSTr1z6aAQPWGbAN/fmwWQIGvB0pekqL6aCrFKJtCKCfrcfmKpKXCK/ZirCafoQ1GYu771zX
0OQxva8hQ8dDn3jtgzATlSdVZAqOuS+iY3ebPXwpxpEU3kUMDP9TAj1oA7TGdiThNsvyGshrAtmq
IU5v++QqU6eSgQa7l12hRYLpyulf7PNMuP/r7oZl8zptBa5OcdBqLuBswBLMeBTF70QfgbK49Gw5
3RyIfw+2hdeHMKfGNBo63nAR0T+gppkBNZAf+Dy9TqGQ65GTAXwN1d1jwNJVkq7FfAUxMeyGu29Q
gNjs0XIKDnJ1LNEl9UmptN7ae8QocOqY5BPZ0+nv1DglkGZmr6DjqCrrsqws+U/LtllwSLqf27Ac
z2ng1kQOSE/MjBwFZDlNaOwJq97dWJ5nYP838An7LsXq24nejFST7AuaSLxHi2aBxKgDpPfXzqrl
0YXicPSXyYYwHMjzcRnUMyp4iRbZefxCAYqtbkjvr8h/FZO9xDJjhVAf+oJYPxLQ/+xQ36t9inap
WcKqMtqZVFxecV9biYoHo5iKeoYn4l9LLQ57L7eKMI8egalqR1+gY8O3Fgf2fqVFKO2LmFyBuOr7
eCwOsVkIZaq3K1cAW2/BotvCXH6tsedrR3RfZ9kVp5JHph0bAW0I0udcrsSyV4HPZ5ysAbJqSzET
CrKsJj5DEeXJ5ikab+KNyW6Z9AF87O0/yQhkzcYa+YYQLTtiJsGqnqo7BfKN+mINF3Lh52Su9VSG
zEjRY4hXwOhJp1zuAAaoqNNlYs1KjauY4wY7g85rFSMAz+gtxp50Lk7frb+2FAc+gT26ZhgTY9D2
1aSwGm3t8UiFlzZRDUmPTDOx65QbUfsnIoApUluUbgMB8FWGprKLmI5i9G77xmuaVT4ht2qEZnxY
fhygSFiGZRlstIwJGtP7tB1r5TnBToOw2Ye+OkT/NRG+LdKFF/i+bor5N8NLSLukqjwQvNf+J8eI
HywSKazWnLV9xCxid1UsAjwn/tNJTYsOCUC8wQ1+sZF5GnOax3cOY/U9q8XiWjrCWgW1rUdaYJJX
3/nNfFCe9Umxf/7h0gfqsF/MVpNHBr5gQVPhwuKOs5Guzwpncl09s4MXPyIpi551vw3AQDI/Laxd
+YChNYk4GWu3NY8qWQtoIplCvcgGpDGEYL14lOEUoZ01on0D2jSsHQmzkgfIvarzeOlxiDVM5KlS
KfdMhwY82OfFDvLKQSz0yBbeSk0Vmvnza+rvRjjQdceJM1Gm9MtF5emJHlLYadL6XmjrBrndAKBT
94kXl7oBvGfQyx7hS0L5HyXrFcF3oEKoW6nEV0C6oikBrTKk3LiBUk15YancBMcKgKDM/8wmkmuP
dCdpFb7vkjDElnd2mzokVkkHXCXnSqw8BMRAsQ75OSxiGxv8THvY4gqOO2yzF/xZhGAj9hHYhgSf
pyMTWPL9DNsNc3L+HjqqRFRfaP/Cx6JC9Zz+poHgmvjmSC5isSAwC//igj9/DmdcnZoqGxqwfWAT
IiY2Q3sB//3T6YtConoSFqJeS/m4RPSAZKwZWlr6EqrBoZg3ZTzgiio8yzg7QJE6bkcs31CP0aa2
OPl4MzXx9n1B8RHhF0eEnlD/B/+6TI4w/tbe0NE6AOqTzi77sGqdXqHq89rShr8jrnB30wOBNxgq
7v2xSArLGk78BopT3SzzeAjw49wTWKvjCzCP1qSNaIynfEOZcFOZ2w7ypb3v5HBvQQ3fR/HEjvdY
qEDfdjSbvMrchxdnkQ5xFW+vaDbB4qyeWQL1iMQeb0U23J9AyyUaV2AgEilG/HRRGvRKdjj4Exk7
zUGcgeZGkJ11NyxwgbybNiy3ynlzKncIn+sXqkmhHtIxH+ny7x+ht2By0hBUCz3SNtm2Vs3Nbrsn
dKy0xyUbP/r+KNhvMhkne4oHHeSBQuBFB9+LEUlOV8Tpwq7XX0059SM/JRl5zNYQe8WcO0LLu7DZ
fILl+ZBGSvKwIn3DrxuZvuffKGrW4VMJ9jPoVy1UXDtasbsIuOeWw4wzjKQG/WeY6tHebnLfWN+D
QYEgBg96Mdfho4vVfhlQJsLQlfcHRAqYNNgrOyIZNoxvg4ZvlH7xRQeabwvPi0YNjY8zc2O8ROJZ
2aI7f0i8yQoHuRj36JWIDw1WolIp8dPg1yG1qO1mjBQjEaVhz8clfAZDYfKARyOt1Sr5DueW7MBJ
+HaaZKaszIaSJ+ngs3xJs177T03BaDjEv48GY5ZmpLLm+Y0KnWEzCfyjokat0JmfRA+URYWPtg73
M/0IAmVgCV/dc0znRhtPKtnq+JtIxzdC8lTlnFOnkwCm4mVKpxVz7FnhwOrmahZxDYmS8fX0jZS1
cs4vYMXhPqlePikoA366XqbYg2l/W2DbmILVlgS7T9+OywkR3lIHEEAUOtAy8J5bngl2KWVLJFVw
GBOOzCGQ3gG++3aBhtelAD2d4HgcC5c+H7YNr4sKzx+17BaSx1KW5GR+mjVXOJ8vAFpB32kvDGXA
WHarWTl5w4GS+byX/6N1povHkdhwl5zeGeM1vJhSIxLYoUyt++2O3Ok76vUu9KRcii4JBM5U+67E
PNFmA/qrDTq42cDKnRgP8Na3/zWrZZfLi1IO2j6zw+tV1qswrHi404t+QQFEcP/zSN/D+2D1mm9L
0sBs8ah4dvxAA6Bk79fq/6DqzkV91y1f9v5WnyzyFG482YYJbRHXt4ce6BL6p3LM0YEkqgo7Zuwr
kUhZ6Xb/WguCJtxsbGHnIEGIWhWKWML0qdmr1yyzd3qcV/WOd67ZgvpSxLKLJAH3KD7GWcwLiqfl
jQWjkkYCLTJrdDPQMWxAxrKTSqJ5yowHmPBgQJhMyGWFEa2yVHm8oZmBD6wRQA0c7GqeNCRVRtWm
6STUhnIuYiKeL+jUia5wNcuQ+g3BhsmoIc5sXl58MgAz6yeiHw8zHpjpFtWdtZoRGya3GVxCkCze
q1VHUAvdBzKFw2k55+xvnCwXuY5pyP0jCNpqF08hUibqBj4VD3U5/D540CyhuJpHoXyCgc9TC+TH
fzi+JHuyrw2N4C5U3H6ebG4qwO0BOyP8yY5bjJCfakecSno+lmnjmUzuOi4UPHyeZYg3ub4XliyM
bIOoyzYUVwPq1OJ39HYZsjgGLJvEo/2dC5Kv/iIkEhpRyHvs3qg5YAATycxDJROj6i2sf6dLHEeA
omddsoTI9fvO6H069d2Q3WqAU0rCiAGJsGUXq+wIk8KxW4+y4pi8BVutncXp3/3h/ryFh7FTPLYH
JT5YNne5nPY/cnWCeK0O8IVQ0RmkHDdCdX+bqMXMD5/U7NJKcCP5n/w7WTweI9oqKwEHIa0Gu5QA
fjnsvG0bmPgA4m/5gwr/ZoCQMYrpH/YchiH/g3lF4HS1UuZPkw9PTHPGpkt9MGV7uzy/K7ftixBU
bAuQrght6oP/dZfDE+0TorO1uQ/QVtrUkWQ/iRuM7TACuRyHjRryaFCsV1xeDMQhIJcAKWwr+gYd
8wBIT4Bk69CL5UgtoBa10ZdEzkpx52G+jdYlVwWs/2rrweR3B4ZohXjvRNstWV9x/exxNWJzxmLo
YM93cKCtPgljUZezGIp5aKkMxiOzGAqgIGMKFtCPJPl74j9ockXTw2EzWB/YZrGdxmPpdDw/jRst
feb3bCMGEJaIIxQwkSIt5BkSDkZkUtno5Ta9QS4E/o41BwWXSFu+XRQ70EeC8xU9RYggljLKeCi+
xXpniSt+MGmMw4VKaLN+/R3wm5If30iltiBAY5I9bEansblN19/oO5ojv7PTBgYZdqwVFUmzDMsy
HeB5fRd1UlGbiGfFBI+TUeGynpEOh7alV+pR14PezW0PIqjk/b05/PR80w2Ylao5bQgT6EFYtPTH
USjjm7O5b8GyjYA6fuzZesCdyTTwrLT7LHycrZucJjQ1roMHPLQZ6tmSl6l/6hHUA5ewva2y7rfe
ZPDjUf7r3YWjSlrmHj7ZTP+O2yaq4xlaPANvJd/CbfWbaxgDAopSa9QFIH5wdF8kitCNIQxcRbah
QJsCff8rk5Bz2s93ZJjWJNeXD+ScMsIgRTH7CCFGi1QiboYTvgovpzlkMlKJSZ41duu4rn3blYjQ
IWvd1nFDZrCml+0C1tku14Mju6Z7YUB8/LhCe263PCAlEIYezfwD1UCbFL8+Dw74bCn2tWAX76sj
LRWWfAj4RetP+BhgUoBzqG+svDP1aIUg4Uw2SPt6sZH8RIKaNhWmWyOaUNWEt/wKM9RaMcxqkTCE
i8513pIn+SKF3/kWo0CDwfOHtezug8bBggoW6Nf7A2qv/wEZmzYlsiqJgjy7vFA84y8MA9zSby7h
y3aaCZxSBNWZLZPyOaBwvdX7FULvaY1UI9Xqojov+XKH6oXjeqOl21ScweQ8CJHoX9jgbPWrO60x
lfjR/ajLiAxVh9ZuLdbl4uzjOOJKStBrmQYtHXoI+OEQHIyQ/77gSay/X4EqYTC8D8hBhYs+wPjc
rWcxMVxvrz7/yZZfjAsLiISnPAf103QUhw3B912Jv9ODuhMJmdw5rt3k0VDrzgAmEjhJzCQ55UrY
5e3sz1Vlno+I/lTHL6SgMG9uKByR3oYJSzFCzDCHXPtjPsl1wlt1mgQMXjbfqPuGyRnvsb51mREA
DYHhKnRc6fBx9r8pCWkzgxV3XEvIUOMstqp1a1x3ylmF2tiBI6bG1pbrlanawqwnnaNErXlU5oez
HMPHOmj8wjwbYbj+5Tem27U6Ejp/LUVtu32F35LqFQqqX/kKwzrxIAjkeoMZHbnNQYOZVtkmhhNu
h3YWNF0PfO29EhOrFMldza+DqsT02eTedxe4ULepZRUg7rikddVmhM82S4Ef86DPC+vjaGGcV2F4
D9uIY0XrPRETTymh8xJWo1bgJb8KGBXZg/fYf+RGYieyg6/5LMurbat6hDZy4hsqmxTnP5H7yiLG
KSd2yUBmuSTn/Pas5eMsYFcAmKjKmdcciFe97Li9jiLgdDhuQSpV1cK82mrZnb1/UgacusSGUgd9
yKoZMtxjIlrYNbMXVTBU6jsnB/crQSbNTPDmwDUMjA/WWAk62c2ndIbufMC84iCsTgu86l+LkBIk
gXzDiy0Do43+xsHJIk9+WxaMbI5IKipRGNI7oa7whPYiSDcRL9hKl1gJ0550MZfW/eeSu6zbb8V2
7Bz42wOKRAZ8KgD2luic2abwg3rtrzs8P9FKBIG1UUkOEIhH7KvzXHhOQzFg4ZbuDNkmZ/7yZHDy
QxuH1JsMyujPtA7DdRERvXdgUoXdelV2RmopaHdcpqBwhW5/wFJiZoKYJ6KvXehYOwzNDH2MbEhN
nHh4XO07dLT4NXN3jbLgv4k2jjZS1nY+bLQSYtX9yblvgasr5Vq7izKC5dzxWsPYnikDhr1TDXD6
2pOulHHfLSzk4ia13p3pCYmWqUd+PTpMtkDYMiuv4+3Xs1u9Vt9IOBG2/DEKptEWOknexlp6Dkdy
BD98M/0y8deX9Yyu/12RGw7X3JwOHsToaNfSdvDkx8MynGynUqc//LoZBEiapR2y/u8bGsO/iueU
8GH463RM/M35/wbGuPIeOSJQR0d9LPTeK/sSIlj6mq5BY7fnIQ0m70Mfrmnc2qJjw/4fJg3gQm8w
7WBkq3BaxiariN3wQNYpjm5pka4n4cDLlk9WCKHLYmtNijPDmJO2ygrHoPxStmYR/EiV43yd2QYC
Lo8U39sDpmvYPYUeyWJ6kFZ1tKStGz3waI2NMpKYUK4pDNC50cHV2ibR4aQVGQl8Slu/SWbw2eeH
pJKRnd5sqhSN09Mc1WLPwa0QfGG/YUioivAAYuzQPyTDGu1A8lMvpmVPu5KHRVxjmzxw12eOn7Je
QquuCo8gcZhxoyySi6CnTgZXVNqTEyKfNxEWVHZr7XG5ATcKtYmXgP7mHTbBJzqcEov8zWPOjQMh
LuIPy4XxyeKQEq0SP1J7pSdXeQnydS87jAFj+z7b0j9GEMDHkZf6bco2fzqMQ8OGIqsiwifDUfmM
p1MQkvumzSdKWIxJeWKnjAVipApVSzaUWVb0mOmVVDIZ4RriJzZUXBNQHSUzdWDxbs+SfCS7Q28o
8roglU8mmIQLNoDT5zO1KQScb83S9Un3dizE7SikYmDsqORvs/kavb6yVeVJQyxIseesk2CUDx4A
C0wXcc1xTxIxxvWvEnlxlxKJ3i+T2yy+upVv4bB8KSvllnlX75VFuYr4fwgmpMKaxAHauCxg9+3W
svCd2Ty/CvtIAjy2hxL6txu3gQcqxfI9Xdd8a4xmxUoUdn2DwdWQjsRM72NHPNZGcc3+FdjRmUke
GKrqe7p7MDgD7PaHdG48SUJlIqgKv8Vd4oEw/CQQDEdYPbXuGrew8uxSqqO8TTYBwpPDmbwhoja/
aIY+i7KaE8G8GMxmhhgksiJRRbBx8LC2bmcr7AlRvjQPtngCNoVARulGO5f0HwDBQOjb7+l5aANM
ahBBZ/10KhXb0/ct4nKC1MBeNWfmoqMNRqCtz//ICayGcArO4MY/234bFG1nhDXu68aq9aWgQyFv
NK1tdFIxwfIV0CVaLC76mipda2T1iLtL95ANkzMAi6vP4PGKj5W/z/KY5vjrlEtBQc+7hZYT042+
SGtMsDlstAqzQjIRd7FNUUe4vNspb7y4igRt70KONSIohiqnr6SkFK5gjSGWAZYXN5eoieTFJdh+
J5MF/HKJBP6iQNRXa6nlDlRTPny82/zeywcYptb+bWegQ00PSilxzZe5KxNaU+Mvtc3GV+3ogw1R
WYcwmEak93x8kpS/d1V4DQZ1GeI7gyljvoRqL02bVAW3axq9aPlGYtZGnG9orA8tHu954s90F3Ad
ycSXDueXeZNvVO3LjkQP0RT5pvbBGmwA6AG2pdj1u2J9kitLnVpNj7LHZBGicqxWcJzOyfT+/5wV
jIVhOUaDZqVnqc3MqhQnqfYV6H25rNJkZMb3mtJoyJXtQnyKpxR8XLe032sVe6FkxJaVlb1VA+Oa
UtrcqA9ZAApENzDev2r7be5xAm5VnpwKF2NG5Oa/sBIkTUzNl1UAPYnhufWK5H1F+EHNz7eQ7y7i
bp05p1HaxmieobauaHkqgxB9zi1mihm9K1SlAUo0+63FC0qxuZBav4C4VPjg68WnIU4tegpqWvZw
TXtEZe5kjOVIoZhkLmOG8+mXD0LXbRsfcbdLhmonfO9W+tStl6AQiIoAaThkRf9JbHy8eRcctpgh
sCMbsQ2eNd7ApS+RKiZ2ipW2Ql0oBbNKj1CzZKdpH42+6LNPQKxKya+v6I613X+6uNeB4BNr30oa
qaReGpIs4yPLz7UzQ3dSfYsQ7AXvK84xPqV11JMUri5nMbsyw/zf8mRWYKVSFdb6d+XQCr9gsCyH
TVcSccC/JznauJCMjSvPfYp6Nz6z63/4IvIRCXMmRWohWLE2iBXlStKhbrR0ypXZA3MQ0pLfurWY
g5wQqo1SAeVlIu1E/2mlXFUigSnzKkuwF4Y2pZ2wQXguAdjz4dtIfPmOYalHqkZcVnx4uqPGgitD
gi3MrGRGQjVYgrtgvK3wfKzMki27hG6hO+tor7huA+QnA6RGbj62dSCRPNbCbQ2Z+749vzOSni93
JK+/teqeYI3BSTJq5noNd1e5V9Dh2imrMEwskYT0KC5hjMQY/eUBzT8te2jPa0LxYj1m0ILi+js7
88SQukGUI6/Ba4E5n1iSGqnhA7eLDmDZpk68v9Gjm4mJWZNg5W63nG30B/5S+e23TMV/LERvSI9f
6+103oLbjGYD3OBAiFhSpO/eGxCVyoXXWEEohmW0Xw/3SiBLKH+yKQhBZpPMLGvqhxhVa44+Vojn
5L8ZsxlsqUQ8eZA+xSUlBLEnGHzLvwGg+3tFx+EcfgLP74e6BOm0ReYGfN//d0LQsXEjrw+KxKgS
CvztvTT2qftYBdHFsJz/LIFiqbUUHK4tW1UrVJnpICvt+wwjatUP61f0I8l8yxQMKfjjTC3gz8XT
LmPCz3NyXOKX0LaorRWzVApcQw/3Y3K2DsYW+Foup7wR1CJrx8IWUs+o7bG70ANe6mOo8sfOXkuU
Y+Pk3bgy1hvBddjswq+wk0U9E8DM/Sb3b7BdHcL6F+er2s7nV5yZazkm1LelA0poHuDmfaf875hE
NlwvaGZ6rNkSW5kgg5rjOqAVEVfbmYb8o176ZuFFQhvoeOijcaSHO/RWhgJBHQXwzXgzykt+XwN+
CsCcxrgf619yzuW8HtkLnNEzo3Ez1yhBH12Sqq3vQkMzd4M+9vuXKfGLZte4IIKNF5GgjJ9mX4t6
jWwdyidmvBDmoI1XA+9H+dJDbGhUD9uqgdw39DNywPGlk4NFFw0nGIzKgT8lNkvU4jdiDtNouaYM
W/iWpMGjqw/IFArJKtHn1hmgm7dg9qvms0XweVzCN1G8/uELqotJqtSFi1oFsBA/6BfbVZTao99y
8+dP3b5r3Y8o9UOhQFeEaKAg3H5Wjpo5QVIxzoAqB7dLxiQeFw7eH/JEKdE/Sf2rB3UVnV1zNOs0
pplq5e8xvdU7oe3hp/WKgq7x7WYpmAsun3a9srrrfrvWpTSBgcIRFILOj1MF+4tcVhz9a7bdAgzI
3gVce35BZz0/RF0eJoLzJ9Ito3hPKsBG57jSXc6kkJ+Td3DmQyEXNlTgAR4NY23UwnnmJlBXtapH
3tFm6ZBfBI4F3gQ0Slj5JaGPAIiiceY5HGYZN1hzTo8kEaVL/9FjYsaLjtuVAv4UlNFsAXNfxh3v
WOwpCQLtwCvD6O3UUkIXI/PkYK5rnPgDq+kcRP7EKfU2m3imOcEz3hWtZAl+YaTr6JEGwMKsy9OV
t7J3LZKwtf1vBpchGfwPgO9NnmVch3YLHif/FZw4MiLOWTH95jrQEVwePmeM2b43MtKdZ94aK6+t
NccV4TGIJ9vYXiGpu/FG7kdyTJtAkKvPIwNGYQ/hhYAOd3ctpW0p4bkk8RqXGqhlwTsfuc1su/F9
j7RO1tElN0h3Mgh/qQCVORBU1zY1EDpuePFWzfypZe5DWFxIOHgikaKMcVNhQt3qu8P5OZFCG2oJ
k77VZ18UuI0qA67270UmxHFJzQ18/DgA3/tE/abCDnQVSZw12gAu3W8uT4Ihf3dp6IqGJXQVCUtI
HnRDkzrdh8vhHu0S+z4S311QrTE0nwp/dMiEdXmv7ozMSBv1rzi5DR8XdSZ5vr5qsDnd5aQ20bDF
52kPt0cHZ51dFYwTY0s99QzGQBf2ErGK9Kev6xjlZwOc4IPNOExGSfPbi5v6d0VkJj4zAMbOjyGr
De4axH3uL129rAn9ESjhpDp+dEX8JBl4rBs0E5tFCPPSPCmN6FucpfXfNeaxDkNBxP5C9r96DDfv
JZG4X1Qyjx26CLpaqo8zbHUahR8+k8R9t92TrUa7NMzBHaPMJf5uM4HJyClCR88QjWTwmKxZL2QB
+ivVGWHxtY144NDUcyYKCkLgOyHRemUj1zWDv987gF2LDYhjVoLxmVO46cPMkdOX9ekdOwgdL2Nq
kT1drWOoXriCs868tKv6yZetu5gGrSDXnwjOXb1Lk3M0NK8oGe+EsmNPYvOuuGDvI2uV3WQE4dBb
350bk0C4LZC2zLfwM4OYck4v9SKmi4PWXGbVnZhwIEoQBkn2zH2L7fiuvURytBFpqih6BWsQosvO
wnaci89HcieDZmlDajQ80RRMOHYqRyqt0HfJTDk0y4eoav4D2wXMOz2niYbOl0iSdqRdasmM21yA
jdHfKW6BMZMHWJkQUROePoW3BcxFzqCY7/Kzch+oXtuiEJEub83UEFgOhPJzNI0+/az7R2Ngr1wd
JyhMs3oTOBK7eYESPnO3e0mUEgTY4U8xC5O+QiDMHDmqf11KZSqKlkoQ5nbxD40YH+F+rou+wCag
43EfXaJLfUcGY0KWTcc9x7/GvDHsh94Kj/keiwBerXOAv9I0vnlIGM1zoBM/pjTl4IfBqQ8m26ua
bsjjCJ+q+zRzMipMj7hGhXXioyyjh4ooWuGpW4YFelg3sCw/hI2CpK8fK5k7Or6OvCi9/yxXfLqf
6ilKC7ivHrLlM7DfdOBzmS1kkYRSdDSkhi7+mRAbxUG9kif6JCpYV0lBB9Gdg2l1tdkSPH9Yj3/k
9FQQdHwmvwzskSlyVtyXuydD9bkEBsdxUSlfVgcrYPkFNeXJ1MK8cE0SVjRvG8Cqi4gyyMIrgCPK
6yOBzuGkFkKtTtFOaYZfW9CS76P5/sH9Elrh3ZdIElJinhF7ZqwN8+AdRUe0Nx+XvCeHeacUdTXj
edQADLGwoKtB/ioJhDImyR1ekclzfC4PNT+m6nttXKIFnqKm3LLbbM3N57ct0NU3dMX02i0XDdXe
HRJFgivONv7CaI9V/fv9B/jwK8GZyiI1GgBUdtZeI6RJ6sd/Jr+aU6cno5TP2KSr3H6jfd7dT4QG
sn7xOBXU+FZawLbqmu0HOVScBeRiAatXTaNnTvm3KXm8onKhdLd0hA4Owj96g1G8TV57WMsLcqQJ
zMOniFKcXn5ImuHgm+BEHNWtbZaXyc/O8J9Rgq4dxrETL+N9hToD558xum7NRCcLA+mF7tLFifnW
BaruP5Fn1Y8gvtqY1zkKkYzlbhElIWAGP4vkkgHEFrXBGU6IPnUo3Ei0SaYVX5qMoc2JwPS1JGRY
KxgjS1OB9Iyt9+dvK3Y5d/bpGPctY9I3O6L21zSJpJ/uSwfZeNtojcqCbLwG+jHiy9Ua2og989n2
i/q6pc+IhaqjoUndnxAU+t/STE5e7isF/rHpMFRcQccsksXtttZDtGOE59GDKrKXP4ue/LZWgmAv
W7mhBhBDFR3VCIHeka8TPzD7XJAuzlwplIYtM3i6ppDdevSu34JqI/+KJUxxjCGXvVYSwiy08MFX
3wwIrqneFOE2JhVIVn2PqpycSBqaUWl09GLDRLQzKIsd5yS9qLu0ovI+qOA5F9nzLWYh6N/fXT42
i8HodphDHia6ODLHq/x6DnJszST79OfS0FZYEF72LAex15DhITn5ix94A0X696R0itvnsWFzCEpq
QXJLGY3sPuSCKlMAlVJ5N5NrapPiz8BfoLTMRD1EvoKiDxo34UTm+DfyXf4budmaTjAzCyB6Gk/c
k5YpZ5V01x4qdJbUzZ7NW6hVDuPMQmUKcUga0rN5La7beXzH9aQriINR99NsfOGpsLaKE2p809gs
0OtA/GyTgG10aFHGXrTcyKE1ukHZ1TUze/1Kti0IUN9QTLycRska/0uBx2hjadkeFTR4F9lCmj9l
FbENEQA9p6ikhK9/BakGWk4WwmS7bsHLcnKnF5crpw3H1/JlD8Qw9v/SvxOxHUJEcvJDsBpB7g4O
Fo35r8bN50LvpvGJtf36jKSNjD2gG7GfjHBe0UbNd8fSJozLxj5JFHS9mo7eOXA6I+8qEdQVlUoB
5iP1Ovzi28rkqeSlt/BbQdNoDYGmnC7WyeFDYFd4qzdL3h0RMdVVSZDQQYQUs/yiHExYRrfqoCL+
HMeUtz2HhQpK+WXO5fxtJErkKKdKJ3njIKrauCgxvUbsXiqojDZX/Xeb5HwBUbkO0gi4zaLB7pOV
EfDonqXvEkiuRpVXhlFXF4VP81rPo/I+L5IdHM9vc0wPeJGZpy9ypF7CkjQ5Nfpvk8TEIijC8+6J
oz3vsDOSHKEFrX060LGCbBu6MnTyPgkGf3U9BlRELEJzlWNfLdqcYgFFVCZeZOqKV/+HT64HU8Kl
OlOEB8fCDKlJXjH9vfA/IblOE2OW3CBWj7aTrUps2RBS1AS/CUADyrcQHI+vu1/YLZZAXfKjiOcm
QIGRUWNOuKPuaF7VbFCLtGV6lSWmMCWcSoef1hAhfJ3rCubRunMRpnnQYKUoY743a4UgvlC+JBIQ
NmlwTxwC/J1GUTWPqwQ8N61zFY61h5r1PCRXtfBFg2Ig5HUy3/KftaflKfQxf+F7wvtlk+xZ30Od
5IEWqvz37QvnjcBjwQvChmRMhvguIFjyjR+3QdhhfZyCK0EM20MQ1/AwBGGawZIP84ZjU3EAv1aE
fAxj+IGbKxC0d5qTW71RTVzLnAVW5xtBzruXc4gro42a/H4Y6XBMganc7DcNchlZcqt84AzKyHhW
Gt43zk04ETWPDj0L11OB6dpXjGA0vQSyn+ErYpfzft4JPJZL5FzobsxbuiUVnLD/vKOTdb+smMqK
5sWk54m//654ASvPktEGiicwusRvX0XgjXsh030ZGcFqMPzR3s+axDofss/y+P/q/ixRT00rJ5MN
9VJakfdhvoz4fKQRrU/ugMdCFFeEY8mXeGfNf/sBJYUOcPyq6sYC+/rQbbtumKWCISZaTmBGSutC
viKfT3L9JvMPFutxGSJbIy0mOWURsyQHmJY4d6pNUgTJn+UYuiZcvmrctNMzuqbEhKNFcdya/16c
7DPuRb9aZb63MDrjp1tp4Ctlp4Q+tiLpcK1ONigATvi1zj+HClo+KMh5chX9XQIDluidiRnzSBWN
ez6hc60O7Wa4OMSVUwceoN6jQF/6ZEoubbnaCGeWYMqhCl+sllQlO+hGR/J2rOc80IJtWoagWXDd
Zvr2Mzm2CbbnFmVzBRaCA8ZtZ3PIjrxFWh+/U6uEzg+ax/79gNz0sPQP/JeWseTqFrOPKdEt4XSQ
IzdnVOHeWob+D3T+qcgscE0g9+YyvATt2PHKs44EWXD4ub6R0lsl+srn/blvn7W1o6CNcDJF811W
BW9eekgaKJ8HRj6ZqAVsfvTf8XCMx9ftl8z6/03JPK7NLZ9OIZgrp82dLRHR8TNeFFgZXMCOLzU4
IkUh8AJmTC7ZJldlieAGte3Q3RoSCenmqNPkkpd/NDZJhy4fqIf3pJLyAaGBVGtM2A5HoqqIW7b9
y+o1NdvC8uLARiFdLZrxi3ie6fzE0u+pLNp+sRiJdLLfyyJ4WTTPRl6RTxp0VL6WSc9PDleAYbmK
ce0jO3HQ49Q6zr5x1Eta9TiSP5TSEV72COkPIW1zYuO+hFjbZSFVMXMIk8wzaHcvh/Hqb4avnSyr
IZfxA4Ukv5Geoq36y4pQEUaWaFc9TSNxtwnznZs8JIMabJmI+WDbCGlcimQrVXcyfA4SfWQ7uIwI
UvdKvIbzBcNZdOCO+BoW2pQhUiEcdmNWxkzI4cyX3pyVLSRemJdpzDPDmPUgSTB5cWcRiPSHwChk
EjcIwG5/cnJV8Cju3nHQSEJ7VvN6FmQtf5ncXh79rNnp6ma4YVcCHV5kQIntkRtDTqbhwcAZoz98
RPINc/xDEh+O1mf7K/3aEz1fuVpqiEgAAGrbbdyhEUWGLvRXTJS0ODcHBnXxkeeR+geK7DiwkCTh
tpqARh9P6LI8uMkaT4rhnnZIa1DxsCl5a5l9wabqR5hXE9r/OcImy30b04upNODyGGw4otvUANEO
Qo17ahLHDL9M9QmsWW1/515uYsRePdhKyijhwSmR3nsthIH1PX4zKVUyFXWqDICMY3d3hl2QM31q
T3MK3/un0WG1vBp+cycCG09iuTSfQejIY6mchGr3ZGzPWkEQdLnn7OhRQu2XVSXafDV4Ep2G4mKi
dI8YNW5VEatfk6e790IVduvDYH5vd41dvXLR554dlnWCglpxqj52rtwwcsDIa96kXBkhnR6buxA8
Ojvy8kN8dW14BySJgKREh3KK30mqTuzTilSepku/rTi4WadVi79m26Vv23xTU385PR0tOYDdgMTM
NbrA8REJ88XaYsPOUaJ1M+IMcoi/i6YN3goGgil2Q653V9jAAi2QIHsNWk7HBcmtXARdbDwuNx2n
DMbGo6DzDrn90sITUfbuqfsk/B6p7lmEerg18Qm4namcmT878ULHosjZfeKgRy/sRKQeDG4vS5pf
GwlmbROxJTpTU2HL56kSbCE6wAsUozV0O/LDJQKrWhIplJaWW+8wEWjFw4vQlC4qoPC6CSmJmvH4
I3U0RuXkKtPhao3P6PQk291j+4NdQU508MHl5lckzfKsNCo1JrjDJWp26fHVMZrNXNlRJ760zvJ/
YeArJ4P1LT1oV7tbcuItDnPQIj8NaM7Y/gomMpXxZ/D35DRYQ/nxsx1NLZEmxwVEh61QMJP9EG1Y
fzoCvUHq6wUnM6PPvnrVYZKntc68OMmPo4i2H3sAiFWhNM3OeOryB2vO5KGESqDaJ8WK6qMO2yB1
fZZkRw3g9uO48c0ceElIM6a7YxrbdX3CZ/Zs8H0OFW+hEnfKicBIVEtXm/phEYKxmTGYe+v246aK
RL/Ruqkmx62e1HONEZ15DdX0nHmyD5GSOZMhl9O2odylNsLm+D40qNU8JyXcgtm18VUjmt+GOt3h
P1Xo9UDZIleYIngH425b66JsAwQGazD67nKDNGHp+7UVSqsjvyAFvlrOD4bz3z0nhrKl7wBcelh9
AIjXCu+WKvlnPjmsNGV2EoEXovhhB7b0rUHWOkA7xpHJUrH6c4YC31vKykALbBbkRrCNuvz3bZoa
pjyQmxAcAiNDyH+Dw8EijdVd/pCC7MjgyOZwAJHPxJtmq+mM1yeGBkdgGOXZySvWIUsBOxnqG94J
IoEAF/XKCoOdLyt4y2/XKksOMfRwtGGEg307socxd84OGjCS799EypKr0n3CHUTy/oZ9bEM32zb8
iMC1863RyinCVFXQa9SZnd+F0dGGiOwSRnunOXuoDjmLllzNfSUFXHZO4hq6CIERLQJSNADg8ePU
o1z/N0Ufa8J90zG0ivsDXMbn3H58bRFKOFTiQvWH6HaBzCF2lOCA3TORpS/0f9XnQbcO97LiAa5K
bgTGTuneOVIhn4EL724C5Mq4JLVV0WAH+5oXeNeW4z2N+h/mpKxIsU1J0OryM4sxmxP8jG7AZfNy
DXNTXNpwxch0RxAJv87bS4WGFRPpTof/n9s69bziryzjNFXNol80TlJgW7uw6/DHRvkdN37bXgEB
TUmgPW+RM/8GnT4P1ybazdj6UvfrUoiKLHnYlOtpycg/w8dyxKdrBqQZflDCt9f5uLlXv5O2mYQg
eV1ry4M1PM5MQ5Ux+6AyphXTYCdilmfApBgXDjazRzGHdaW+Ckgc9ltePGFU3iaFb5xrA+wS+BgS
Vx+DtfWxqG2YJI2nMABrIWyjJHecIBStc4QgKGXGMIitJn16u6Nl1dgjdOUdMXZGQFv976hLRwZy
ROPO9gRHjIVYYbAuR6pABOONVllMug0GezZrd9aA43z4fvRVr+PvHXTct5ivCoSG24Ix8DsdYsSp
HsZgL4XDKuUakFkHa1VAAewiSaM0YeLFEcTIjNyL43IYLGloNCK1TEvsFdtEFiF2QcPyXY+GZfaB
0ZXdQBawtvEMOb2THXY7J/nigLDRMYGZL1ll04FFC7POtEJ4+icr/l/ihBtFTu8UDh2pGRejRBsC
Sg8vqtXR2uRjD3iznT5KeCKAtoSMRVHmtn6SmgouOkIz4xSkvSLS5j7wWGvMz+SXJCMCIJG2+t+s
BPRiZSqw4hyrniNZMeGRI6uH39Ntvr514CzYncF+Q+2s8VJOmRoGusS/a7EOe1gOaAGwcr0xUAz6
q1N215ESBAcCOk17fjPrSQTc8fmREZNHBxNx9UNvfN68YzXoySJrgNLjTTEy/7L6vH2+URqyCArw
hujbnbZPzz2FMTLiohBRgJie1SjWwjhsE1U1FXDYajZ/Lcd1mZhf0Pwer+E7fEYzyzeQf4ojA1ja
eeYXwgOMfxJSxfi5ahNPg9wW5TI17Mub6NvuCB7axE/VfBGCyZq3U+9o2Sw9Vp99opHk6rO9A/Vg
KH7pe1ay8IioQQJW0klHQf6MsWm5o0WEXIkd63Oooqpa/EILSLO0ehz+ERKaAFAq8K39cEUWL2GD
BKWzZPUGZSXm7LJnHtpOtRG4WpHShiZb55J7AZGLuT5sZP3caUoamqKX3O+h+WKIHgYBVDp9Umml
EYqdML5UG1mJdoLKgUKEhNpf4nW+WODRHRBFD8EkAZf3oSpYiCpbY12HiN4pkSYPUmLUUm5aIGDt
zDZUyTU/LMrz5ZI9TUHarCu4N/cNQY0DakJ5v+65p1ZFS5hcpey/uiNOKPuEsu5Mmc4k6IuxSJe3
yFT29KOBNIjpD6mskj5MByIYYX+1Pus2muACkMXyl8CxEWVQIdKtCf0ArUaMYeu6GKV4honzLu62
jRnnF+geRqueU5T1tGxhnuRg5a7yvaUTeGpmwiibhbyVR9HC95ZtHAhcra4HZUkKnjBL+XTihHbI
6aKcbNBijWUp4M+tfM0HIkXs2ZXmjO0uyaUVboPYqoQwVZ+cU/6BKRmJ/r7pY4s5eto14WFEIDnO
1a9Wg/p7Ypxas19AILweEOaP1mZN68S6RxbuhgelQySoKKrEB/dtt6mO0yaNssmWezPOzcHYlc+6
SHYKQForfyXTikQYujQpZ1jMwPh8Rs+VchgUdf8G/vtJL5jdiMvzC1D0H1nCAHjHH6dxvSbENwER
P0FTSEJHMnkJdjLXXwpbR1RQ3puxs8XVZ2PZa0pYl838+gzCvqt2+CoFDgAVL6KqUMBoHblrTCE7
QpeUnDIYoRC4x6/9YngIZqi1bswwu6A9a1WyN8jFgXs9SI8mkXvqdGWINc1H4I2D/mf4VpVnStnv
lgPgGJiFmDSbxQHTLAcqEsLbyQyrKzglMT97QEJ3X2QEryez6vquRa1EgSPgC7NBEjqv/R5klfpF
+5EKqwoAojayqIzXTSkRWcy3VDPpy7sz53JiYWAME7EMEUv3k+o3Jl8KjE+P7a38w8XnZytbG1Qo
t6cZY1vKgSI9Mp8HEyQKbKRc2Y6lmA469WR0h+DLFPF84FJW15vV2YDtLdZ6XlPopOp2XCzyiTRD
EFrtJKbLlk5G4iTyx6S71nHkmPujWu003O/8PssTzhDDQRPhWPggNebuWJE3WBWgpsFaNZdpuJCS
bi9ma3Zf96cCSz/FizUSoZ/NkMtvCV7CHUUbm43U9Sf2mcyEuzhKGw+4JTmM47SZSf/+iTh80rUQ
CmPLPGNGabp0S/YqfPTWyB6z4gz+yK5J8au1uMMDka0ymVo9QjlI+aOwQIG+Vu6kZXVznCmmFqan
1eJ/W/opPuBT9/xy6sQ78dFOlFM3MyxL/zbWh3zY3MO04B/lu7zm9SxFCf7zv2rKIs59K1KrO9qS
pVF4xJS68FHcO8QeVvgJtdw94lSkIZMQRtT5H6O82qRh7vpms0G8LwdQAZNyJCbMMkQrr7tGTUCC
Ofjxx556JNU5AYWSG8lVkEsmjhgQiukNV7Q7odN86bcWkvfbZjE3WaTj8KOkxZkmJIz415UvKtT0
XfkzBp3Gtl44oL/5Lo0GdzPci8ZooUKBN+LzIx7Xafc8ejroqgTv+nb1IuB2/TXxdHrtytT6CfWR
J1pnL7W+YjrXWr8jY600eMJb0WfxO4unsMFdgCCr5I8F5PWj5fu5DlozXlf0MDygrKEGusyCw//J
yFTIxHuBZgktHcpaTQEo3JDKi/s5v7yfBZyD+kXBG0vkeiy1h4qtg4orf5af+hIWHjc2xkbYscs9
ML1kj3wgdfkzOgjNiWwVpucaapNttgdO7b4jLW9T8Sl1P08qTo+214zXLAKaWDD7YXXntAmSSVtG
tTt4xH5943sCDLZXr4Vg/uDHy7zztzNB5hRbLudb9zPPX+YFbhHXc7eqk/z5tK8TTAVcdPvGR88q
qh56q6xD/ByrKKIbEzermdCMLO1YmYe0/j5/iEqMUge8S2JNx+v+Ec1QLw2aTvQb3k6qrYlx+1qw
bNEukyzZ5fIgqgAgEnzQ7LDaQLRioWI5SHwwircF2Xn8CLvo/5x84MUiqKjbWvhULCspuiKWQ35z
FpJXOzX6rjfGTHdQoU3m3sCAyPdVNmpyeX1PbV6Gx7RYDktsTy7sm4sC14iLZ54EL2mktRamvS1i
84u+X99/hFlCZfLrPzOPbMDajlsN7HyhzvUeslJ00SnsD1kCcqwzX47PsjoFIgYkNK4lBeQjHd/f
97e9/4qBvl8UGUKOzUKvy1UAH3fcj7ghnl4rwSJhKuOzcF5ijW/aDYgU91IIARKI10bNi8n0l39h
eTSAKRFURtxLeY6vgSpoOqeArLeIqqWTNxh68cu9cSgBexrw0bpcAeCY4B9XmUU37Xm4rkxyD5+V
EYJE5K7XEdNqiFX8xrrU5cUjPLAA5rrJ3H78mLolLBBdQTfA4Bpj4f8oEVPHkNKNhpwjHCP2ppoL
uOGHdXd2xI6QCoMFifycxvTAxRQA7PvVisI4CyaxzPv9A+VFCjukyWKOOMUroPx6iNJMUldTCJ5U
ioClhNzPYh8FQ1qDo7lhPyhb1ZkfEGJRlvH11ENlGmSi4z7rojiA6+0i5Z68QCJGtjK2SVI8vgDN
HO4UiVOYGpcV6aSPIUgqyYhjRy+h0l2pneXy6IlQ4vn+XvUnGRwqY6IJNLwb0Af2LGE8ju3ZlOMq
U3ricf63PVUuqxhwgDXWgId4sEcohzG5NhBV7OqSvV7VoI1zkbvgPw36KjCvUqHU/LQ3flHN5/sV
hrdHyvGCI4U0ehn938JfPtgeZPmvaJJM4a85uh0QDDePh3qlV8pikrCkjNZyLkU82np0Ila0reHf
FY+gAszlHSiIIkscDhSgRuk8Tka33fBLkpWdD4HY8f8/lkEwR5iBnrlyoblp1Zbf1APElPmZyBqL
a8nFz+btc/wiOpf9ZZt8j/UOIsGBtEJSFBvcpgafz9hKkdG4nRDD9wzsSwdBsO88AE+PPxKPbbvt
WCuRaNgEEdT5pWMTHz9vURpJ1HHMcf5rnSgnY36PYsc+4O0OA0Lo8tIDi6J/xHFnU3UiJjoQ4hjt
BIXoQifMrYYyV8/0ixqd789mTS2tdfWnlSnb8oiUNwaqSkrDKM9tdP+Yan5mtEAxdd4FCLKD+kXR
ym+SM2HWbOlk6C0vO2mtl53n7uF+UEWNzDsGMsU4nl6NaEeQTsBjMNLxRx61rv77ieKxlHEUEVFW
r64v9wMzi7cmaCPbl7/x/nclPAnjd71yMvwspS3oqI023HGj0DR+F792aFis1mqhNZd/XfPjOWF4
3/hEpR0skNEqDtap52EVKjVw/jtPcriE8B1rkwmo2UgEVc1NTwQEEWSLqr0bb7QZ5qz22JJ4o5t6
fbnh1e5ZebWP1ntm1JhdGfk0eFJE9vqKALM2KYbOgVeQH/9PsyOXhpnpxSSQT2tRBLh6ytE1lO0B
pRpAwvxn73zkDrPMVWIfS/W1vrQAEh7Nqkkd9k7Wz7ewObHOz5SZnhVkScJW+o7AcPGh+tXsp0fy
OTFTxV3BekvRFHmZhXAZL9wmKvz73HDMPgQidWzSpIgsivs8gJ9fb90J556W9TbGY7epwIhOKWUY
SJXK6vVp7YO486AT6bcTN1MHQzhgQDlt9N+IvYyukTCfapBZEvqsbBLtcDF5cFV+xyCTYmidzArm
+RWG83Rtkj8jqZ1XFgrKoLmCgPJlmRVuPKv1TZhr/K9Ys8+crK4Bx+lLxkTiNZ8jsbgjuRUffn4A
i0VLaj3n/C0HECNJ7Srzxo3b5sx5OBqch5XqJMoOBOy58efgimTkQFq/AmGXdXro1fu8mchkMpbD
jPAejV3/BdnCKmOmU3fNL9XwakDXk7te1WkKHhhKo+1eiO1BISRasxZNfBQbQnb6enHzz2SttGIH
pApZ8GkdNyXM22iyJJrpf0hlvLR8O0QaDQG7ReT6+wLIHyrBezJCj1n1rf0xujknAPbEO7GNxLN0
JVEMTpIRaW3Mlr6uqvK1wvg8ovevQXH19m5+Q9Qg6deUjJIv8W1qdbzQfFMm2w3VwprTbG/StuKz
sYOFHWLjNTRd83QFiKvy5ZMKWFLoA1f3uaHOpZsIYzsGbwmN9siM0GM9suOYDFqaEEiIjWF4vkUp
B+j/XcHiKQl6D390/975+rUlx53zoko2U0YXDNn7ymMpJy1LA/4aJT0cGlj5ClejWsTQDbHCHgHa
qh3S8BrDsoG+fg5c3SgvfVX8Bd1GMJ6ZuxTmxQlEthBCZAs9Z+GFsanGtWpbNMF6nthuhwN3sLPl
LX998mSL3bULWH+dhNSucF2iM3e48OvbekRUa6kvqqRZfj5vqOqyvaCf2HHtNertsa/UzQWRhNY9
H4MfFW9Ii+BFH32PXvpdgb9EaCXgQQW8bCIZYwceSG23OFUkzfs60MTRt/1H/JIDHHr9uAkved/j
GtC+mHwI4xB9TFuK8BSR1sUjQuCBUnzCe3B5UXlu1TOXyhtr1Y0U6+aqWCGrzcgut5asHSbd/72S
gFHFQNAQPRqs6ZWgMoaH0qKC03L/j9oCf3S580J5uJMHHhJrss43pOncTMMEqeuMgAdqMTKfSdRS
kzFbSJNa8lBe7rZ17KfFeZnsj9FZUA3iIpur5PpVy3DYqKRmGnZEOIYOwkVx8Bc68gvAEidzNe+I
r4rEOBV97NvILqvShEt/SjPZwYMjKHCfsgJz8qsgzupqUpCsSQ4fPI0T19c+3sR9VUmEnrIzzAvK
rpKCuJuHgXEZtDZxgazZu6L2gL9melRBZl1DPdy9yWjU82/2OCb1xUahmGLdNY9L7kAmG3/5tLh9
BWOWyuub88jC71WgtOVYeq8L06PNItvChMu0fpy+I1/r34LBGaeFgdgbBXHbMLw5Y+rnTsa5ghXY
BS74g05wWpFdn2BLL+Z5yTS0EQfz/CmbGDLgtQdOBSOqBklBh8qy9d5+c9KVmUy3wsCbzmPx8vCl
al3DWIhC/aADcspO9ETalvJBw63v94c7QcGIfXSJqABw9rEKSfZjYCFUwDLv+GVUIvlq8l9ulxHW
o/3Z2VMAaxRM3vi72WJEEs0xLSRpAvVtQilA18+0jxIJ/HshB1bhmp13XNxDq53PfZdMVHyQ0wh9
oIOZZRIrIrymvja1MfoWCHE1wGmDJyJM/lQWMEiJKktQamkd5QUkuvAnAfvSifBjTJh8vXbordhQ
PRZppt9CY/o6TUvE4GA5w4ylaHRgsJwkMPxjOugPs+KX3K96ymQhsQQaIurQcSxu1LwtwUrSr7B7
ZQte40VErTaw1/naA+JAROIKo1ce+Tkvwyh+rfPRg+khX1W7uSpAHBj1sf/ZsKl1TkFmIzD5ZPD7
PxMVXp1krcvcT7cTYybg2bm6sHLi0D+W9iW28Z1t0FAe5L1BHPIkpYfWSEHZLwtSltqVjTjrgNTR
t9HjPshLsj31ndh9J//dDeZvz9NFs9AOoWRplCv5OkJ7wPmtnphaaY9tIZAFM6m4OKmlW4e1z096
srW7kXFB+3nIfemdCUSHypx+5n8Sn3twAyUfvH6FULl208j1ofl/xxk9ii/L7FwMr4or6trWlIK/
Ur5vCEd3AnuyJc2+TdmL2JESaCUyrDH3QD+eYWpu5B0VuMwfHUlvO/TaME0o7V9ZF+lq8yFK0vTj
kle6J8pZDhD1yGN9k7vcsFE3Jb7eEnv/hD+SocHgTiJza6g+79NfR+55wq3bfNxtl4rFBhEljR/k
3lQAOQrSkCLV1OcYsZc3Mi8pZ7ALkgm81aRcL1J6Nfr2VUgMSzhP6XmRAdLRd8zI0VPbmtcWzTO0
RzG2/KY32uOFClIkDe9BwE1UzfyxTPOLCw2cAK7qc0noWibfLqmVpCbc/mGY66i9LZULF4Pfytaz
ZGXuYq4M4fHaMa1F/Nu8F5mg9mp1h48lNqHdtR92NdOkxxDnE6vsBI+kO/QxrEEG3YFi/mAHwMCN
S3CWB/oUcK9AOvuyLqjWZMU+B+6ra2RSZ92ByLB5nj0mhYA5N3bvFGqQYXkwlj+JaYlYtwRRlbs3
tjkGOZ0Oz8OAa63GkBckikl7IfE4JCWi0e2Z7GdhJ0G2lVMMVlVL3Wo8sfl+P6gkbwBGaLUhqST8
ZCtILT/Mn7ljL2Bju8bYXAsG1KoYsiW752gtkpyXYA5D6/TALjEIZxdPB+q2/yDUvcnbClVAgJUi
SlK0ySjAC2PxlSc91Zvm12XXlz8E+qta+718csFAsz7zGgOPq2CaLm3C0IL4Gk8q12GsLy2WWzxh
ZJZDTPeLDztsmwho6PZ/pXb+imsU+MYsE+A57MLQo8uaigFH8UQfP5sGycmY+qr2GqyIAL+Mx/Bk
g8WO5lFRBn1AW6IBgjQIgXvVgoxGiXEg0mB1mwtPlgFvZQwyu39oBGKvyeY9aNCWxjhhY9E5ZH27
VIxzqguZHur5R0+L0qtNLKL0l6h0DCKxueP7sR7ohVWR9EGUYKXBh30orSG5XgTqD7pQC9z0nVVS
J3UzdCnTxcsM26tzjiFeg7Wg7dB8juB7XtLjLYDtweZrkoYNWoePnxUYz96HKIrVv8MfVtHkUnH+
IqBo6j0MOWcT+6bN7Jq0oZDDZ8M35ckugoTnJWDMyqGkAj/BO4GS3u4xn57SfkFA5zGnucMtuKGG
eMNR6rmbdALm6pyZhWa0/Mb2qD+aa2r+79Ihh38gWMTazyEpZdtPHdWegyPoTTFbAIcF//JYIN8+
jzrZZnzlfjPXjLQr8I4126xbn0SNTc5pn1cjCIFS8VfSD2fhk2pArwLbHPK2/kLSH5FAR8M6GH2m
EkceQKxH12NR5B2tdkOmKF3i2NTqgNxz+CSytJSMWqe4nIfcxdRLyaN64Rf01w/YtgTPbMWfHocb
spURFqKNVBeeNy6K+OrPFprmi37L7j5pMfhfzizZxGLDM6lfv9x2Qxu1g//iLRoI0pYXSrtWP2r5
PH9js6DSeKfDZomevh7hH2Cagi/KPDpW4yGv3vvfSI2pMXAGqchwRNzhGstpQI6yDdHRatlD8Cxw
9YpDJWntn+TKxi0GpXSY+7W27Rc9eaBj7Rxm79j/bddqPnHpk3hzx8RPyt5i/4WEW1x447TKHboR
AQnXrhfxv11uF8UC2zaUuk9el00/N75GyGNrAjzr2Ze1aAmEFbtOduUlaiFCFs0HhctkYC2DDE+Q
i1T24bix/Z//txCXiapXpf5FpCUvrOFrcyHpb8mqLI18uHkIDzILtD47a6pP0TisTdZM9CQerOUp
8uCVT30WsSpVjojpS6nzgQkupwvw41nKZ8A2Ww+I8g4+gTV4FRL0/NXsxFeL0iQ4COBgJhPTX7I2
82pqYtNIcvn4t/1xqK5361jFk0CQMsxZy+kKVJZqX1dgFP0Zlei+qt/bsLbAQT8sEqTqarzeRIcR
9DzvFaSzTNuenKq5vo03Gssbr5Lea/FPMWaeKijMyRpYX6bBH4ZjWVT3wynwDG3neqVlFQwBUNw7
cNFiZJyfG7kITraBaVVSz+e/hHdIb49ZPthHQdoEthVXEOvJTfmFQSMtTTCRI5rI53kgbCkLICE6
CGaPjVxUG+WYMzD8gGOsBGnDbK1DNP0+y3EjrcOdM2p7rMTzormk0XdscSdttwQHnkilKI6PSkzp
iql7t0Yspw56lLYN7NvIhuFx0a93wT/fnb7rR0VwryqKEBdJjh32h1bHXfIdKwq0AhqQCBQzBQOB
ObiLQDvivj4KXfdAUbCfOGXvihXXKj3jKDUT2dt2oClG7OgeyZrZsektnaMKwPfWV3s8gZ/HkAE7
KDQep5onh2wJscGDRgX0aD7rPpvyMhKgo7DRtF6+N0hAVhs3v3G/vul9HB9PO6NHWkajwi0HhR+M
eDqje40N+XcICr2HzGdhxW6dtEArko99n85Jxvot4yxVJckgPdL5kTAV/xVNwYtbzTzKLzIfuMUI
LbEWlBKG134y+RABYEHFEBgdgVdxDmkvsNUWl859ZGWbkBvehacJiaQFetmacWZZTq1HYGe4TTWY
dd9Cpeh9RW56fFUVfYdIRVWxlAZIgWQlGP08xIfd/vkJCeqOou1Tn9rmJgW3Q7/umAMTni02LHkW
O08EggoVC3zyZek+ZzcNFLSE5VJIHTMWxFjuO4qv5s/EnRl5zCes/AWz4K4v7BWwztygZ/GesGns
tFpnwQOuC6/z8sBKASdjzNZrFCFh55C2j3EwZ+oV/FgZlYD62hUmaPCjpt6tqf1HcaFtuHZwFGnK
uT9NlXiKDFFLBkoqsDIKj5jaygAjX+y6r3fZK8WWxT5TfmD1B3wPQ/OJhpsDhmN3cCAsYbweniLa
UzjVGO+3VEigxSVG3xZ24jOeeQ+/CbK3qDHqnRNB+oJ0YBaFQ07HAZvduy1P9jRJR84kI3aNu1Tv
KVsmgnL6gLpqgmpG9WE9+fFkq0LgxreZUUBqgQkf0mIPw74EYRlefgLm3+P6V1t1ziMcgRgYSxxy
gwDoG408QEpW6XuwtT3uyTrBIjFRjUl9DOJD3vCBh/Y127g589gAuor95iYbiiNW9NGswFCIEljg
G2MTt51gw9yZE5U3d68m31fJnTfX/8lunfxDoBWl2G2vds2q/WwovUBtkgyo/nlEWRealGsoWyaa
Y1o9bb4UBpbfN/S+87M0DOnIYGMqufN2Hbsabn0mmNCA3GLLyEMkNKaX8313KcoWNQy2pq+MKUrm
NjUXdLyroJPkg4C9tt9N1IGfqSfvHedgijQp5+rQOia91U9s19fMc1XeTNCLCMDMDplgBtLtJosc
uOazJxhQJG3LBTmi2Q+H+ycht79jwDO2lnSclZLS3O848KuAa6lyUT45UZ9htShzIXqwgBXhevR0
Z2A+/tKVE3IwpBcht6J69MXZPcB37BBUQsvse5sSc1mKBowkUNLeRRos3iccvDq4My6lzNl7Wr/K
KleuFgIeWoBly/9YyKfgTd3ej7BSBkY4MOoTQwU0Y+Ua7dSHGqzM/z6Xm7osMQGfV+T1A7xioNJv
6nXGp78/DBqadoWFphgQI0IL03ddlbDKJiQjgPjQeWW3xnsSNQ66IGLI8vHgz6I2rGPQ14D8IUAg
mInB6Ws7bj7qwIfS9tNDKgqKc2KmOZJAyoD7yid3tZCCw47yYm0EEIZ8CJ3WO6kJrBUqfwCRLFUi
/11zumuyhdq9WEQKacpbFweWZdjRgxA3ZYGPHt2s+3muBeT86t9n9aXBN7ys7ASs2U+cdPvaJNNN
w8qUKxOBsA+YNJGm39qFWAkC6JUvDNebgxvM4K0Kdx/8wGSAU3twz8HHyc5epUz04tZW6FKJF8+e
dXUlNkH8Brfedu4DWNNfCHUZFl/KxBXMSJd92H6rr8nUqhFSNkKMB3SkE5/GeOB4zfhvOMYJDqyr
puhHNS+PpUs22wEhUJyCOYC1qS544d+t3BNXGooqic7JFYHTZJg3CKMsn9PRHf8Z+JzTZAB8ACNF
2E3yCkmTCpL0Ofw2gizseMX2O1Wj2HxwsGU8t78LLuOcoytSs8qXeN7PrhqoBE3T+ZbsL+2ajr/5
Hg4AtrxX6Vou9wNw6USE/vluByGXifhGrq3IKVqtmwlmZ7QaprQqza/iX4vQAXoqetTF5CNjURqK
dAG6Y+EGj7ULz+MPO+5a1seAHxP4A0yE2ujoacJVQRaf7LApbcPitpHHkXLixxY5W5IcYe8+Zp6n
MpyCVgSfdT6GfPdse8cyXF3cMavyPGLmVHMMgzVhPHY+91ZVBYitze77xcCkF+A2samVYoB4rph2
eIzlX/wovNiLUb3Dgkk1JMzPNlhyfxQxUA9RgX6jftlZp1GKuxGMi5KpFglyLdLxkLjj/QGBsFmQ
TDeAf4iV7QCJO1VP2WK9Y27X6C/JhYM7Zq9rESHM4h6x1aOcE1u3d0VeV6LVPu7RkFD+p5C0OlKB
FFW38yWUI/5LqbYzBT+3t1JinwLNxDu6vodNHR/V83/09eP71MNiF75+aM/CRVokvqnInX8L47Qr
lJiP2fhedAtS+EsTz5Abth9p49E9+LOtcPdvoDb53Pr/gFITOp7sD0JIVF4bjqg9l6jzd1IE395J
+0tvdU9bkjPG5pCratlWj3b+chvgqQFNmjD+98uCA1KT/TUIIsXY/FX3yppeQn4lefstQEdEWT8A
1291dwhfuUmrQXr/ACRvh4QQ6UPuArBnggsbyi3vB4su5BN4z8lhe04BMF1H4j0QmW9JRIezCbL+
6X4g5XVQidgRyS9mrU0h9j7F831qyymPGVqcs33keY0U5SmvOHQHREbvDT/aUZ5GsX+8ML8/DLz4
MCRpd+tzLAdo5yEUGyiARlkyONAyai1tOPibD+1Pcb2cJaYQXWD7xXEouws0iTD5UocEumnegPXn
q5Y6dP2K7zdfBuv2MvfLw1kYFrnpmM/zpYej03pnZgf+xJGhMKtqEiW8A4X36h3rfAil1j+u8LP3
a1QyZqBSloT6P3lTTOvWQeDsBzpNL8R2OktDlPqQIUBZ0XzCtV06jmPNYvBqILyIPj82oopyTQEH
zKnzNtkcR2z4u+E9JT7iveFDSf6sQ4vE9/kHx75TwKZLkKD+uP7dERwdo17iLxbffORdAijqxbBi
7BKZGKBlZp7ZgqHe95THLE0yI7MDPbn15Xs9sbOKfCxDkGEfhqteHDbEjqY3SQl6Vs90qDGBdpWr
rVaWZQiKqzjYL7EZItlxo31fRZ+GVxZmyC3s7xX0cnwQxyRVgFYZzhpCBgFzx6QbXvaT97bIBiwp
OJ40m6gsUsBIO3QPduJfIA1Jhh3x5HcS/1R/IQ9MzVqNTRl5Z4XElnGQMpPnR5x2jriBILyurKT5
O82j5ETgsi3jMgk+yicUKE2e+j4c5Jq/AgQtlnERTso2M6GtSAb/h1+Aa/YZb8Tjo8anbnf/Z3uB
ScS0pjinlj+wkEgwJhgQ5irzK4dpZn1n/3flLzUs7Q9NrVIMXHLAMMx8IlNinWVtkIAprt946jUH
uLzdj3KDuk+sxrGjOWuiIVO5z1jpdWH0PjTtv5OP8HwupYqRA739G0dxL1CpL+fpRPOGPNh85oVU
8/TzuEuMVIBXLAURqjI1EYfDrdQHHi8ijLjNwpL56b6/FuuIVr7Y1Xu1ThVzR5ahEhUEsvN7MLOO
jfJ43mpCrVVpzuSkZxJHTypscu3F91J8crS2RAqbZqaJaVFusAxFmZS23zsdiS5yVyGxvjs1ULyc
YdbPrRc77Ra0fTe5web7V1WdoRtCDz18G8u6+KVrdsoou8v6wpOeRxagYkHLbR+g6DsXyIUWv31I
kGWkIiws8Tlpxb8nlYrPr7krUboaz3QhzcU9BRpqejiYzPYENvNgsrsQNHxmgBsWGUOlPtoS7ctf
iuM4Db8/jX0qORb9jhgFozmc4Sm85Q7E9lB15LvonGeJX17f6JybRMnZJdPJle0YF6cAbuwlNIY7
u+HH8cYhA4HtcErsLg8PzXoI5jBxH8ivR2mtY25WsMJcMfm9TzLcafwBIrIXXoo8yIuUREwA3AH/
/+hQ8xK5S8pGOFgTwLsgMXc6JmZKgD6OT9bPk3nD9tm8HVCFLV4UpAgslYRPvYiF9aBumi+KTZ/J
qtadT9nrHCXPIm4ZPtt2ts3A/gcQBjdnryHNzUguxW5RMhtThy8btMxCM2OFrr7/rjSXtYwV0mbu
HGgmeh2pf+6suastK/577jh/y+gbjIcx1d+5eCqwIvUfoL9BYOkMokuiFGt55i1JUJLXVMPjxGeH
7UDCQ5r4UDVy0x2xuzv+CYKhE+XA9sLh09HtF1YtfdAfQzEWsEH3C8syZ1RAzzOqK07aR788t9XC
Kyl1SQypL5C4ixVorg6kpfu0V5VZi+MOiEzxeL2WpiQPC8RvoZUQOOs1YhMX45mO1+4XdjgDuBKk
d4hUJErKzGtvKItSd2PJHXxPLBUqx4EY1Ynjx1xZmeeFnQIuNl6wczpWbZapWK/LqaGUQJNTe0Dz
RLRJl2HpeNCXEq+y9240h7QrxzChxldC7KEVdI8ryUh17ThqyvupWquMu34QC4pmqHEEcOTENHqN
bTpn5QhNmdNsxOsbf2tIBPCf4cx4HuTpiYdeALouFCVUlazx5bM5J8hOVBbmzKSO39UcTyaoGAAQ
np9OO9IiWYygt6q4nyQAN1hM/oXJV0/dFJHHmDwNQQaJG4SfQ2rhJkDkKBhE2LPXBU/D5pQaN8nO
gfyKsN6plB1HFkYlrUMzR52+yd/fEcZnxu/+qrb7Q3KJfV5YSCBQ2DbDKMbFD/uO58hdPJAbTOGl
B7j9AZk9JLDkZbqqsDf9SQYVCbFqpnyFxRZbngx33ptkPCDWgx1Z/sLycl5cB7SjZy1Tz/vNkgrt
AeKwlcfaOlxBeMHen+3xOdx5bEVXMMHi6J3DJyIjpSnHCBI7uSron/k8kU+T+4LthCdMC2iOfFb/
9iPY9t01I/zvGpa/urH9iI627KvX2Uc3uXmVSrEKUmn686WMZpizJlSkWFhglWPFpizmY91EVi7k
ygFxJxElNmcxuw2FPqtkXR8fF4U0M2bC0iMP8D+VPuya4Q+IUKt/kB/Y8IjIjuK0A2sa/w2mBwEi
TcnOz5Uin1NgxQokJd1EhySdZpzZ0h/FuGN0MFfpmXbfpRdKVdzDr6ghyMNxsv5hx78jDGmdJyY4
uRSKLxiF8idi8MyClPcVRNygCFjNdAl1ebKCt7JTCGd/AreKgNxNAAa4sTFQBa+y7nPqo/LdKZWJ
UXim9HVk7pEROMpSF84q1pvN+soqE7ZwTTmtySYCiro8+tMSFJ4fu+EHXF7HC/+iCbGUwaXkTTwZ
l8qoWR9fOqsh95Sz4Cnd5AP9fYgr013U54HX375QCylt9AlvcaNqkALORXLHOY7c8j9ynB4xr0mt
QAb0GwKuETsKXGK8BA2uzfqSU7NgmueSHA4a7xrr5L/wXB+TG4TwVpcTd4K+oOr2rxJPsjolY6NT
O0Cy0Sf5JuXNw+LP8rg2yjb7BjVrN/XGIPXxl43jOYxm9MXLlcFxSph9aQ+xCDE78o8FwdU0ex4z
u3d/+6ZfAdhELtE5HffMilP46oyMSLS+ZP8r57WdDQWXMzTuW52nfuOeXA5oxU7DJmMwS+C63xJx
MWmHBVFjeR2hoY9p55dwcEnu11Rv/EocXUFQXIY5etQmdshnnyCDTlmMhBY0kUpZMnX0OZ/2F/Os
cobDUkvN0ek/dFQkDrIBz3KflGhr2lqlxjEbvJ8XeZ2MR7WAuiEWHDLLRoximCkaPROJ7xnyG8x1
x63xyKU5JgT9i2XEsft2W9XfA2B1eNX2UijdL4ymhFNn5JTCBOFcgPATwAUlg+xhOR4ZsjEDxWmw
ht+H+RTSPVqKBVIgmRRskkhCWbIbA8zo+pcdhOwTm/MgzBmhpcZ4bXKWYhrFg+81y+2d/oAHHtwO
rsycShL63IvFyD9Kv8RLEcd7mz+wt5NSjHNAhaQo+FVkxR/YFqF964cwu4HalmAowuApJs7YAkOt
LZjRJebyWb66lAFpvUDBlj/382EfeImQt0ZWdZVoo96Wjq7ouhbjPInwvdnh3xRwof757fgWYeQD
tEWGPbSXQWodZZkLGZ5CB3wLnYtP0RPcB2nrnydtc+GjY6vpc5YUbyc/Y7UAXdbTZGaM2WVXl0my
z+iGJH4BZxB/0K2mxKyx3cwKMH5ByooytL9aCxYvRszQSvKL+ceTAznX5Njt+NuaNxW6Z5WIDQlO
w23ER5Zj/tEgcq/sOSBiFLtjd0SKS5njwIY9gHIuIcbH8AhRdHh1SMlkY2SU+eQWViMIpMrNeKSR
WP5ym0qbpmnoHzLXd1JfMuR7cL5C+813qZasfPDyhOkaUeOAVVZPXetDPYnUZW8C0HjyyhF4Su9M
Dt4WFmyf0WHNpq2dly4HConGklDdsrmU2qnBX+YzgH1Sb5hy52ENmLHhw3TCVib0jF0eotJUAJO2
3IwiPVODcHQYRPTvrNxN3gnvI3Y1KuOePpCPkv+5F3eYaFXEOCth0pwi2d2mfeJc7TdNsXKwB2CW
MBajx+UMv4arZSKufLu19ZsZokroRTkM4C1N4Kmdpl4z9fxaWHrXtmzItwJWsLrXchCm4f5kGTv3
2xhyoy0TpjHYaWgottaCobZIxeqLDW073Hynv8TcrU5JeZb1BParwD1x1m+HCbu6Zflrpm1NTYUS
RQVc0f+AELD5pxF9qcVJm8PCrYqUyQ/YHlRYxtipmeYsl8GqBgV5dDYhPyOkf0EWVm2R9oiV4I6i
jyxIlkfHN6oQpHhGJBYRJnOSUHoEbMe9lqmI7CMEPt4M0ERrclNIzmQTKfoGQ3uFXGoFHfo7sRlA
x+mwTvlhp3+Q53xBA8pw8NjkOBqfKZQ25+K/2NdFu+Wy8hR9Cv3UBlIgkxx/PBTB+yhM1ZJ7s4gj
hafH2Cxzr9njslcoz0pyWlEc6WW7gCQt9AD7A2sU6G/8kaIe5Jw8RQ87LmIZonMNZt/+mBrBfYyI
g/k83kNQ8KoRI4hmqcU5ZYtNskAhDKxqOvPjvca5QPULKSC90hmi+zIm2ZXJmx2aOQsLRQ1IXmn6
lUhx0KRqT8eUq1G0KCeLPKD3EMXbA4qCBVcLa+7n4CUzpJRXn7YpEYmrsjZu72gx5EnnEp72fVIM
Y1bdvihfwkgxqaL3umhutcMfIcHupA1nFedXgIZOs5xqU49Jn9eZYmcXjbUvOrjNgyyB0JqqVrAK
D3O6IVVhPzSOg8NI0ULbJkS3hbIyeSLXSKVhWkrixymeglCkc2nQ0SLcyadZgQlsYlQ4/oHloI8u
UMNna5mhttalLCAx+duCZGama5Jn/mvsXME1MUip0hVl3oUVgSzstz8kl+9FgY/lwAv2yvaeKbQ1
gcmVn8YM9cClCpeFq2/Xn4l2gynrWUk4sfvZM1ySBzW+HLiegQuh+BIPgCb2OXnfYdA6XLgYhv3X
6F4jo3nNOxCHZYVklBFEAwH++mkcizCFxzKQeQwXwdonP7XAffO+kY0hSFaqvIrZXNfO7T8190sJ
r6hmg5xrr2shkOg7C4EBcIvIoEli0Df3l/dq1xUEiWTvDbjS+he6FDmfObwoCw66T1dTuxDTMNkO
YBqcNpl+1O9VeYPiojJ2FlHPrLkQe3frjEDV7037etHzwADxW3CklOg1ISGpnJvtv82wSWbDg3xc
MfPWaruGAJqc3l87+q03rLSOi1Z1sSVTPWEozb4r7WGYSkVLWrAbigU5/MQEWtjw4ftJRN9LxwS/
lOTnabYmOwSE0ymEQRMLBFP0JaDvy97338ajhgiqvxpuhJfuJcfoMmQp2VVhJBKnmrhuSNC13Vj8
6qcjtT3keiaaWI0rGENO4HJR3KXYWa1srbEOdTkd5bMaAXwc92ZfckiwzHsG2a1dBumze3yfaaIS
qOn1WzrkpoSWdudV+bswzRpVor85uidTM2CIsrSLt9h571X0rn7aLOXs+A7Ay/KOvOpCUkl3sUof
j3aZCfAxIMnPALGTh65DD2p19EntJSdIENBFMA6ceqxoBQ7kJ+9OnPdBZW+nQTUTlb1wFdkFQ6FT
rI1cJmklK9ItMH/5EGXwRbwhoj7nfb4CdPWhBxtZxblvAArYe/PmGG7GknBE6i46vuYqEjTl1ukO
5cnB/SFR6ldx2orzfPe4uym9Q+CvsYi8vJWdv7Hvp9T7tAAhVv83liS6GK+cmeaIcbd5hQdd3E8j
83ah6VQbEHYJjmoouwBd6tVqo8kvZnKMEBs6NOMZtD0rK3FPoKWQV9/iv252wYAxB+4o/jqsVFeY
ugroKRI/RLyk7MlQY0LuOkqEwC8xalbH2DPiYODmmKf5NNgqhJQrXpLP4l0H9bgDCvNRfnYjG8Qn
kgNs4EmCYydK6MzhiZbNhUZuwbuZT68Ue7vRUEALyNW3Bcy51guBE2zoC5n64VeY6rwRzV+0ORg0
bc8BcKanV7hsVhvYi0dmuDcmPl2JSekovvtvE7sg3/8mE1wCmZZTmyOqI8hmPbwApE2onH7iypCt
EIGBRy19cX4tdDxwBIwD5Rm/8E3Do05FKMUg68Qs0iP9mvehhMIKw8M06Hb3L4oz9rHvRNTf3+3f
8/pQNXLt1tgkPXg4kZY7QxK1HOj119UJjybmoKRta+zz/x3+SM6Ip0UdQufs4xiOIHciT9oc7qWx
g7ARPoGHvmInXno1KkbutnyveKHgAqM734L3ePd4KAkIEzPe5Bn6S0fARCmxsx39h5xFxuMZIMQZ
impov+C5kmcBC4iLloG4Zc5m01knVJucUQ50KAsMsm/RvJSmE0Gxy6Q4OJGdj2RqyeKZUK3H3xjY
Q02iNx4cPyidVcKx85qeqd0FYcOPZvODnysRm1faWFT6wXZ33v9vJI5+G/9hYz/gg5mQONe8C63B
pnEEzVknvN6Q5GICQtcY0f0ZlZjl5L+4IvddSByJ+L4T+ASXh352FFZdqGeN/0eeWQjsu2zKOB+I
bug+zbrUBS7y5qmGQNFjYIzsiSWcOI20AfTDf2mTpMQaeyefsX5sRrTKbYDc9JmAQyt9FK2QgDWu
vLtujY/wgLQdYN4SOFkhL6S/2bMxLFx32OXrHvNB665IWDdbiNuV5d1oEaH4XEPLtFHV7jsecgM6
ByU9zZiPF6RbEkV2JJMbx3UWRMMJ0sUgy48WXK53zTeXF+zBvF4r7C4Vp3uMYJqYBHi6sCC6S3BU
/JsNXMXJDDUHoz7IGlSzCj5mU7KXYA9hVRQ5PI8xz/w6yFPnhytO2yV3S71aSd6T/N7n/uw9MWcl
aY3ZEfeEKAScZLLMWCpG+VzieFVDb85XmtdURQcOIB5g7d4nwFCmO2HDSKEp2UKpYA+CG2Vx2AC1
+/nOyA3xv0Y+oQntGaOyQvVVE1qduNXgMAT8cK5C8aY9Bww3FqEK6VK/75oHKXEJpuwPn5f+jg2C
5GBBWeLQwXoF7ENTIAfI7Upk8SHbXs9e4JOToVIn+SASroAzrNBE4fMdJJZdLHiotfjnRaAXiYkW
bTswHeTWS5ercPVp6todCZrevu7Xr7QBurVjzDYzZ+VKFOu0fg0VyLlj+vVpZRbjDd0mn91Eq1OH
4x4uc78xE2tOdHDcre4kBaB+Tg7d4wY2tw1jIcYU6Gp55GjkJeBP8+2zPlv+1S04ef5Hj6QN/yDe
xhZAhcaRMebkBC1bMglPepTS+IT6uV0DTeNF4i7oB9x6wjfJA2+Eo5zHIunCA74wiRVxmMxdaJuT
fmtWUuFWzsQr8bAxAr95gyWggUkAfoTJd/jcC4xSrt7IjymSDWB4VajeINvJOI/CxsqgXKCsudRr
zxhdBfu3kyrv+M6ojZI/9dDPRRb7uLxjwV82YrWXdCxDeN4o5H75tYUzCTuTjNO1HmZbWI3HxLC9
CLrCev5F7vsgNYbUBVlto/659sx1Wo6JBefKPtXWAp1q+m5EuPOWTevDijA4OP+DT5SuxTmXurwr
rwCerIm/ESzJ9l5PhJoKKmhtNwPF3yUgyj1MIdWQqYZBxoWgTd/oNSOnFVDk8mNiE+zPAmNscElW
ObQw+6Nj2bq+JTvciqQfx2eTLfmzrwkuHrjUsotQUuIFykZMapsxbOyRC+Qw1UqO1pFDUQZGFoZk
4QA0Nj8jt/oGiQivnEOl7FdBI8Cv1hYggUzc7/07gR4P5yiqFQHSmsnwFaZRTNWzBmHqm4cllUmC
0gUKJ++ZOtpbKNyEwFgvRcLtLDBd5Tq1PvOd+5w4Tf/pvyBwKsf9VL2sOn1PVeGZXLQ4OyMQHUaf
xmQnA/8MS9ksZ6uMjf0X/hsPY+RU73C7ZjBMd5fdXFFDwtUnN1O3XScKkIilVKVxEjtXKGiOX1OU
PZH4PbTQ/Y/fRdIWhtAmMH3UM0z7nDqrZiosYM7ceNyDEpP9MGxNo/H2DwoBtYWOHIZV3G99VD4E
Fe5rZLycgVBK+161/Lqj23FW06R/wMK/WyVn0Q+TwJ+Bb5syzj28+YxBiYtt+BnMne9yoF+UuDJ4
wPq/Muvnubd5q7Erut9tjZT3nBST/7U7nrp2+EyhTRdTmUVi2TpYMn9mdU14U2cv64yzrTcX0Blq
beQ2J3+Tzfv4iQSQ/UTWLTnVlytjC40JBlnTLWcxqPAcmwaOfwTp2gg31TEWVbOC0267jau0p6Ww
XDIKehiNWFaWXKiHpB9QkxnrMiqw4mk95ubNLCpSNqzLzuoP0n/+zAi/lepBErYDrbxsE7y1ScaY
jW9uiI7Cx9PU/YJHQSUWpm01Ab+rlRrYGcvodl+8f3AEKryspW/mZG3GC1ovhGuUpr9pUiqppPVy
FPys90001wnhyI+7ndmXT7/GvqcveXlKqJHhKenKgRJ0UkqjT9iYCp0/C+jIexEFNXENvxKFxlHA
0PwWYHnX0JkyaydLm8NCNehMA2/m/7IYKGu4NT416kjFbpcpBIT/nxV++RD9+39dppp3/PC4kcGT
eWkMNGQJWunaNE3JdOiDEaNV0LBaMiZvn5fbVZfZS6NnJHUFUI0AZs/lkyOpz2RyvDL61IxvvMMi
SQMVhjQKNDdcW8xw0nfmG0lcUPcRK8/DmnTiq3OYoq5kpKn5lh5mBK0FdcE2eN1ZcuDgRTUu9/7c
sDczZzZrMD8JawwoDGXvhUnX/8TLu9owLBNwXVFdw+BunWr7ijWcPkwptYhpGtAptk+WR+/DuUbN
cd3rSyFROKlS5s6TCNSIOGIESlRMS5Hs8l7Ds/XbbJkkNwGAeIDGuPshNH4yHzMOItEYUMRd4IUh
cLPmePosgjcBbm8+UhzrzRe37zjsYHoZHM9wuaKhetnxsNKvDbIKdYbdbwnjyb4oeI408Ag2g+Jf
OB3PqI5EAAYZzlTs3G8arwKVqiFUMZVyReQ+e7CauuCWf0xlQTkGCu5Rwx2lnIdK4rGeJuLVwEd7
I9NNHWcHN50CPE+FE8OVvDTX4C/aqAgIc/XlOKo9N611TolrK9UNEz9finrvIarS8TH9SEZd0VFN
zdDeXjOyt0mHwPzclZWem/7h4KVUCd91GUK8Nj7Iqt3vSQ/o7WIE/xNSquaX2M707v9BoI/4T2if
URJwJND6SS0iV9OfgM90GEcuSov/kFSxfYhpfrf4C7hjZEFqpYbeCWnaJNh+l0CEQJyLZP5w8uQ1
13z1wlgZ0lr3igvocyvHbrkkKAlfTjJJCkGSXYR6l+VSmzdpT/X7JOrOH3gFhKGNoj9zeyAd7lzd
a/o6ByG19ycUXbe+0cnDrN9xJzTIGRgMQWkZGjJdnjwPboJAnXfDkvAHz5iHVqcXO2lRpuu7R7VM
qAORcFaBn68lHMvyYAySorpmYIJUD6gCfEh+PttgUCcNWtNR9UdlU0Ga8qhZnIomgkb1HK6CpLED
/ILliyJe9i9LM6P+moCkkzkGKPWNTibgpAkmZD0HO00Bigjy1huCXvZS4Aj5BWRLP+V7Z4M5zqgQ
5poPxvo0d4muaUBaMKMwk6hAvyJuL7UE4DmdSJxycOaVrSSlPf34+5t2YXzFnmgMeOEefuBkVG54
G/Ll7FJkP7GhI14Gfa/oruP7RWWhY0lpbQooUvyTdrxPql4xLfUlkG/Vx+2p8+FzstHAjaF2pQY3
8iwR02WCWOwGWZ900IFr29XfvUd9G9a3LjvH+WY6JCqI90c9a2b3Oc5VRc0Z4hjGADQjq2JJ2lX3
jjW4EKOfmf/LKM9QN3HGTgHU77gddNWI0dDARpWnJSBF+OQ1DUUDrgBiBThwdVeAg5j9h/sm0TCq
EkABb0q11DY7CTSLhBn2iP2gHATQ8aIMqmLNPILO/yKvTuYGusNKkG0E4LZxdYBgcrbdv9snY47E
fWtSj2xixiZP5uJTJo2IW1AgVN2vOOjcZkPyHb4M0U4h6sARuX6s22BqgdEBu71KR70OgtiSISD1
QqpbEhjztHlczq1xAZ8JZGmEvx3jZCAoiVao5X3Lpg7BiUGUYiNoc9U2C65S8UUUMlSSpxhzPvHr
Hj3mTTsdfe7kYavOF6EilHPw4Ft03ZeFA+jGFX1uZsX8CkDIFLOeb5RXrCez11a2rHDac7sXAKKr
+kQt5QmGPuIIoZBVI4h/+xXDY4rrQTmqtzi9ArAWzedO36P2RiyPrI9cof/0RnKsIJGtalnzeWYO
u/dBwBxG1w6MLzc6aUBdCnAVgL2i8xkV2xyTvpCJC8tzeHU7Fide+7AxHQAvU69CnXDmKifX5Lqm
8s4n3irum5RNYRXmOyVxL/R2NJxigtf4FnUljRohncn+e2TGXRSmJ4t9wNKj1UbYPsCmLKlx6mlD
XUng8RHnBkyw3tm0ph9O/6R1pfL6k+ptvH1ZHYzF+oh8jYOi7V5kpQESKWe5Lcw7t8wzaCRMEJqK
9HWa3n8Be7VylNSe0nNhT7iabpK4a8faDOkqstKGYdlq2K3QUBDLcrBmRR1HfDYs9j3rV4MoUhU6
Zckh0jEN2r2WAsAaXNC5Scct5NL9n+Nr0UqTkVmZK73nY5NWd2DEFn/zq9FKfu0B9v9AEbxUYHD0
27/bmBeQNeXY2ecKOCKqkUWDtoKE04Qwnxhp/kvBsNWET10K3QVkOlDR+33kqoFA8FWrQUrz0vr0
P+xjsz0Cn+LI/FEGjFLJvlnRaW5Z2+8mpnwmfyXaL7xJt4xhQ25l9lrcVXwnUgJ+eQAJ7uISKc+5
T6BsPQyQFZfDRJ53F8eTKrIWCBqFxcQh+NZHltbpNS5mwGMSlhe693Z0iL2iy4OdGVB9dO7zukdE
13PV3T3Q3OzeFyt1s7wXckiENS897kvXZZbmMmYlxFEQJYr+nLMyKygnPYViggrq8jufNADgZYqy
5MU5ZJj1wx2BMU53/AgajkuIhiYCoEBeoAy1hA9XbfN4pTkqjIrajdbryawl/Nh5dXF5fQ/sPBf5
3TtrJyYF9APrftxjg6XeTAXny8Bfi8UBTu+KZVQvURgde9S0aL/RAQKCnj5K9ThZK6LNPf8w08q0
sgbKc8aLwL+YRgYt/oN9btK6OW62/te7VHerNvWaO20F0IB/PfcxUgy7RMP1rVB87i4Z3OP9xY9R
CM08fpq5TXeBi9Zxor1z7f97x1/IuMxdSTap/pt8gu65ehgRZmToygzlu40KoGrr3rU2U+KZAGhA
ZIwRiPmFF2uIHHpyncJhWR8YQFBndNrFRcDCy3SmAz3tl6RyCt5yE1ZPygcgDDFg1T6Vn/ySumfn
sel5n+ZDBQ2YdgKeJEvq724bWDSsywZoV/zg3mdzu2fbh62qLc6rUqO0BXWvDxtz2KSDI0uM9Kh4
6GzO/mRe/gSOORdKX80DSLv6ZTR0Wb3gpfsyXiZmdfnK/96FKe088NNlyfdE63D7lQ5Q8HD/wu+t
rO7jICEVkJoDxD620EAeQHF3vRG7YR/FVYFSwhU5kIqKbjDefcwwH6PivHNrh1deBOhXOVfextuL
YX0bOOzE5kN6grIAKBj/6jG0qn1Riz3s8SfMgvWVxNrmE9m/FYh2gkZ1WyBL7Uuv9qqu8mClrl+e
1bRpJZ4Sm0VpORD4pCevVfXDa7ka1O54d1670U9Pblqe832ci87RFdfFNscBO32MmUF6p8rS4WqM
qfIF37jnBM77JCdk0hnEzXrDa/QWgx7QwitUeEwYtBUh0GdbOsGmdVByxI5sLdSrcwNNNXC+EoS2
pLLONRd12w80axz1O/ImVy406bf/VekN2svL22lEfpfRv12kn8VZqqCnSIn/N9sAw99UdH/yY+2d
0Bc8vwQ8gwzhRORiyqThoCiY9AXzHHGADCyrr8NhqqVEMKJfWfzj/Qm+xpfaQ08s5Xy17ycyBfCH
wGtEXbTtuiBjnXv18fdwSnwY29gI90iQ1uxoKJWqnzYmO4EhlOmOZFhLKFLEVYfXPl3Z8of8oM9x
hfhWN6q3En9WPxC1whrk8TEZqYAEs+pjaW7epbCxIW8mx8hNYaIMKrZIn8rGIO7IMGK97/n1i3D7
UcrfejNJKzX4EP23ER8CPugjx/EK2gzQ5Ti3ujGgnFrah8XHGJDIcHtIz6Tl6FM5I2GKsWvFszbJ
GIb5OEpwmRWurr4jIW0MzhPDz4eZWmgKII4E4Z6zQD22OZKVYGzns7wlb1NvCOJ9/kU3h/Ga26A9
F9qJwjm+paSvjvnQknhjkNZE+3deyi8P5Qujsq8hbWNLfyVzN8ck9xSXFekud6lUylNCuYgbTBbq
aVXbtxdjl2tGTueq5dS232Rg1dFkcWfBjyCeWxYVRYE6J+9wVMt3kWsn2r3asxVDVyVxZ9NzSMB8
t53BeFa6l2R/q8xnrWzoLXZMWC9TXmAqrv2vhkNRuiJfUKyjxgO8esW8Lj4K9qvS19tvVKOGFziA
YxBirhnTetY8rMolsOoaZ5Wi/xk7xV1F3LlHkSMrsAg+AdfrrPgwFlmfcvBlQgcSQCfIq7WVPgjr
cA7+SNZUF4hoXsSvBYUIIedK8u3ASikyIX3A3TVGVzy1iDgXeTCNoga1/28eonLjRThN2qURQgtI
wHbKsKXEcQJ+OE5Lg1+92W1eX46Pp8MDyRvIb4qhUHZAD+Hb9aqGQP5veikgqtt+z2arYDvIQvZz
EpZyet5cNo54Xg6wej+8nn7yxQ8fBtro1Ul4aTDXQTsHaHYYG+8LnIQu/v9NRcJlcmgNHedT9+qn
UkoRiqua6oRmnrxQqHaUPDnsf2xmYP4VMKZYz2M3bKObsj1FQOao+tPLp4wptprfGEpuuok9c99P
ROuNGwkKGAZ3BnD9ADq1Sjxh4/Gj/Y5xACf8AgYgvS+VFU1o2wiqEqW/Kiu1HVGDfmpEO7isvUT/
Mdmj4OtMAtWygA5zu5c2/yJnzIXhwlmWJ8HiLKgM6AhZK0+YlRHu2z8VGy2Xu0gGMyLXfYzDPoAf
cDruYr1RfhUAIUUlP58krhw1pup8EvTzcxhJdWjoYsAgXZpC426iydgpknrhNEYJUfjvxAlDBmZ+
dn5O9zupYX2+Q3JumRWPZN+YsB1r7SHggIjSwwyuXw8kmscU8n/hFDOCNdlsCE7nH2hn4QNK6pK6
HrHlG6jGE/wi5WmR6do4UFCwd0S+FTYWln5B8CNRZExYlagItgsxo6fFXtxv2NlD+8wyQi5PbEIG
Qo4QC/1WLEgHLag/OAeM55ZsWoZqcYhb0EQJrcrJybfOJwJnQEnVfWPkjorINT0WEOhLsVkydtQQ
ZTKlTdLSbBCxMKZOgd7zR0hqrv5fZO1tXHDDm+6Qqy955l5smxya7Mh3tNT/uoX7LdKida2/y6T4
z1DhiR2/iIFf9VexBMG9z0jPg1cZymPK1H+yGd91bn81HwS7YfoxrvoAC2+XpAia/orLO1+WrlKK
DMpYnmtHEzV1LyzuUwW8WuFWAPp1zvjhvTO5qZ6nFsxj3FUajXUOGDneHbOv4MHx5nzeqTDFN8nZ
xW7uQN1IhqPZK4973x76IhIX0ZEVWYNpEdpPPb2/+D8iVQCW/XxZiNspDxcqy7m46cpVaIL93YfH
TQ7XhN/B+xyf5SFw4943GUH9GidWDLBvZOJp4q7IeYU5NaUNwLjfTDmFuA5pwgUp47jw5puGwJZM
J7VIWROGsP7xkb6mw/plHnVKdGhg9gnEDcgI0B7gjJugcgmjp8fFSzW+fWyPM6YUDZJf6UzSFBk+
t444YEAWkEG76OBtU4jGb8Skn/o1YvHrbc8hqpwTjkkndmw/jURGWQW0jCrHx5ofRFWfH6X798Hc
LsFquZBykF58EIjI27EuI+AycoTFmQoh/lHFgmzT28TZRcOfpoHBqKpqGlmmFHdEE12/Ho8nl1o4
I1oKEkpXeBMH8aZnbXcRBEYXeTcReKX71ZfXZzS/LIslS+dJBTqH4NBkrUsjYFOHeBXDWnWKpCG5
zEE9YfaJ+Oq8edO/8fYIIkyLJIpyzb+dC8OLxxba/mfQlVVzBjm3ct6Epi9gtj3AMztIoM+qfrkt
L3Rxt3oDoyPBmnRAPhPb+V1Tj8pdlLf4HXmHO3iLSBOcilWw0jHNUebm9zKfORrA1EG7U+WaXIzi
Ctx+QS5OveEsmB5Ci3C3x932cH2I2pm2Q7l33LPShJi6Y3TIpYJE0fqfX8xVjXbY+LUMHs9Ed/3v
hhEGy690RYZnIGUosE8mMWqbU2iFjSYYcUxX1bt5y1kIg9n+xpKgRdcp8mejvg8xs0Mu0ud2mJA4
ZBgkJG/hebUcaUSBlrPfUMQfRBLqaXnWYvBw4sPvwnGBfnISkVfW0eFVSSJ2XbGVFNTZuv9xIFWT
X9USbdc1ODFT6RR0UWKABS4Fx/9y4txWs7FImbNm5btH/A+siQ0pXtaXcJXaNODMr70xi08fTdu2
2UFowIMC8OYyyB+JDeUuDI4LjekaI6n3K2TphYlOgHvzbGWNwH8JlgiR3+p2cILsX2ULaTe4hjd7
zydxk9i8yS1lkUj6UCWwDG88DgYyGbB7fGf34lvF5XgAt/0BxUDpoFs77B6OOfXVCUWhnOR4KoDt
h9TUHZcUg/XcNBRWD0DllznDc+AZ6As9cthuLnWJDjLKdNpuvq3oJQnLdIXJsB1Vn0kDHPB233st
P2go7aAMjDCfvHVFF1kxCUt1OU6TKX17jMBGD+yJ7ZziMW9OAtE5anZfQ7Ic4K8H0rK818i6Goox
70HgkX9RlsAo9ArC81sZA3sPG8xypKlicccJ59SupfDqJYvRZhNy8O/bCj0pzF9KYURF2TmO5S71
chQ+0Jq1ZrF95l635UaxiEEfmygEpVXkS2OlDxSf6LIMcTFGQIQSJazgeiWmO6LZiIjy5Xy4q8Zz
j57DK8lPPa0/8b3Xyd57lsns++ta5vTHg9PeVeHTSECP1LDybxiGzbzEsLziis9eHX7d6e+weR+F
P+O7M9NTBR5bWpH57gFeaMVX4stBPYYNC9Mf0UUKzPXiOUreX/R0yBrkDbfcu5vqK/suoL58UjUS
Y0tnlaQ1HTP2ywiQrNhpx/J2Zm7hjwFZSO+kuRfSCc8X1UeIcKVMogrF6Iwe962M+9BwOUG1fDsU
TMyXaTiKcq5fHzekBxJxbqLw8wC0w08K8v888wY4i4t1FBwcM1fCGPSSAwXAD9rbpkXX47vcpUBJ
UFtBaHQXYS2GngqdKSCA4xhTukq7YodaXFTU4wDPySuAuM2/vqO08xLW/bEPmr5m8uflmjIVydAK
eUFI+ro9dMGYbUZlm8qP6wESfngDhhKe6KWrYXli5DxwCu8YwfhSzHr/AMMikXNzA1kpf/vEeWur
wniABOlZkYBGipgMfWFOVoKEIrElLvN+bWSZr+/oBJZUGvE0ZeYst19IqDLSuqx6XrmHKefC645a
ohp1IznyXapGJALnjJBOpoq+1JWCdtBRZlerZT3NyCQJbuJHy4s151u/ql9WT4A28cgrgAI/Ysqu
lxPnbH8zdUiw8AzCXypJ2u390fG3/vnCdn0GsTafchzk5GXm2Po01TM8iypJ7fi5ZbgfUnaAJSzS
kxDYtXhTrY5P09iMLTg9ccNfh+UyJtiQcU2Ff3qHyoVoQRDqJAdYEbcQEdeNSGsg6Xawwk4un0Fh
kA2PVRMcdOhTaOVY5PQwIfIKn0al5a6m4hKTJuj30T2hg/EengGs5VRZILE5mE3Ao6Oe4ym2sh5U
o/47mRETT3UHh9sUZnTh350FUYLarov4Y6XZDVgbYBmGyI1haP35QIC5v1VtKCwIApKyjud6TYAJ
0NujUL2f0YKrcSBaSueEJqGOPHUbxRkFbXsx9K+A1JB8VWMwgEESGGBE+QWjTuEFTFrGKd3Q4H+U
R3zFpQOQJustYItDNzFzBlyTT3VVseeKIrSXzgpvTumlO2sBzd0JafGdhlfVvqVfsuRDwnPTG64r
dHbi2JaSLEifBNbefNQ/fJrlwVqsy/WK+KOF91P6zxJeMTSgh5HATPy7dk4BSGSt433eSmVNcy8L
lIWDxh0e/D06nsP70Dn4V/08ZtMnerpwpkyAPhX2BB0k3S14mivjpmbs4PLBGP6cu9vGPzRTNSK/
xVdzPghhW1EvK2DS0G2Eg4PS25vueeeQZDj38/k8IsrntI5ZxvQY/SkMtH0MUUyiI9LyvpEdhiy6
eEsUwXQ3h6doY7LCKVchAi6oy2KHW4nawV4cJR+c6AaMHPsKV0LCc5HwJjmIGQxsuYffAJGmMwt5
Q3hgTWNO00KcRZkLstT+82FK9GldJSTZ3AawoFNQngIlyP7qVjF5bx/0H0ptU2ei1D71J4/sSfc/
LOn4Rf6fkmmlBsL+eFQdZzfE4JAoPnIpCdMUnU7LQMgpwCEXFcwB+cZH/Rc3Z4zED6Lo4aTLhuHs
7hV8DjuWXDigRtcjjFdCJMgTOW2BlBZea5MlDSI2HBx7V/Wn68JobIwthF1eZwMkyC8D8Dr612Qu
FaD5kFMKUN75QtjRK4a1CLneTtwC/Wg57o7+QnuEvJaJA/Ifee2paF7UugNsdo4QfEdWwmFg0g0P
yCf/2WTDqr0uF4TfhIC3FjS0mp3Xb7EiaaJZCWi/wyZ6r/mYLHWPjwO2SDaazJjGRR+cBEP2vjn0
ypCKb7l94cYx8RnePir0HXPW9K7y47t6MKU4SNHEeBcUSP4s308I6Eu3Kni4892ojzK1yLdo8Wpr
WruxCKvQIqX+c0tLnXoyCyV4cghSb3x25Ci0sASEPWg4Y3jzsuMVRJCgVfhXa8VtLUl84/Oo0eCY
6UHQN+YS13WUe89s+JIiK6OK8KT9mn8lYAo+BrvXhM15V3ntKTxbq2spDks90fHpu8dStram30eO
PplB21sJaEphKORHhoK2vy/c/7RDGBWRVl2uv35Aak/4ecBUhgq4b092Mz5AT9Zh98TXBVxKzlHl
ss1pV+wXzN/SmwlIa/b33tVBtn0aKy50GJFAuOmMKJVQz9+hHNldrNfBPrHcc+6bhCVwCLqtlpRZ
28Yl7ojYwbcmFVt2OH7CiAvTgLCVaU44XqkNCfMH58rfFZY3Oyx+wshHNCF0H5OmCclRCKOIcgrf
8jyRVeWmZ/4DXChkGfXcUkTmJVRK9IJR3aRhEWj1tM9hnHgk5GmUcrDMmosNMiHIIkZtWO61PeIf
hls4D1/ZbDvRgKnKpCBdcfABWj3GZhqCd7Ce/fXdlG08xCJ86J8yfNjz3SnIbmwain+0lbOX66vY
n97LoPKqCWJUc3OmDgesLZUjid843yo+k88dp3+40cOfVN//PrXYhoRxlDxDXXy6InAo87zBW0Wo
p789KQ6qDN9vNFVb0exndnGO+luq0ErIhvjjHiGofaZNTm4V76YwZCnCv42ZjD+zechbXX+XBKVU
xbhI8zF7l2rY2TINFTDK5BY7aa31SsSR4l/DC2brEbSddxwHiyYNLsfKxcyJxcJRILVYYsS39634
USx0AeqJN0R3UFXGSTUOvOJg6EPH4H0ZseJ5NghVPiulWJau1UrgjFG+7DIpOP4oS1qCny8xuGAr
EKMz038rbqkocl+z1Hg68VdOJKDmGxs9AicAjXI1KHFw118UIIQ5Hk6woxtCTFZaCyP+8YYOMh4d
eIYxQhdizbrSULz0fEfnlC8Uma78490sglTNY1Cw42sE0aWoIzTI60KC9nQ1hx++GGqY17lkppgq
m69DN+YJnGAKDepXZ3rV9ZdIa5jAgd9G/Pllx9S4aHSTY/VRqRXY18Gs0eJeGL95yDorAjnmUqZk
SD7QUNkERJLxvEPysTl9/tCPfaZHLm6UxJb/3W+PB9kSj2IwTeXBW/eBNYH9bqK0hqZ6P9oauE05
qVSHJY758VpErb73kfcDUQ12EzmNYxPIF9WFQyDUM4WIN+zNZAerKP39GVNqunUH2/Okay1hOaQn
GzKJPw+K1di17QdYiunfbdK2XJB3xtSYLSiR7DIFVy6OkR9IH67cZ7dzFO7mRp7LheQ9nAkWay6P
30EoDIe6GiWLqaZ+F1Yeq9Kbyj5GLbYLnKHkxaR/mcvW2PNI05RR5dHsY08Q/HIDi0j80RREsFRy
4V19ASIGaMM5OVwmJ13KjaR4c6LJRt72Ve/Nr47SEZG30bIdpAt8v/ln4SO8ex0kZAEAQr+0340c
Jq8jDbeTewaDEBEzy6xqBB6Zm+f0klR5DE1MxLxeLOXPNh5FEDWU+J8pfZHcHm1QKlICLYWS/T99
/tDNZNcOFx5YhULV/y8UCWo63pXj1e2GQVEeeO5iNdQEzPPOoXvrz/eJ1wfVNN7eIptJuAG2QanS
IjRtWu2B+8AZqTM51sDULIB6wT7VSk403mX7pCgibn2+VvyFT6DD9fASvJpVbAGucQ794yH81nNR
QAEqp3uWZwVvwNffza4l8+3bKnRH2oBOW4pAwoJoOoyqxtGTPrtqTYY4mIBHLYbaD8kb2hARv92M
J7yWI27VtgJiP+6BQHN/Z7ockSPhxxG9mIhfZIfEZ1rJhuS4s1m9E2nFlfONOXGCt29kkYn9BzMZ
ycV29PkITnIjMOYn8w2L7aIx9yH7koWRgWQzKRTbY37YoHmLngRoRqPuZkcNfgsCSPfgzRERnLNq
NQAzFOPrCmNqgWfnQFcgW6rsHlFFzc2l7ng17mEt0Rsoau+tmTCm3bQ/H/MLVbpTOgZJDs0St/hy
v/osyk2PXETS2ejo5ufBMTtJQwdI14VY8+UGPgnrLl2HwyYYmOqgMQy2A1vhMVmZ0M8su+IpaGwh
ETmJ4v/5zELZw+UdSVAvDxrrO3tic4VQenRxTEZAF78V9B4ARX3pQhyaPsvG4mjPP5AG9rV4JdmT
mSEHQfS+/q210J/vnn88lJt2EzvTyGVgGVb8gJdyG3OMh1PIwSeboMxzYSObt4i9/F660KybJdUK
rz0AsLQTbpzHmy1eYkhMJkl+cXyYCP0Cbfo4yQsNuAs1nTotFSQmkRfbUCavKEIOyBIUitJXza1v
xYJ1M7BVEQ8fze6Yxbz28BBpOYoMKvw/Avl1AfAOnMXIiwwr5KROwGDcbYRTiMzUubvEfbkeZE0L
VcN1l7DnfNX1NhhYHFjhkvnvTMStF1jFktsYVplVghBtJVNaUyrQ4kvQvJzyc8HbHqrKE86fu5Xu
4kx7s8clcsc7KV6XmaF9ctzsIIwX7jsytXuTojFIw2bLmuebQ9z5ssZfXE+dUzV+ICtAEyJHM6Hb
1eH4MQCPaE+nyipFHUDcJqA289/sx4fA1w0aytLGkkeoOwUqLnNZLG43cCkYcsRMP4oMJJvEsUTv
mGfKrOCXAr9awcepsq7FwzucSIW6tW+KovFK3d7ptI84n331140zPSWjrx/Jg3UPS3/aQjwwLiPV
1MeNv2hHvHb1y8oc0uHA6loFD9hV8zFsnc9ascSPM/iVTp/5qVEAOfukpAGu+r51Fn+7OgB37XC5
KoQNONQdxwBqW0OX+HAPlPud7cSrXvQr/fxUQO2LVwhY0ceRkhkWPCYyNFRBF4Kr5yxqll34hqXN
kc55cYMGd7m0HPxf3kS0TBHn6TlCjzdQQ+/cPXuT+uMOJqWf1U05kkfmbnqWv5LpdV5HgzwIVYiQ
qU5AmBA5t1K1386bflvEyKnAG6EChbQ9BK16wJOLu0G75WNY8cItRlYoRs+U6CChZ2YcW3avh8BO
Jiw120aFXSZSHH8zomVshJefuN/RRUAcCe4frigrbzIdnL+DFHQk5xYE28/mYt4G283bTjxFmFIK
gwvd8oj+4Gdl/Lw5Sf7dviyonIZfN0e5UqwnPpZ9ckn9tbR5PaAB/7GsOlCKZR6Rb6E9dFna/WCd
KsIHgAGRv68JhhOeXJeWKg5QcbDKHk+FUS6GEZhD0a2C/CjmnREfBcIkeGNkcRcN4/cVesp+ErE6
D5mrT8bb8HzlI4QYF293uxdDdcaTYDcBRNyfBAovUu/s1RjOsMPkt88KlG/mVazAQEUl8wUDqPUX
XT8wKTNWzTNTQ93UWz75oFBZ0fFAdN+fPXqLlYr0eB+2QlhSJ+sh4+J0vH6njrxhcpOXYPfC68Ct
9jrrNz0aRyB+rtnTMyw0LH1JEfrYNhjcGFKUTnyI5kD88C6McRSJVl0TkwOLVUaKi57tq1KeT+2a
zzeGnRPZmT5Db3juLtepnyZLCurSfLKjGX6IZKAlSYN3ij+HrN4qkzNVuFJdwueK5xZRXbHd/Wpy
THtS5FPMP/uIeWiMoYWVQSDTPFEdHZTQVC1G5en6BRnu3JRrB8pPbegTAmSEFD4NA8dfd9iMjM+a
x9tIHuSpDqggg0nrk3hO4Iv4EqoRgRioTqEaNWHs4xEPZdwz5FTBbxPvpHtQjhr3c6W7cBVqmphS
kMaREcZQj5JDRFP+wA1nHVja5WR70XgIbPxAlYFyXLhdUtN5nIQCSbEBNS1BxD4yb5b/u339sCCh
abYeluQpUHBkb0hCXwAYs78R/hg81Q7Ga/+mAUTPdt58enuxZ+dJ0E32lZ3jDVRfqCCF8eoWuQo+
LfUcdaifhoWMoRcZcJFKJ5HhzOZRoN5ssb7iD9b/81Gz2ndacVgL1PHVow4vIoyYC8Cm1ZTbUaB9
f6hNtc3cnGaCYLJV+fptYP/BQ1HLBMoHIB4SLyt532Ri3YD0kfqRqQhMHRs/RjucJ7sri8Is0+6n
rJlv81cAXDfi232YbnJL8NxZ/Zhb6hXCLWDEgTJSQH5qaodjXzfTLtDGqd9swM5mFbZgLBObTkdy
DWRjeh1tDnCVBxQdyVYDLls4aIlFpqg+4ch2GSoZ+qBFpHtrPUhqQPcfvpm6EDejRoNSMBZtuszR
2iav4kAkRvlHHRcM2fJUpvUhwWkfFD9rieQmPRWC9ZZteJJyoI7iYLytwj4s7/nqmmicDPmcj4iv
OqkeEUE0pQvBG3Lsqe8YsTiXM1icIn6Glkz611PzDoLwbHj2so5aae+3G+9/kdUE4Qw90ornUPXM
h94mTqF/bR0drqy0RHOgBoR3kdHEEu6w5ITG1H/8C8wow58LZBNMKpcXbLQlszw0v2D7mKUB1twJ
gVkjdocTIkQa01SGtEng52vfLUx6wuPNwNZ6Y59wRgxHAF24/Lr+P1m+qDYr6TxIKvnJe1yE3CY1
hFhvzYb/BIjTUW8dpLBwcivnCtRe0+h25QJ8+B97RjiEyICxyD4SOUmfyXMLIZmzZBncn2opz0JV
qauOHmwyYGKt9MfaVFg2Ie4Wj8OaVzJIxvugPLthFv9FCRPbBOlOzirYYt7i2GCqHh1ylM1m1h2Z
BzAMC0y96r7o9LlAGfhmjQdlYP8k997/bJGf+ZUXlNU550mP7CU84hpBVrZTnH3XOjPLMucwv9nU
YUX6BkN3mSS+Qi3DcGJUsTMaJgdk7ZA/4jQxmYMflwpMY9Q8PrOoVuNp1H56xaM1Ir8zgCP9dSqP
zdSTLRfdPAvA/rF3xR5hNs+Y/reqYTaVgLriQjUTbXQlP4lCvvTUSIJtsFBAmuLFg/kGLag5jGCS
BuqOkQrhkRckg4MxHZssJrasmouu9ZZfXTvgppxrL3BViAaganLaM6DJsMSLA781+Z+6AwKUmQjQ
D+OFXG8dwDgIwyXg2v+VgdN8GMu/xz8Ka4HTwReq4LVqqq6ufEIuYn0GxCHWlIres5hP1uvIJGB7
VFTIBlIGjpUpXWId5Dj4RrL1b/DOxRTUfTxJ/d9QhS5OcZ7XYoeCUSIxTAxkXfkkiZrGPjdaQoGe
otJ0f2f3E/wGDr+Zp5CgGKZWMjxjKR19v3FH9HshtmUhHIEGd8fFI0zLkQ6nEn4bUr43at0RFchj
2q1two59Q6ybvHyIZZ4skNNjcTihpCu/lzLjoj+rFLiCdd6b2Ds1xoYNVmA+eIjqLlLzaNLOU2tM
7HwsdBpUkw1GDGQVTWQDD5twZZeFgXDASkdrUmEJesLhxN+0MxBR0AqTqn+Bqr8K5HdyIQ7c6bDN
aWg50ZqMw/j6cbrcuyuUsI8weru8UugRBkS9R6urYOjUa4gJ4bW+9k83XRdZP4Tw8+EsHtU8GD/l
3210nmWPyUTDS2JAMxtHeP241D7XfleYZd6CO0t5Z8zHwLNKNpTu5p8280Tb9cJc0RagOAkbu4SB
lnsYVPiSEvgpgCFBdmtbcCiOdhfsQ1w8VLC5DpADdHAAmmULcqlpUfx2QUblhLgUEpOGjuCJAc3a
2TOkntHCWdm9IkfxvBEcmoJxqQswJ0gAyZLeCmIMjZ/8AXBss2OWUYQ0515g5PYvFI7MbIBY5pHZ
2NcCwbe5h9q2/H6tHopD5RSdELHg9+iSrfC4zmnQoySRkZ6BSHqor2X+qGcVmaCkCl9QK3HFz5C6
GA5yuSbaTL7tRZI7aQ9eVSZux0Ln9EMJOVm+uVLivlfRjRAh3x66r0e6SCQt2AsMnt30DN8lcn75
NdbrempTfxFiqDcGlroB+lcA5LYttE6fF0Mjgzr2tfMwMV0E+aLNxuoEk5TCjGMelmPJuvYWhF4/
z5atGvPgXj/+/6llCRPKQFreZqaG/MatiVoySd/2BnGvFysLemDedd45bJYrMYt1XLR9GizHE/KA
YgPDZzxGHYrGzlWaImqUVJhA9acAKQRg+f4+0muBpXaxabDRggx3oYG4YF3lhrQtjiZYdXUKOQyR
lUoT8fZKXvW7dvudm+N48NWXY8fMTl5pUUbKE6xVG7maUSWrpZL+ysKzQsWDe67Upd27aXYkXns7
3v54Nd/WhhPJg04d5KMSWLI3/F049TriSgiMaVlwFhLASyR62B+7OL4k90HOPPEE0uG5/MxZCBSY
SoM5BocUltTIAE++0HykVl1kvq3uh8SMW6qR9L5EUj+fpIxgJKM6l3jXJSwC2sB5iPvrGoYjU7fq
G65FgKk+/H91xaBm351OK/IZjuhB0s/lGESrl7cJR10lb3tsvgO8cH+p5C66s2Ao2CDoYOGkiJW5
U48jLtkjG5INmdleCcf7B9H+yTlOhFy8VcffTFih/bvOUnzMMcA3n9rtpKxWyyp+ehbVlcrNUGLA
Yz4VUl2yPb1OdMQZ51yoL014X+tCgs3vqqpmuXuPf7eKktemWZbWFbaszQszDUiltyBL/1vNbmmG
dXTXQH4DcXnUzLgXzGtXHj/f8d5YATO0glCBWob0uOFrKIIhWM4S+g1/gDbvXsndNuaNBnR5mHGL
JIRrQDXCw2L8gVSCbyyr7bBcnPdHoZws57rWs1/bE93P9P/z0O4BI3KsDL54Z227tOY0pkFVvglj
vpd54wFhJT3nG1WUf9tk7oM0MQIWlFSA/cfFD9AwuvAPUAKosmWEbxLq5oyhN7z6H00UPKNkmvtL
Kjl50Zq8lMj8DFZ0INiLkPZ5Qbz/jxkzVo7eAF91wLN6XobVYQKxVrXu4Kv+r4L2Ha2lL1Hs1b9P
hxFxNkjCNVF45Erj69zF++ef/yrwEvbSqR3N+qduUAW36ud1FUZ08Lkm+qk20EYbSsgtW3bZUo1S
ZdjtIWaybnHyQPIZ5JjfNAEz6K37nWOUy4dyoKnG12b7vBNFjl2i3Ad8yWrZGkuMwQki0FklD2S7
Y/TlieCUHufmJKdb+j1OD960llYZDMVYVB+Qq6DjJ/XlEhd6A8cwn33JQT69xHNEC3V5Y/5WOvAN
ZKYS/ge+OBK5WyhqPqkVltyMjpzdiaHlzsthalsLwYtPCd7Qtij4m1fAjzS9Dk/Rlif006zNzjSB
lfd+yDCC5YFvO1PzRKlzrACDdGsAsbSInkDorHlznnNarypUKuBl9P1oC8XLKCmbODtEsgp9325l
UsNMrz45ZUicUnuEuY1WAB4tjb/kEQNGviNkcNgN2zfROLdUCXItgigzipT7TrvXV29tVQ2TtqNK
LcUPlLh1UW6khcdaKqMuqDdozu4h2s/x8zqgiZsTByRhSU7bCx7nLdRgr3ZCt5OAblgrWnLjmhi0
HgfAcVZyqGgaSbgUJW8ust8x9aCwPFus8+OeRzlM89iq1KQEZrwwcQ4sUD5xZDF5XXaZvj7VnEY1
REr3DLy9TMJwGtKs9//nq28Cay/3Y/vFyOMdh3/qWxTXVQV3uId5UXGuWF9nxt2XkCJzKA0qPf5n
soejgg2rfL8xLVfOrSw6F3vKf2K7viaAHDFqm25oCecELd+ClIegEY/5LNaxOR+30GK/TpiTE0aF
cW4h91S0DCKuIyRgUk6mWv1fA7rOF668bU5iMm7whi08v8ODvWTgkQk1yPVlRnPb71pS3ixrfy5Q
bmpN7iBw3NnLbXt7O/9ZLAvHeCL6UbtIOgmBH/00OX80SOSi8UzouAt4M5oV5/BTZ648i0p4v2XC
zJMUUj/4XeTYKU+xv7yNvufWFy0XYUpcWlXvhrl0YYLNyiXQufkIAd/RrRXq1dLkGwctDcJ7wAdk
swoMZbgh2bJ8P3tR7dRzptT6ihpf0t0Z2llTHr1LTj0bxpF2pjP4xsa15LmKtW04o5yd78VQgfW8
4VKQz5NCztU2uESBZu6b6obvFJBaLfwcajGyIsa/ey4w0hr7vO/pQZp6cmNJ51vmqpGuqi+VG0c9
j72i7xX9gdzNO+JeMuwlvwWUIMTuUHNI3jXFaDg+4edh8XEe6K1x2hDu+Hb9dP29arQ6rhhtGNmU
EbsoFdGODfSixyda2Au/baOHxFKZzIVJOP2J8W0tCsvtVU/6T9cB/81rqxrLOiBI3oAuF2Fu+g6X
ERvDF7/JFW9id54Dg82YKqrM3sIdrRWb1iMyG3NSy40wlt2Xs7M5J7FH2yPWoTa2WHqZBMObZwxk
nr1e2oh1jiIsbc/gLyxZTczoG9m2mlGi1Zv9B5tAh34ApcC/Wa7IpLmzzLJceEkxK7VICd9V1pV0
GiGraHUjBxmZkoDwnmWJTqiKzKaWIT6PqrT1iST9P0JPQ49pvPJRf61EyNnjJEiK7TvwcDa45Z35
+4CLXW1AR8qFHMzM7ZVTIuxnpobvuu/wHyAZlfiR+uQXwsX9u3PgOMhZoUEXl1bWzKfMIhUyyV8t
K1teuDqt7NxFrBxkRIbFZwN0ql1UnYPVuaMzq76T9YDoqrKEAZ+ow3vwkbXzMCeGnfU9SgRwKJYv
GAnvJUnYes74+o+OxO7LTHFUuwmPiQgMv9mX/OdPvzV4+alSOsuMvqud4LVMocxUU3vlLsR65cVW
BczY7mzPN2Yf8rNOtae8JYGr7n/QQJgGGkUNIIFU1vNSu4/rUnk61YaiXp+LN+TA+Ciz1AU04+ef
aNPfhF61gGXFTzLRvk5WrhG/gCYlE3nl/NZUaAhdyIxHJM2MzhJCe0TPcVlEODA7Pvwz20O5SfIV
JuWBiDcnlp9Vj8VopH2bET5UyjGJnVpgccE4jlvnA40g+KhGswsLOSqV2AYoZyIkP+7e0DKlQx+8
QX+EJUOxNbLkKsXIYD90lQEm4IMEU8P9cfOEfGoiQ3undqrj/9tFTJt/Kf86nVjlknU0pZz1m+SX
hTEzqpASQWn9e+yOw1pUTeWwXfvmM+KcGMTum8S3eKUjx7ghfaSuvNgK6u/D/J5mzVtMzVqp0sge
Ch6yAsyBQolIvloSvX2+QqoyN8jcYO3Jtsvg0GyWM8MCB6cG0qYHHeUsbKbQ4PKWh2m/L1y/FDSq
n2BWiQvqazousZWQj0uen4Z2Ln2fogGXdOWp+ELkkzc2mOmSS8ZjYHoFETth8AlrlQNlYC3QbK4q
5wc/9FwlC2L2RT/fVOpA0FWzQP9Fty56L1OYVLjUCKoFJZafIF8391dQMYCfNG2SURHdpTVqwFTH
QmC0qIhk2zp0RUQUBy2TIt7PDzgp3qhE9t0ZeBdDOK7xbt/vlBpBgQHc083XtV+lR1n4RMxcGLjf
iIpDOGtp//fbL6srllOIBxzdS6QFxT+78Ry9jbADcB8evVEy5bWbT/CB3E4FhHFrjhHdHTqAtC/h
/Og/2aAwFZ3jeMh901lllej5thDZ7r73+c+NSM6I3pLK8jMeuHxixcHrCNHZlMMvc5jij5xw9E8B
Tehbi2qb/nGidKFdxe9yvaFKPdxMEIFQBCczBRhKBLusVdglox3cqWCnNnb+jGHc+1vwt3IFMuLv
YRvRV+HU4xmsISPSAJc/w/bjU2TA3AHJSeSZT8U/l3RFYUccZkIIkLnUZU4BWzD6HHlAnW+L2F5G
Vfl0D9ek5yK8tWll9S0wOSxbLTaURlu0206ugr4AimaqTo0fsDziRpbrO9useF9vT/sfA9lirHaX
4z8NOr550bqOMqM5uWuV+2g+Wmpk/hLjDSUmP5ElNn4tH3A6FWxVUKfXsJGgRu/ih26o/6BDCvW1
kbS61s0ZRJGnyWIN4mnhDSZkmA7jbvrMf/wSoOw9tzWJ1dy+3zbYJUKxdDl2Yxu58ZWeG+ymsDEV
lLE0XYAPZD1F9gY6yVeT4FrcxPBrY6SYHvDodd8WE9yLbNY8HRSbbLsprYPS17jp3WieJ+8+G+u5
Ov6/WUASxINxIJsyOBY6SucjidYaDepX2qkOf8lLGmSfuIA1DLPrGCX1A7oBrtHyKYEaYCQX5L8k
4OZ1f8x5BEr6IDO+HDvX3oLs59C9EMFL0guinK0xDzcycpIUFQYoTm6hmzSKPnMGUQeyEdasULIZ
ftHZEnPFtopYJgXlQ2G4capg+6znpORYN5qtFHng7dUuODk1zxhbQr+TSyc0wdGsX6tUWH/jk0C5
a7PfwFVDVS0NolOzKjsmKdQKL8D1aSDUG3iLiC2BpzkNNehApwJAq7HKeOsSF2G5SuAmtzMNOLUV
RtBwJZaCx8gQWRkcjrHD4xFE/P3v/c+0u3QFwwz6Ti8fUrjvj4+bt0TSY48IKlitxfNgpeisGFG/
khbWhHxVjWfk9+HRnWWcTDYkXOlMTw3HmWMlk/xNlo9Qk+0imBrnnWYcwptk1bmuOKyhrBuWg1qZ
ABUn2iFEgTNW5tjFRp+kdtWixGmTPfvciQwQlCB74bjy0HKC1ckPfa8u57JCk4QfepLRdkPMp8AR
B8oAu0LURjLBf1A76Bnofaq7PbXrroYpA0lmnVNQ4EgQFuM3WoBA5WA1Z5wg0Jvixgpck+JUmX1T
qoYqU5sSgqQf4p4PxThqLPGEJNTTSyxzbMmUja+fp632anjC2PUu84qrwwtlY/SIYsrQfWh+ilMg
2y5415IVlWvXASN7s2LhfQdkKqL+pWKlE9UjrnNTybw21OZsZ1ZY1QWZ/ntPbxcviYaXumt5Gmz3
WxkPJvQDMho5Xen97DI7irtfcorNXEkFPZygls+N4fRMhyadIXUGBNxYodlLJwseuL/d5cVla6ME
Y7lQ90GhCL33btzSSHmRE+myDmvI88zjP7LY7z+p4vLqXYOgFa4iCrc3ijItqQzKLfmQdiu1S+id
yyo5fAlMYGebBjKkaMDdWkUEjxG1NzcmuoXvipnDyLi8HgmiE07KIZ0oMxp6bnXZceViMRCBvs4V
jW2Yp/6RtMLy9leEIHs1Nzogs0Z9lC1UZm/tTkyvxqU7B5Pya14EbLaojk/KRlH0nmxmVtD7RUGu
4/EvojEmz8ReYUMYKYuyHFV+b0ON7j9hkO3sRr4Z6b1zJlZddDZ6NRJmXvOo/5S/K8WSwcJydhaW
rakSeuFUa+awHWyVRbEWGDB7W22lqg6nw4yGOZ8VC3vppOCezvdjbuDFHrkh6U+7Q4wLUFdDVW4v
UGtzOw8GOTjtHW9o7kBN0gMEQpXb3UODcu7p5L6RyIIZZVndS4+NcZPXLni87N/+yjjEQ9zB0Ur4
hI7fG+iETk6GmpD5eVZx2NO0LHzwnJ4zdUwEhs26XsRbAmBy38a51A6EkGvQT7UMSDpS8qUiWx/k
i394o8KJD7vmI8zTJskEr1uaBlQhbOC/9FdXLQVbf+JirqaeqDaU9tjBROSbOLg8YZOTT2/jP9qv
MEqaVaItw6P2cNHjvdghlWAlmIMy1RquEcQbDAB1U+aL4+YbELJJTev3BzY3W9JxD0nAqlEc2FD9
qhlkxwDZr28Y5FlRsfLciZmauSCWQsKVvquWHvHhvzFc7m4B/hER26GjUkeTVtEPmNh1cftQckrY
rLKw/TGQJNNndJb2HL5kr1QB3VPs97vHoxOtfX6tMYW/a+YLe3R+0sdN0wpOBxrOGXzlU0ibVWHr
C6zUYu4PUYpJiVSScRYaF3QXPrrSwY9MKOZkXZMCMcLOKNKd9wZ+R8H0vFgFH6bhy68EYhIPJviL
5B5G5FRQKXRZjRXEMkggySx2crohH7eVVyY3XV3FaQNbaYIVZE0BDY+Zscqstdu6tqe4FE3tZwob
dWUPOauzBAIM/PFKWniKSOM8eOyoTBjU+PyC5OBE7RznVKOJIRWXsnZESxjWGkBX74/JqxZGDWY6
uRHhp04BhCsDuYkzGU+Kkx+HOpa+NT5UpLKtn0uz5qdJXEK6YlSqDH2f9UkxmjvkBCiAFouukmiG
ApuvJdjaAy8gmNT+K4YhvqI1v5QSQ/7vakw0t4h0H9OZYhmPOEsDWICGxlq228O8XjfxK6WuRFEG
WfNyqAaGr9tp5pn827/ociff4MX7CvfsUSUCtfMIg1OdXRlqqGB+BfuAXY/2/rM3D3M/9wTKTSFE
X7524e4wfbDcFDfErk7L5cqkblcLSvhqA99ippIlzmJeJFgiTJ8MROGNbNXuYkqimtehuhcGSyVj
I+hl/0uOvxFuWplqVYcwoWGeVdDYEKO2WFKYbY4tvJomk5m1/8aBEMpeeom7FIKV2fVBiCUbdTam
JqFZVQ9VKlzJJkNnSWgyhcqNFD+Jl/I7aH2cqBpKQzCjkPfXrFVeg72Zeel24b77RqFEVnHsVrBk
5I3P8fxF5OTfhXegEoEWaPutwwu5C9H0Uc0S8DjW3CS1zD7fV3G0v6c7PVI2oUOsOVwW6QRRksfo
/J74JPZ9WBf8upA+K5QYYe9mgV9XNKs48i7XIa5whUQYfOm0FuDzajZ5LxWR7vfSenhRn0lEbZcJ
s1uW06d0A92igpfQGA1DpoN1Xxwx0mh1Su7Ann2IEI1nVeQvPMBTwq0zvsB4eDc9r3eskSzcqHVu
UIiXFrayAIRcvDkIFdqJibM4irLZ+QsyHzojkaKhVF+n9MPA77vFiT85neIoYcInJ+zPYv2T2RVP
5k8xIg8L/ptoNG/kLzsPlC+FPK2qA1WGGKBFgnBW10DhMdoOR9x8fZxcAxkBRH1infQzSRsDXZvd
Wwls7gd1giTIetb5QP6DSGabuHXv/Mv3vuUbyFNpoHM8aT2XZ2eVjQixsYXmLRHY8gXyWjjCWCRD
5W6CwqzwZNufB1+hEPQBTwWeaQEgjxKy2Xa27/t8OYl2Dq5WOnoGpVbwb7FedW9gSGZcxTPLGdtO
L+I+sb5ZaBbQRuIFdEpnVQqXnkAOL6Jrfxx4pwxMoKYo/NVvPhwrzkb7euty+t/WdK2lXBbrz969
scwQzK2FVCGULDUp7bW6NAAF0t6W4UuMWoeA7+bpHg02z5mB/uS80Q/NqGGdk4AmxXnXm83DZAuB
D075+F8SU30XF16KzrxRPqFI/AWb62VB+qMP9yp1v91P3h//pVdpYI82TeXiktX6CKg+AVsYuIAC
M0f+PgHltu4deSqsl0LRZ/5iAS+u41C/4pk1k4p77cHuz3TosUFAUDZmn1IeTATsEbXZfncfZmLZ
BvDTJoPnjgypAAMK2sqaviXiMIyDChHZDD/DSzloC8b5NidcGxktzl58N6daCwjnwKw1CU7WPBMz
Nrn66V9owGMudI3GQ0bBvlnWEGDT3ne0Tjn60hATT7nj2F/RjMpJW5fXCr+tYQb8AdkRA/onskir
4DD3DH9SoZB7NKkTVWXmJBDZheBJzKVho18KaWdb6tZvNEDLFe5L6hfHCnKgY/MWmJoG/uTZ3Iid
jD2NJAcWesHfC2tZGMF6QcAqjmO7lyJquHbSWauzw5Hr4KAy6yG/8dpt+1UUKxMRe3Mq+fZigKpH
RF1/WoCzQD6vSf2ZgfwF7zGXgizLVzZgzU5SAsVr5OUbpLZ9MqJ5nd+P2GdNiXMFlBBj/a4z1iTe
Bf/qUK0LgFsM6IQJuiKAmRXzYbq5GNU1xVRRR4AvD29vB5rtXdSof+JJ+QqwG9WSbGfONA+JTaUU
3F/oW0UwKneF/XivGnkpAOYvsIXDo2qi63IiLOrajJNKKc58xa/e/NqpTLa/8Q8xLjgdzf0l/WDQ
5EwlsII2caHb6JFilQbOHYvNqAvl3ahg8c3tZuENIitUuEBqsx/4stiCL/nxkxSFpVNtHEatYSWZ
rRaTBjGk+0AO0g7/x/OgPnU5wmnKCaL0zYoBHbX1/cnf2l2ZOnozgUmFFFg8hUGoAnjNZpZFpuvW
KdnZo/WB+vByc45Azt2vlWUiaLWp5oNMQyFb3GlAXAxi8/ngM7f9B+5+FQjx0MsxhNNdaPYcDLjN
Y/76AkSoEsxuAf00pX3HCLw7l/wMsnPNStQHSLyFbSJtVxOd9yhHqiTP4Vx+9YJScpIutYpiaZpM
OzybGI2dFEiis2VoBYM/pfRhPrYQyeCqYV8TBSucua64JcrbvuflNV19/dFMEWQ0MsBpuai5JFC0
+j1tTNFb7g4wfM6JX3fYF8mrMkM6DTybppg/HDyuEUWdyrA1thID/lTEpms0Eu3wRoyCJalYZj+d
KutM0mhDZeUgACrEI7kkcHq0XTDhPimnOWkQK+L5/ue2HSUrgnU8+W0jmI2v4f9NnXaavkC+3n0e
jPfzD868tah7hJrCitY4rsoWJH4n+wy5MJCbyeE/0PrKvW6tln59pjHshDyvgZJCJ57KWDWEW2pk
ZT8x2qQh3Gb7kpBXj4q9nrYgo6DuwtO8fGk7Xrtofna3Wc4bkH5L+56dhnW93ZidENJpm9tcqH7X
0/w7Ve+Q64Hot90oLMgqv8phBAEbSXP6nQ5k83MdVuKvEw5k3SjXBvZsYATe32Jj1U2zHl/tnzyS
c1D3eD+23LcYvyZr0Q5MdheswG5R30x3ccq9Bs2VRiFedGgMppaIyYicnnPK312Ykwqz/U4wcQsS
FBtJErtLbOtkjtjkV4wUdXBmAJtgY5AcV5kdUSHch1OanivMx3tO/N97G72SsOkOMIiO39IE+hNU
/ln1FT2OJqN5yfrJdZ5xw/EBzAh2CBELzqOUzFh9n+u9ZhIDiMzPHuN6r/UliBCiPCOmtebrCY+U
N4PaqPeqzGWtp70desWloWXcEp+/REOgPlIHjK4c90KqqJhqlGFcB+vmv/4W/zLab2ed4OeDx3FM
ljNyTczDRK9gOcLyTbh1M+kMKBILomiY1rN7JiUneZn95dd0inmCtsJo3JpN8E27+ektwjpfceMf
nVQvEFOO7KwRXN0tKQ0kYuZfUt0ycROKqpyYzZ6yD5ebMUFTADtRSgQA3zHDLynWD7LEVIaKSpaw
xlsrRAEG1Ysz+Ev5Wp48fIxivM4KMplTF8cbZtJlujusohxbbOak0TBw7Mf+caDHRskV4o29PjJX
59CKkJkSKGhjGzm9bwRutAefRu5IxQy//pdCeT+YHZS9Phyd2Vqtf3zhVzJGZDjwJfhWsKMFyvxt
/ebw5pBiPyL4M09a/fOYQ1RYK1SSu4Ipjct36zdxjeBqykECMmcboQEqHEdJ2OX4/ihby4LqvJqp
IrWEjU3Mwo7qua1MFkZSoSS4v/G7aVXUgPQ3xF5/Zp6UVzWe5aMzhZeLORRD+Buoxi08tqzkZ591
Pwm58AefonvkKh7ECTcS9TYylZLHVYkDJR4AQIptNgszWnGWZPXjcVUHCHbHXcLHHJSTPLsWP01v
yIWn92zSH8qIsvJLbNMf3wbu8L4bL0ArQvMijEh+KceKYiMpiZCZCXwC75daIzvydCoYoKo7Nf5H
dnOx2QrFx3z09kpYXHiyDwwT8mEeZy2Y6eQCOZdCDpj87QR9s0WglwSLCJjMaK0zgNKw/gBQ1jmg
yH+ixSUYCGH3vTnl5GfddBHN7s18zbb278rNycq2I1XkH2ByDB6cNUjYFFJa4gO2yD4tx1hGdw0r
ReJqFnbu2/mdYwJHHvdV+F6enkpx8FDctE/xRyTWdaCQWTa8I0TiT5z4i3qXclg/zBqXsc/pGhOs
NXWFaDKoW3IK5zLAEbyq5VSA7ZXtM+EAJrUpiw+RIxSpfEwY4tkBgujINorEm6jZWjmVEOzk1opY
4JRhgDGx59x+tnZ8gv2DNg6nsEED6abZ7ERa8NBV18SGLKucWFFg2bINopB32Uq74jY8dRawUNoR
CFt3HJ/qLm0sMu93fRlOgNONrRMuRtkvnTkRG4f7sVA2qVwu9lXHp3B5o2H1BifJ3KFxnFKEfOD3
Bn6xZt3Ye6hOvxjz+2CzhUmYJqcCO+e6pwUt2etdTKIjLF5OQu0xW0y3oDwSdqic8MF0eh+14M/5
nj5JyOnmyswJxqqeFSEmokcx51IWaVN9RJxI/va3l4XDJlP3sTPn4KHIgT3iptYG0vj27xodLU+D
/MeizL3SFDSYqJfc4A7s+qNwUYiH8G81rUAyVkp1GZ+Lb3drQxY+mA/XSk8IeOtNrWGKHF2/ADlv
7KDEZA0qOCPq1f8TBjjDRdHRkCbS/8iHq2seWUik1PO79iGYhXrmR391gvh3f45e1AxKddS3VC6O
446D2MwlV64fKgqoIjruosWeRvrlbjpeDgTE6xsXLKEW+gdxzCiffU2Qa1y+cSXxcirkI56M8wCw
sXAvazwfBN6tyV5CtfXGrof0zvBYCO0eEIN3OEYIAT8ETC78zjTcI0Uzaj2k36e44mZ41Ku9WpGS
nImVNmklxKk62qyFdf8NcikuICM2DpbkT2nDYJqdTfF9mm52Yww7LOpPFRyCDw3nv+jns0PXKg0y
a3jZB+C82TMd2a1EVUGtbX3VPIJmQqhwIll7jvJjkc8LeMYrnxNRbC1OZYd4krct9O70N+nbfEAp
lo7U6O0zHYnMKi6qp8BatzL/dssQLb7EsK/rrYrDYZT20Itu8Ici+FtJeTxz5Cp3TYcNo/lvsWz6
IFBdypBnlidOOQhlCA8m1uBL0D+uqlrjLekIO3kwJtan2aI5aUrS5YPeIkHeyHDKJ5rO5/+NbaHk
fgVmzt8zNP4X+lH4QfGJ1VrkA4blxTWAMfcXfBaa5EG6d8XSrH7kffTlUdsrfR3Z3ENMy3wXy/Qa
R2I7eep8ywmY2/bdb+7PoGAlCAt93IacPkJBmpoKb6sEW1XXyTjkoqAIzDWzVlIMhrt4jUy2qnIk
S1K73oAzjuE3QaF2f7w1rp+dZo8SyWA2wq8Lj5LVnZd/RTlpyHJvFZS70cqbcSocZ0H98GK2v7j/
3tsVlaqjBotKF6Zxhp3RCiK2CA2ZCILkllQvMWWMwips8fzN6nPkTS5tjrsqnjLgXthNvi7YsNlq
L9AqzWqtdNxZZtoa9VQyxJYXLLfGEFX0nURrAnoENPeteBchlKuF3/C0qCxagu1f/5rD3R2E5sg5
craPU+whruZ6FiPdAlZtw8FN9/8dGtW5/VUfJPyoEoZ65Fwh2aZmgAYK0+tolyscqslmIKXjGTO/
lGU0n39WgDiIaXAnxpegaYfC2U/OOiu4kJMozXF8AGczRjkQJZiZnaNjfp4VXv1m7usLRdsK+O4T
Bb/6WL6w31hwqIS7zUwWkaQRb+1/fkoIfCwOzkMmp7QxBgTwY1aRqKU9mdSctiTL064W8wBfsPYl
uqtB82ql4X6BPH5t9WjEOXhsL4aNYFH5BO7r+bl7MlpXT/jUx+/P/P4Aik0rD3/zRkp8yMCwYqWD
aprNhAd7JWpeeF6w0Po4j2J0kykm8Gi+KwcerZf/vQ+REGPUhAivEun9683uK7b5cnTriOEu9VCS
Ey8GuWcPW2ih+m6IJfeGoVDYui9T3ALMcX8qYdVW5pSHco5Dgr/E2Vv7xIg7bLDaJPcYTLXxI2g4
NWSS8kj+ixJHC3KiE0kTOvBQjc7j0p6VX+Nh5lKAIMulvSzWrw2PfKx3Lholae4K6NAnMErIAeJz
TCvey2YfGl2NDVYS1m2pX/7M1clTUfk48tXLyqSih6ssKk/0x4diB4o0zThGOZnfWfToblzAow5f
MQ1m2SyE/3VSozVTIuscXDkxymSJhi1wAkFr0RzSzJLKQJPyBBjLY9w+pyn7pPFemEiqICxNjVS7
H4DAVO9lG76qAqPeEzVWeJFFOHx4tpGmwyXA2BJQs909Bn9iYUbFcXyHq0xBO97fl8xxtIYEzhSd
AMudyUl0yD7wHAIQyfgIEv4BkNP18zEzVCFk79xXCG92pD1rqR8thIJHIquZBt1D9NDgKDWQ2KN4
6ShDW0a7l2OiILXBiuU5AuOiNWkLOLW9MITg52j05dBnrIGL4tzFxonUbeLkfnN6UmwEPYJoXhw0
39omykZOScdGasEipUnGcmkwVfeAKoa2UoL0picEiBGHGGjWizpvMFVzBT/B4uN6PElvhxie3xTg
Sreld0XootbHzlp+/wGXnDMY4Sjx26z9oF/uXBgW693NQjscbG7ud2UCJl6U/sdA0NmvDrDsIskL
gSBti7fBs8jy/bWUCWoRuG90B+y+NbwIiBCbFGB1yg8/wAGU15w4WfLWBfKhJe/+qdByoGpceIjB
xoh2RCBt9DfZclm8yw5BZOCj6VJOr/AR2fZvuYjsau2c/8gwF/FDLIgTrBQzjV59g35XdWbgudyA
T5byO8fhvOprJjfHDRY7HLuDkTWVXa27U4fhY1j2MZodkTRyqUvoeuZe8I/SF558pXNXTeBMybvL
wgE4EsvnFaTd6ODxbqPoayP4UzT/oI+J70xdBGvGYe5F/qYf4h3qJNZjoxNY5gesPqWQ5E71Ap/G
Ahrfi7z3SxgQLvQMVbwEVG39H4H6nZsEhJcwRw4k/+8x7g6ZHrFgmP3KnEq9mQxzBvZH2v92x2Ut
8aTDEIqEBDS0LfkgQ/DHcNf+xB/KIbExCR04u/wROJbVs4tir+OS29gVdizJtTclfZCKtLtKI4J4
JzCNUFy/Bdwl3FQ8kJ7fIKFyvO2GejdZndk5ZlFFlsZPolkmeYzFYD96/kII3JuL2RVomyk1ZW3F
5NN/a3w5jENHVEepRD1iv0uuyDEttFUz4bji5EHC+sN5nby4Vu1eJ4CixdXwd+ARxVUSWbpBTgLJ
x8PS5e2eARvV+Ry31kPQftyrnQvY4bMk8B5gZy6ryeku9qsVkNMGUi4j3QCuEEYVWsXKcbn4+eDH
337+tSiomtM27PoABAO7tP8NAyHouEt3GaPzY59Cvr01QO0BxF/367Vwv51ykabQOA10vZ8UEPaf
6iWpprsyxT8QpEvbkpyjPvoTSdoAEI2mPZamxzU0ORqd9YwBSQrnithty5KgXqsQlBg0HWWSRIwq
aM7Fu9465hIx+g2s1pndIegJUGlFTku+OCYwK8WDpGDaBz47GoHlHUCqmC07lDxhgRdrRlE6JH7p
VQBWuhRzOLS4TCXU+0w12rybYnOFsfm248smkIJElVn3PFHDCjvHditCM6S6Rb5uR7UcRnojtnFE
scJm3JjZGJ+DxktRU2Q4vkDjPX4d08W6+hSi4L3Qd3edMn5B6kNuil6SUAq1JAYcWYn+0vg9+BLI
QrBYz0VMBxJZnaMtW1pr+hgMYAss74ugUwS/ShzZVuhe8qxIup8KWJo6fGDQQsCEW6j7ctLFxdjy
oCdJfX28+4BwpKbuEl4+leLMG1Xdvb81i4lL3BI2j1xemNdqZBgNSr/2KsmBsryHnZkLklqOrvyo
15A5XNOIUYzkbjliqG65F52uKtz/TxtbzMeJPifUlmrLSuz5Ag+ioncqfF1zQMLOxSP/VQJHdG3M
JbQF9nTQ1eFp19rY6ZLmG4O43c8TcwH6J39sJ5QER0YYCYI/0VaYjiz9LPPcVulPiiI2WzYGXVXN
UZaJQx297DHDq37D7tu5kYdtgM/nYnyYN6b+TR002w6OAVJlugfTLFGZF3VJK6LZN69XvIsktUwP
u1Palho7O87XNbwQv5P0lwq91FPuREfoUekmuBLKR9dI1zQlK278bXygYnQZ+iwbl08vHsT2A309
FALQz5t2tX22HdDumK91YWvFOGql7qDT493JDRAWOxF/+AM/BaAZs5K4QLP/T0hM5GIzHsccZt//
XCSiSV1QEzxi5z82ERU8XZhTFQMOLPMuyVQCjoilwHamxxFGAM8LQslwpZJq6wCYTiWtUkSPc3eB
NyPuigVJZd0W7Uwubfp2GpVXyaUltvMqdMgMWrJJ2fEzva9JNKjLikbCXgLDAovFnnsXUjEyHwd+
9Xs/vGZXxT7Zt9ENc1moW5EJgFdnyraVC4FKxPSxtQMwdA5JdkXDBsBKo4If0FO7IGkHEMr9Z47R
aIP5We63EYtZKEV5Dnum0HfXfBr3OEnL4MxSK/4Psq4BkZy7cnzzp0o0Tb1DgyeEfQ1Wq8S/Vpcv
kIo7SBETtyyzHvse0mv7LVVYsCqgKp5PkhwwS2givrTygcyY5WTw6do/C3gjc0T5JeCndd+5gDtz
EXDY+8n2OLUd+MMvPPIzKzc7Y2y7May/zjie4Js+FacFjc38+hH+EsDDM3pPuUoCU7N1dt/ow7jd
7g/u46GiXSB4sbRkcBGVK+Ku6goUDq+kMeTiO3e2ly4dJFSuFX9VfnniRAUwvUDrUGD3diH/rXXX
ehqiYKoR0etvsxq7nVJeSWXA469l1l2mibIUOFVtKLc4PTKJwELWMBSD2570x9wlTkZZ3Lc8EJsj
0/xvJiatMTqWxf21PHYKerIi0nLGtSOMrFNa8AOgLkp4kZhAP09GJ2Rlfh9Lw8UBH7UR6FwtO8kQ
P4geTE855PAM2b7UBMMPoQdn6z5XL5vGt9/6wsLHE+h/LvA8zUvqO1lQAo96VM2VqAXTR0Ue6msY
iKpy9tSia+NhBL1XOMAyEScMqcHYMAgNwsfosrxjTcTp49LfhgN3LE7SZv44cMP7l85RnkYe9VcY
pQsa+QGsm6ysnW/5hnj3E3uQ8EwwphGQfyH4x7gOWNu9HdPTA9h6Gw/Dx25l9vaFtjnMdL8F78R9
bS1GzyInRZQ+6WTU20UKMfsk3S8Qe2Q2HDGz1PHk7j39pF3VA3wuL0ZRFt0g/ZYBgoNaG02HyAMK
/NMBGWmelSWCJ1K/tDWm7wQlYqP50ow3P4TccgHToVZNYH4DWYYYXOH/IH1mBsTx5flYawoBz3pk
LcNpxeZXRpSZq62Jhf3TTA/UQyyNw7v8c7UIzuXxIzZALbpcxAgFitv+FqUHlnqQ4RG6wJkbz/mM
HiCTz747rD6RKvmtCtwYNV0tHDDp3TBMKdLKBXglpBWdL2b0f5u2ZpowCwWidBFIvhexdKTXnxcm
I3P57jR9hKTWPjZVDM3p8OVSkrvBX5n79InQtLwDaq5qQvkYZAcjEOPYkeDR8VpvsBX1RVwoPAcF
voyZrY67svIbta7NaDmIq0B09TRfOI/dl+StlPg7wLpAej/2tv0Rej66SQ613B5IUh6+UjpKaLSJ
eWSy0GrcFhK1Krgkl8hfcevmA6tI/jTwOZT/41X4/27ZJtAZfaaK4LFT7GxM1Wr+zT4hEbsCYsAt
QmM3CVil6HLSPjf3mS8rbCNGRHRH4M69ym8HaUzWOLa9CTzuV+7BoeVYwamDeZp8rEWc15n4TjUM
BAvIkOL1PT3xvSCGufv3JS9sbdQMiY29NeEyCk+7+gQmkt5u0qWeOyiAVOQ09lK47auvNYFeSHIX
35CsDNc6bCTYQak/IY/lq4TakTCe2lagazO8iz4bZHBaogFHEL5+ZuKSonbjtq/vNLPKExXfsL2I
Es6OPeurscajvmiRtmpfRS4Mrtr2yQCGu+gbXcFWX4HRy8pFmJ4X9jFoUDOQm23ATv7OBeQAYHC1
WRD82VcMf5jyWCIh9XaoEuI3/qL/4T9u82MEHdAv0gWgbMwz/vqAr2I6o3fsFKKXUYxw8zaBviQK
yFw+G3eTNcpmkiI+vVv4mXVXW71fK575cMu3fu54HtTcRGkfQD62O+P5FXoIa9dVyJnakFZKUD9l
Qd8FrbBRLIxIkpmpuRMDGAeVPavu8Tyi2WrtvBj4kw3UnJLkO6tCDA0Iq3yHugqnNnyWThzxiYd9
tzE1R1FBOrBedfydPqcVhap6NWS+m5wh8HQ6d3KHu95AnmVwsPeICE8B7q9LvyUwbBzLd12ON/eN
joZkx+ssJtr8WPBgwIRwo2JotsUqgRV43zlslgB0dbrB3z1ZQSvLUJsrfJsiXyTYGhDzLspwByQ1
YbQZdkhJnxcZW+LTwdOLH5Qoav7n9wSiYsbsMjebembUh8Zy3DGI97NTxA0g0GbgTEGS72Wp7FdH
7U88mQ50d01jb9eamI4XrEkR6LbHIt6L/XoTEKOHsXZhulI+E5XwmRWhY/ZMPReHsDkvvj/TW9YV
QtCOjhYouxrHQwVqZyMhhrGyTsyA1D/r3RVEBmGsxterLYfaXhit5wZvJA9lBGuv42n65jbJfboh
L4P/7yEyMGy1+SgDPrBou4LDalVvbnXeEE6LFZPwZnuDcc3IB1nWG1PLCwP71ogii6wNnsE8hf+O
/flvqDUx2qTaElKroVs9ZiRaWcs9aCgLKhpsglXINlCfbAYZJZZ3h7anFvXqUbSifpTClzIMlPu2
HMJqkN/bH2+gnNTeZFX4wFSi+tRJLbpRi7edGP63AqlcGOzOH7JhSVX1SvaBfORK2lTf2UnDujXk
GxqJW5cGwUMFnUDjz+Nel/D3fZFN9G576fx0x4ExwzG0t/JpJ3m7FM2ZOX7l/6QIxIBjzZg8fHDD
o0CgcmFLSqrrIewXCIOtwdI8Rmm7U3JisIjMB1xC1I+/rfCRVjsS+W+R4HBnDqbXhIZA4VmbszpO
+bDF3Y86envF/3JuldYfbn6BHGMAt3w3Cwh10G5d6/rBKCEYSOom436rWPN+bLb5db98ezuo21j2
bpQWQTR+5ir2e/UfbejIeGGLoi5bcZLbwk9giMFHf7iaK907A2z1bEd5Xred5UfiqhjEqaaylGoV
5RC8nEaxkoz9IqtACo+U4zfLVkaSYzNYi1ShLNh/+GX9RH6cLnqQm+g2dSNSHQk+3qJpTcZ9B0Ux
UTdexVUEmWatMFNbWe/d79ugr747KbUDLKF9u8C1a1+fwagzvCFqsk7DZWSVbAGrbj2TIUzCuj30
oG2wiGlK4sGkyPvb+HduWNnnvpma7hX2X9MlrUm+5JONngCm5vfGNIwDY8vEmC/OXv2q9lUaw95O
LRwG72stS8D8cXTUwzeKy+4VN65n3j3g31uNir5J6tkXT2+53yYaiqluIGILQOR5yakqcG1fYv9m
2iR0tjKzmTXcy+WUeyibcdpEp4Iu+78ZDlVi/znKMyzlthTkYbNnThrGiVSa28+VWp9gkf3XQpNj
TnkfO41E8+aF430LGOzBOWXq/Mx0t5dycdT/nQsSqKYnEFFzYJTW2NplMU8I8rp4bxF6Bz/5W7CS
i0A/HgWKXIboaNpQJI0JlDhG8w+t3PD47QU6QTn6OKIdjzJMNaAATp065p4GasxqZWfpdZVrAjS7
+/PiVQAOrmukPtiptVmiXmiOZU53TXPtmk5oUgj4gN0caPlZsqln73u8RIAZJGhF+4FrRYefdduz
NkYVMKc9wl6lf9mxd31IZp1mIPD4MzRT/vzXmWVsnpMoiH2pe6wsVI/U8+F4rGtA0l2FBEmqEesN
F59Xt6GYD2Iir+iJem9b5CHMuTMgqJ5tPQxHFISgLTeSMKk7JKIp5sKfJsBIrJqNZXtkKyfP43Pg
C5WZLIUuX5lJTAF6l5VI+N8GDXD2xXzOMhwSg1W2cS2T7qMQ/klQY6FZkN67zmfY663qgGk+NIbM
YBDdWpJX/FVbmapXGP1hB9nOj8Yhe9UWkhFG+A7rIDMoPYEumeugny8ntHFGVYOEj1ivr8Ps6OSB
9eHtMYIBjlOEn/gsurC7SFFgD/iASMTXSczbP1HkhEVDuFkQQtxjNSJ09ILUIBE2bIgWci/YdUHo
U7AGfP38hfpJnJlZauHIZJfmap3NSOS5KYCS6pZA8q4OwcduQfnDAHAGYOZf87SG60sYvcFg1seo
hinu9/TDktfFcUg/x5iQWqjhq7qJ049O5cdi5ShckCWZLK7molEfsZWFUwunCI5mjiqUcqOyC/Z3
9rQ/ZqCqMCmqcqg+XuY/f0qgYqSI4wuoB3QmwxJbznBYBPesWZYX5LmPfDSMNKVFmWzwfeZrjlXV
O4p544kqRa+NKyC16jWsUTkjsXFv6q+oYQShlwyb+Zm8OFzqRAJHV38xbehf16egQP+7xybfpbRd
O5s+ITsgclqGWPzlGf1tbOEtbp05Iuyw4grWRUrCVKU9o/O9ym0cTW2Bom+0faCj1s09X/zhH3IC
8PkcXoB/sk0YGVvYUVoO0xdZfT4TjOeZy5jHPukZkUBe9ROVLvMqB4RgQcLRWdlNxtbQHH2HV20C
7VA95gTNQ1ocIZAU4cdJpCbq/Dy0OzfXkF2iruy08gGeDOHYNkRevXo31pHAUI/sUz5gwynMn7h9
QiELK4L6nMgW7WGYnBfq2zrnk/mhv/BHUFnKsETRyyNDjVkkSvIXxulBXTE/uk3fum7VjV897mTi
aD/zUUMptCeLAenE3XXNqA3O4W0lHcUXPlVnFJ3yWZoYhSY8/bYuh3Oilgeye/+VWrQ7Kg6ZCUrC
j4CnXHeoBEYm6LHotaJp4jv8kf3JB+MDLCUUYfmJdvYPNgpNZAmG8VJQxGjw9Xe+J5gDeag+JuNW
Evk+wro7RC6TuXPuNiJk72ham7WJ+m1pU7b1ghDmwUb85aZbnbJO3iJYl5Ki25xaEkpvZysvfP9h
BPtCPrsVKqN7/fwlmdhksFkPDQ7OMvz+DEpRLYx2aD5XSvvGmIq0OpERjGqvf/cXXEVrGAXFxxoC
BSIVuIijnL1pBNirTi4FK5APRo0qziyz2JvBO6xnpRYzspMp0Rg6ET5yuWE+d7ygYIhmRqlL++Kg
0Nxed3SHbShUaC3kqJsrMEk7jv0NROgkK2CEf8EXx7knA5Rky8tNR2igcI5Xaff/bVpIkmzEPmTH
zKgQQgGiwrRCbkx97woyatIMVdmjPsH5SMDr2A35UBN6goW6B44v+fdtN+jQ07GXriMRITVyaPRW
iR7R9+7pePokHqkR2rCyHZfjd4+nHa25vmX0I8rVPnTMCPhbJG35yzj3GsIQ9pEMMgg75eHpUMui
11tnPpKpYIKXlg78y8opUxWQxNxqoa3tuEsGK5OI9xbhnfm8TicoAU6UNJHLp5XV4bdhHixQg8a4
AarNwZEOqViDFfYWqKOSqG2V9G14KNq7FXWyIW42/MaZpWkc7tTNS5CndyZVH851/oijrFfF+17q
9lA9QmBNzM+QVcOiKVLsI2LVZcenC1VYu+54cdp7ggj+FyxEB8pi5WCWafPNUBSqhotUgjpepHi+
2Slu2ksT0xOp08lFoRsaHw+kZjKoxdE7CQE8byg+c7yKjUH/ZbJgMhL/7cJFSXAcjs7LQgQe5qxG
MP6NaNFJ8RlLZ7bnER/kmluZsaeNnUV9hFOJF6AUdgO1Oo4TWCVnF9j7c0tFxqu0oHaGWN/CID1I
gAZhlsSUNo+YKdiUUI79rg8N82PZePibOwfMyDS39cn1UA1q5HTpDL89+k7k/DCai+8TTFtijO5e
KkGE+a7OsyCA8waNXZzE1zNoK89b13RG+Jzkd8DzstNQY22QctWf4iYaQloBqPdzKXPPjCcLCD+m
+JJHBJ2adV+48/chg9bd9LiZGKy3b27xdI+ZO/e+0a44hx5POxNvEkgjloDsvmOywOAtna652r2Q
O224azyVWt34FI92FxGI1sYeSSxzk0nRm2AQKe8JZ398j8rFOZSruJR5rAoEAV3XaVsUY7J40iK0
EeG/lCtpz9VotDRMlqLm9eaubC+zcRclFzmVafKjCQUjjpywj9FAhLJmdHbetShpFKE33b/CRcKV
lV4XE4lssIllsCR8xb6g09W0wAGR2Oimsf1jzdB0cM9zQGC/14GV+qf4GVxANvQ5iRuY8Ri+HitJ
hHh4DTAwFAzO6WeZndTE1Lcg9J79gYb3I9UqIgHa0NcJ3BEobjT3/IZXvjF+qPSTgx8WZWVp3XfQ
fDPpBn7IOgFqu9g6BESADUmQ4D9evcOYCkH9mIEDWlL8Wz7mNFf8rCBEYdSUb/Ah+dKpy291jTkW
QicZIYMU86nuK9wrkHql+dkYQyBdnSwZT4oO7KtMVqcWP7e8k3VNGQTGi1mdb3iY91olLEmtMcEq
tJV8BYtk/QyXIy7AUFcTLZnj7Bf1Ftw11PPxJOmvemXqAw44gfiuBrTeMTwVoKXMHCJu+ydmF1F/
3hUFV24EcVzrzDeynFHsLWGJhgyOaF3jUFUwHzeVhhHA6JQWFsSNckpKL7lAs1PysSL22dNCzMvC
a4S1oOjktqCeZPxEZnnklX7KG68R0oHMNxnbWggzFVY9CC6FdG+E3WYbWEflRmhSqq/pZR1PRrOH
4nZaCkNwS90GaB6cioDvvLkSruLRUA0u1HlXtRyu53NJSKmb4FdF9JGjPeEJSLzx5HME+U7U0M9C
Vq0+auOsEu5XGaMQ56IpFTjA5dSMGnd1Vo1By/7UIB6D4DfcSwTJGnwVWqzFanhL24qWtcf31KHc
zfOdPnFK8wtV/TZ6zl5KBorBfOwwVpG172ZQq6mzDM0/b3ADOT/sYuHWzlJRI9/k2QU+xuCu6wB4
Wk5IVc3FupKcWe1ASgJhRs1t9E+brjlIXAL9hjeJUjtXxwae69T8I0WTmc1lfI8UJVWvtJoWpSni
al0VDjeg1Wi0ejQcRKppLsEHYJVoxhNjQJikOtqb0nGP46wrlPrwNnwcJ+J2sQTNSf69dQpn2jXk
OO03OS8LjsFnz0nlfoAZjOA41/lQo8Z6w92Z+A3JT5TJiMxTZVWsLdv8l/2X3+8+12FHbb9DUMB8
t+rLDTtDx+1a6sEcBtcmN+SJfUieAPzZobdGOqu67b/sd1EHM0Wyg7pWVO4a02zqS3QDUmVAJquz
EMIQvVdINQ34/PRerRLihd4Whb8JzrKJGFnBuwIjvaEFLCpOTNSos0emMoSc3Y0l46Bf3JYAPoqr
gorD7frlEhTEo1LSAPVhLUxug2RjWZEt7MLyl4ulS6t8rEgcQ68DchkJs2ztl9sV82is94fyUPwO
ZJp5CKFqxiurtuHQ02g1WuGSWBByt097P2BEZEQ42j1RkC5sBUflDFCOcBTiST/XU4NCBGsWzgmo
3zQQA4lDvmutEXd/jhtGqg4gc/IpG3v3IY2naeyIdrwx0hYMcOmrT8mYILwbakyFVsCsYnoqNqod
8H8enI/YLV1OfnCxRACr2MPOGranKCQ9xIUm+YyMBEF5DUnCwySvCHK/RdH4h/L26hD+2bmPPi7E
B3qAteCHPl1/tGNheJUqwFDe3wyLINv8OCPQGux73wzWLr4rI7awtVYEAqYkefmKk4CsDPd321JA
PwIx896bosWhdFEymmJ7pI4dUEngNgKcEY9Na+Hkz8HcCh9Z1+yqXImgB+jYDnpMoy2djTIyJVOR
P67HZuTGzoHaJJ4azLJZ246iUocmqw9GpbhpfOO+O2P4xsgJlv+12VjjJvgdFxwzw1xS0IRLDTWf
mzoS6+P2W/yrxzcRldFP/wtKWMj91dA3NB6jHK5mUaakn1gECDDgqbV3bBXY4RgnAd2a8Kyr+5mL
SVWUIRUQ5Bq2Nh/fXlodhJsXx6AYRZ0Gz/01Bg8FvXTVzRHogWGAhIYYSvktDt6Rd6kX/6UhLKDT
cGf8CdvBF/rRc8trhw0BozXC+X6GPkBoBN4tHRQ0VRpZFVAZuACKQQoKhQ3lTBCwttSgh+kkNi4B
d32RCJisOy1mN89UB7pmhaqP2d/jaOGfjq5XzqJjHBgbecwsk2+R5PkH7mzwrq1i2WITsMRLhng0
B9B+UlkZLaca3fITDiDBLvf4Un+GkOFt7Kl55s4kxHDLa16PUPsPmkhNcAqG9M4ogrixCs88oYgn
iC/QKdWboPSnCwNJyxylNf1yIPWplaCeFWdcXVIBGFzcF0T5ZHu4G0ofwEIaNryZYS2sZoYKoUmn
/6naV6Aag8DXtRtbmEpsoPlDEMrG3PbtmVdW5gWTRJrztOk0m11KVvRhPJiAmVACrGDCu4G0kl5Q
zVLw/pFqCIw3WHNsQ7LPlZWM9bxAAO3yjyU8cA93JgBJvlD7xaHZSmHCM8UOtgvsnx3VnMmC0Eod
8pTAOZCaGjt4e4saBfa74CXjfYKv7oxMN+w147p+nmxx8txUO37kPAiffKXyNNFEiaxyujp5VnYB
JD6wywOEx4kOZSSSKBCaWWNM0g9APbrAxMjIdwf+XVnZP4ZNVr/VO7FEgekXleA7dCf/ChrNIoud
K5SrLwmABS4lHq+eyxHrjyrLe693kEBd/QChtZvtMQ4SnBBH+wawplG6NY8Re0unNP4EOj1RLTN0
rvk9l6X5OaB4kri1/Fe6Y9xpotdIyLLoF4uSEZMcy2HjeUdZDbvYCnJG7KIOeIh/ZmPaj6z7VFLi
Z1rGXxIKJlICy1e3ct+oDu49AwWoW2XwLCP1n1Ch4HxfvKXx6V6kF8B2y+6QCDv2EscLRlK1Z+tt
twMdYWReLdKm+XdrSvSGCl7V1ZKQEuIhY+mwEZ/9aLHa4sNHCTEk0CCzl5sfeuLsGInRd8PXb2Bx
ZR3DyGiC9GpRTM5zItgfHa8TMIwaC9lHNrDlPU2y/n4ZvujSdHO+E1YzFfVLsVq/8XQMu4fr5NEL
MKWdf6CtFTuetLGc6sHdER8RO/OuCSolqmJXSYNRAdNdqY+gIZlRk7oNHZ28m33KqPQRJXc9C4Bf
3OMS8J7qHHrloBOmT6YT7XTxz499Tfmn+ZZbOB+1CTD90CU07YNohP8DUshPb4AVGf4x+iUg/eFa
W0o35UetHDMI+QdlhkirgH9U7YSPstiy9BjbKXTAOVeHMjjifeCgrzlu/HzsCba5Qwc+rEWiFou+
mtycgakl8zMHpzp0xI14W0s0WFE+FdA+NyKHRrhRo5eUcDoRbuQ+jDBATShbBkz8Paf8dhhRAuDu
OZ47alrCcURGUBtlB5g0m+bPsVSkbxQfqHTEfxEN6b41ydkQkhEC96TlJUH/S0YqnK7QC7ALXMe5
NnHUY8DyAcRPc6MQzDfGCuBOZdTDoXOEcDv8VJpdr8kC8U1zekg+92YdPOYRucmZSog7TK3B4k7D
ey4XQnsKWAFUAUK0DUXHDdotE7lyhCnsLskkViMKdeCG6Alc46lQXd+hK7M70I9LhNLiLZhyzoLx
dIyskIggPDJE8yIKjdovMF9M9yOEwqA3orQ9OiIbwr2YQeDs+99Jgmx/sPd9J4yLIVo/lGVKrRjh
TTl15RCifMFHgBcJWYXaogJVPhmAsrCqD4907j9mvgKoBiR6/hPz8XwG1YBVAKsQHXBFz1zEQXmp
UzgPq/WyvH+wvTifc3ET355I3cCMiZbaYIszbediMz7ixq9uo1ru8067pPk9oAeDHZyyqE+zgLtj
mR/7sEyetYs3j4+WgvxqEFnx0G6COGgZYzIVPU6+0xiR06SzhYcRDBKXzJCVupvRADa2LGV8VCKd
9wHh9tsfihbN9+ILJeZh3XpF3lRz3RSHyF5ymNbRKQtBBhHNYi0ruOzf/amr6khhYaVseJhVDxop
lYdmULMyEOyGXP5LcaOUig2jAK7lo63qcqAjAUZog0e83LRveyg7dSIVxhbYyORmpHVBkW4zTCL+
57a/Ow4qZ8UXa1m7pz6dB6rigy9rcrEiyKpW6Xqong+Gl2Z4KMx8VgsHV8rw1hQJY+9SNTi5hxrD
BYFrnBAQUx+/B9/T0DgtrDp/1a/81pTDBeSTVPQe/H2x/ubdvt6NEOhebhx/cmK72/69ofttNoHN
piS3i+fYGiFZXsMKf7rvmLFq18ABh1KYMdu04VyuugktfbLASUzSP3gTPu7CNuH9Be8U0hsQsmD6
FRndMokYfHvivY5+jdk+uSxwBCGsfJlRfYKONVhv0bnGXgZCVioTD1bqZNBxA8ipLyJU2NfI6zCz
irG5CKVbiMibqXRXjH/c5CkCbpD21xfhsi8+CBxm1yzphE7J/2Py4YG7jJZl9uo1xYDK3DA3x1P9
cJzcBopoyBvs2gXcH7MZTREt2xWUVzPZp7H7+mQDPOIYcpagePVFi22PTKadAAmZ0k0bwNwV4t3i
I4kRNgrPf+iFP/GhMeuKEIGI/wTqJbQdBNT/+tddvO6rne6f4G0yb1FXqsjDfrzGkHNdrWuI7PJE
yR4srH67OjqEYn4AfwrX6yqE/BVA4HkARBlxzVfj7OZThAttNlPbcBcJ134hOVmCrlZf4U98HT1w
HlQTGoBSf/8EtKN4cQZD4JsVbr3G1//95M9xhlfNjJuLE+pOvTK8bOh4feqqclHJVXPTHmDOIOJ7
A/nvb9w19FYptqY6h0ulgbOUS97CMdFvtObRpkfFVfhnb6VjWm31IDDj517EMObzlDGPI8gVFKD1
dR6U3JrLbneDM0yHhHsK3QqH0F7hYBLJz7D8YqWbkPKxsG7L6a3o3OC/AMycml2lR6elCchS/8I+
GWqdE/bqp06SZkkMjdOS+gSUgu9K1Vyf3SzR8xmaL2Hj/7fEBSBksMhw5rTQ0MNAxAVYczvjaIcA
XZN7V+AvAH/w1ZX/5yg2YW35VNrBuHwMSDV0b9c9CYomMyUANoDStL8JSYg4YwDUejX4IrhKh91J
Yl/zuNEEqEAR6yXIaiJNb5okD2odgQgiZPHwGCRLbgDvLOlBE9rtn3SsXHz4mp5p8bi/rjgG7QKi
17SWFmqrV+grQkJfH37qZe0qZefQ5pERhTdpBAz/lJr7+WYg7pCaHj5/YZR0br/D9n7I2vTHPdHL
NKShNOJ17a7nMsmAkFX2DR1CFVjvEZHB678EW09DP4r4mA3yxPTc6PIAkB1vB6zStjxQFxrRNGI+
A/a4Dlqu87kAgEolQMIxfOTggl4qGwCSYRjltM+p/ITBT8XD06P9OH7B5LoaHy/2RgBpfSufV19/
0ULC7AzHAWd+qFPsaRbQ4ebZTP8oySc4uVP7gZ34nn8DLnZs7OEIjRSZi8aw8+ui+7j8D6KnupRQ
fWtGs+gDweCzU7PxquXz4QS0+VROSimFrw/c8oJpK21uAfDK4RBkdFu9WnactuOhR6KK4EMm3hlE
Xp9i/mIykflYEbHiC402IC+DhAihlcx19UhRuXzr//5t3ISQ9BCRN+7B+DgE87LzpUDi8Fd3iAwl
PVN0vcuQTwoL9FeIKnAxna7OxxJ0fhnJjgnOf1MkkYVpTyhzoBcO15p97o9nx8eFaD3PLUX/7A+C
9MVsfAzmkJrQTnfh1YxWPkMqRrCT7U0lpp4BXenLV2OLmeo1FwE3PqNMg5ao+NYD4qpuJ1eZOqRa
fOIrP+J7z4OqiSsifWILiVj9KqSuHprXbAWybF6evnUng83dDWplQ2s1kw7AQfLcUT/myB03ZD6Q
4yNQphrpaEvKDb4w70xqdS1iaAJ8ygOLNgOmEZrNrfZR0IIRmcU8z1BzulPssqYiaoZvECQa6v37
Qiaoh3M6hXXZxAjUL005iINtC65cLjAkVDYTtdTh9udVbjh3LRcDHICHHg7vBkexP2YCkXVRY5pv
BvZURKpAXgpYJNejmWA0bx0xoiWo7KrC86vP9ca8tONfAf8fyyhKRCAJCEmPhYk5iyP9RsXcqD5p
x4C3DWkYkUVSCRA+N44Eiq/HNXO9nYKNasAWOB8Trgi0AQM6M2LQBkiLS1f6T99bArmmiWCfNABT
Onqoe/8hLMNFF3uDqut1e7nUmCjQB5+brDhy3J7rZydjoau3m64RuiBqRNFWLJAxpY6WTOE4h8hn
xPNhBeHBqID7AKj7I0rnDqWWYB0iZKPFIHxNLolOkT/beJu6nLRRlbJ3kQwUlviNehX26YVgDOEm
skuzpcQHInDjTlAzrbF1DF52udhjKo0F3atZACiPS8y30OAXlLW+wltRfuVt5y3+UHUAhkQNAiTn
lbWkugj0H54uxK1XcmkZsgzMDc/fY+XOhpxGEqm9jGFiBlHWyrpBjdlMpl0FfEWNpQ67Eg3vVl6e
3q3yc9pZaABj3WkrjI+bZPvrsXN3mGhEfw9STMPrRKsmDLTc9DNjzQl+Mn4YRH/3+0WOUiUZ50uo
x86wEwD0N7FBpydivbC/R9RPn4Tq2rI6zHcd6r8K7Vrm0VrM9HjpbIHDW2+QI4lf/xW9W2WUuou/
gFy39SHm2/yDCoZxtxSk1avOeQ+M3Mvu5qdJd1xx7Xcnrac8kDFbLDMESfcDgYCtPn3Gvdmmx9NG
xLk/nFFugPjbKuka8rLeIB9O1x8QCDLV7yQk20S65WRQfCdY/dhsm3ZiLoFRAHqVG/ldjKJqCglZ
7t68TPS+LCbQmJD5uQ9rmEyqjc6Ud4kpmrz51j4E5vaAPs9ETDOz9VHdJG8Z6nmn0xB6jczVTY1k
pAhPTb4NmmFvcKgqARjxTWEni8Oi1Iqs99pQwrRiacndX2ZfgWJzHq/AVUYR9ts1ouX5LvI4qTWw
2OyqLxhg/GPXyaIjWf6sAb/deVSc1kMW/62DtVB/a7HKGD0X2aL2lakfZOjRhS0aWLP9htQeV9t6
PSU1hR7xDBDphAhGMXwBrF6V4TDyDvCrCV2Hcqs/t2arzrYdHOSZYWF8Vd3K+2s9ZyakI1L34YXT
Zg7z641DjJrHgPc4aOOUwSnuBKRI9ytdCuD/pELxA7kFIe18uqSPBXptDj3O1kxd5tWe5Urc9FEu
c6yOYcMzt44A2mu1t7lf9809Kj9R/onoDKt/WxWmYtU5TamUZN07LSbU/WsHQxby6IUPhRzdg4JI
ORv5lqSqW/WsO5e3d6hXUWi5DRXzFLAVLO8F9fmAvA+UbgtFzPZPZwV6dBb/goPaTKlKoSknS+1O
FzD2QT3j2tWdrvMcPSIeI9R/AHwL/ZwWHEBwIpjOTu8zKvqYBzX8dP/XXrE0fssLJP46VtZe0znr
V2x0WUi8hwFLMyng7GX3eIelz0/e0fpecnyoqgIDo8E4c0Lphrx+DAPliF38Ufc8BLVkHXcuqfky
JcZjo8QG+ytdR4E9BYmcWUicTFrTli3enTsti5GMCxcMplHhWjWumQvs4oLtCrouBzMcCgagtRIe
gA7axqI3pXHYYMPIQRVPL8Vg5ALM42i3a+2K1kC0YYOQ5pQb9IdOxxhhvNPjEQhiWaaCn4ccFO/Y
4DnjlNTXzptkszulCFLWgaW09+N0St8fQvHiOxY6jvRLGzYlHo5XwXwHwP9pT7gELT/IQoV4fsY4
mMwKVIGWRcMglixsfVq0Ii3to5uZs2FkUoA7v5S11VctCh5nFWBgnlUK804DR30Sy0v+e/nLDy5i
/5Ua2IyRbZmQA6s+RGqm/4r5541ZawfXYafHx5k9X3X0gxJPNlBHMwVgQ1jLgbbuG77SsSWH2Mgp
QaIRvg3hyRTMaCgDTpPXEJt7AUIy3AOveUtkUwtHBlR7VHRafr53DaPDNDKznIYXfWyQ4Coy6ahC
e18Udxm1DBijUlOTgxFfWhOfoMssoDr+AzYzETyx/Iu5etVRpGSuILJqRR1loj/i4IH9DvSVqGlQ
fbpka3F9kBA5EvSBj12FL3Cw31M1DgOds6dc/+iMStmUjLVzyc7yyGVqBrhVsvrbe/T8wRDqs25Y
LfEZpm5SvV9EIocbJYxPPe8kP26uIMSTD6GdnNwBLAzqteLa4bCnCAWF1y3Rism6M7pAt2ECFKUr
mUrGxKkCMxw76nepF7paOtoiunutK4/lrnvUKtUclAWNKjdSk6IMurjIW9YQjVU2qN2cDX8Vqc+X
Rbcktgv30fsbJ8Quv50xexJZeXIDgL9kKYZyOlWs9zl/7WoOqb4RoTh87JoPYWGv7BUgKMjBK9jr
hS2IXgTZ4YwIaFKibk2387b1Ij7td3W9ciNurSkA++PVVi8tKPPTNR4WZp8SnUFEv2Ok2CNMfMG4
afXTPsMQRY5Q+FWT84xbsX3Sm80WGdlTSAR9PuE6unpSzTepPCv7ZFsW1vB3l9uYvbkGOwc0z9NQ
EuEKTR91lfHvu2samPUOzbqm3irw8SjHEKU+eY1tpiGtrPo94ypcnlrbY/wiowTrATLY/xkIG+U6
YC41c2c/7CY9X6WlFdZfHAiX2FcrTr8w9PYwXdPH9eWqaQ0aje0muCOCsW4A3uOnXuts3iHQqZrc
Lmm06dHRlYg+RxfW1PJre2J+nsA0lWcwIKh0i/2XcIUU2BYj6yFeGkp7EUjyxrtmoy850qWyD8Yy
hFrkCIh2JEpuhRnotetJKcyWuh/sYtXoAWUMKXq5+9B1iAI52DIn6OTjA0Xj0jcneZ2zkU02fJC/
NkcKiM2NT/M8sfI4Iiw5jSaJOgpu8V/wQLrudTy1hdxIosiSDEcap/gHhJvnFn1B+ZOg3bHU4VIY
y0DutK2j+NI2pkNh7jmLVKWa7CeT3dy7cVWOU5Z2PabR7Hhyx9Jr6oqzwvf1HUC9H0QExUHHCYzy
7lPW2vEKoAnCTgnRfCib09TA8ZhSSgs71gXHwzxhPSIGzIYwbUDIMDQYyVtHn/L6Shewi6VIYLmJ
8tvz6MsSODYes/+iOdd92OeaEDjilsL8WV72d88+mcV8g7yuz7l5tTXBJ888UbHAy44sAc4JZIuL
+s939YnMC/8H6m1HzDNWVMpnS+HvCtTZNyH7bouJsPfseYQrAecV3CSDAyS+n1+Hkg/ITO1nNSLI
0K4voQnGHvEddZQDsZ9VLcrW/IKbxFvSBoCQR4ijH88dMu2p/sSslhl7+9az2vRrAWkCqGHjw66c
ndsSGu6beyzIlKhmk1hfTBB5VLKmDcAY704vmi1exa6vyyEjzRdXAn5Q20zAaxUHzqOesv+NhcOA
Jg98Eh1GEDqk/vfWy3IXwKblFTxkdPhcWd9Zzym9YCttTwhTGC59dfMyNqe5OPZco8HNqTJOQnni
9XXlHmI3TTfqdFNQJpVcY4jCOhR9heEy0TLJarX3Z91n4AvAz06jI5nO9HMBxvY+UZ1/8aKWhZaT
NxOTmnOWGY8aEmSbyGw/AX5FbKF6hG3/sklDBMW70ZqJJkGkewSPIguqqaR09eqkXkRPwhU/ksGJ
czXXfoih7L1gNzLhM5UbU0y70IH/keyBNe7VkLCgApk6DyT3lzpyKaQOCb5BBgQwTiAFgBAGVX9l
KFFclEL2l4f+BE/Wo2/3fdOCOJnm+t6rxQitNT2iaYd5pDWbRuv+8LL8q1Z8s7VxXdZUHV7vo+wN
dTskn1ZXUt+WveZPYwjKi6UyySI1THtcUE7g0asj0CAoB+jxE3/qVm1+GGdgX/0+jtssp2c4BAZc
KPrrY7/Ho+hAhcNHGiIIx7KAzWZS2nuCuBendvgSEdLjL1A9zPe2vttRUWv7xkWYHCDSiGhnoZqT
Jqys+r0pICWYlzEqgVRHBib0pjXBbuDM+gDkC6XUeRUEqDhS5cW04elQQ1ReqkpFYpH2t5wgGeBj
yzPx885q75SPNbJS02cEfOBGKBIAompYDQWIWx6E4ecWa040Dke7a2qfIymQV6vYfXvUlPupEuyd
H1+FGqZi/4gvX0v67+p5iuJyvj5dcNsDueAl3zmCpnMjE4+Sas5OvKQHlORePHIX0p1o+ANYATRV
IyrA0cqtUkbvaJW9w+S8uHLLD+GgjJ4S4mq7y0GaZoV8czhr0l5AL7TAaLzqRuEO4rY6KJc3LI3l
QO86JaUMuNvaj/r5k9D7yEqe1nxJzzoeVxvPhKP4WUBDgNtkOUIxebeoCHi6LQlzNg+YfaUBWipM
MZgdYChdQ9UvE4mYpAGVY8DNy04hXRwpM+oBuv6Wx125t4vBYHBCc679laAk30GgCx25WmwZxGnZ
DwPWsznmFyrz141yN0CvINPZBOjBqmcFBKfxn2gKi/UsQ1j0pSFN2ARyOdjLd/QRxHUWl8k+H2U0
04eZWzdWLwHVHLR3WUMEfBD3a8LEDiBsbiFcg6MQYl+1KOP+GgxjxHSfrwSLtXL2uhU2xF7Jbjwr
td1pmGEp58XsTFkbtv/TOWhV3R0cXgNLeCGXkSE1wZxvW2nTpygV2iZSw6jxzsabwH2UOGTqNUUT
hXuRASgLIcLl/eN4/MQMwLOaU6FzKSkKCllX3gTyw8CzahkeRq+V1U7IIh2MgoPH1VIoauvqg9p3
7AGFEwmSbJFPBNTb7sUk/Ob9oEqWRvg/uO702HpbK3gY2lwWAiik7VzNrgu1/rQ/1F4y/5uzLTbU
LdfG5dqMSa8aDfFDkI5royv+dfNkX2gi0s4Kprf1N2NUiMbkhe+XSk73FmhY3S/wQ8LlhsPFhtUh
mNni346cIGgUoSwhZ6Bq67m8Zwqz5bZcCWdodjbNWScCdq4XDmqP+VtLmImPKXwzTN+DYC9HqP8x
tR/yq9asLqXMlOWIwzF9J5VLnIvq8y1OHSlEdqSygT3VU0sGriVPT3cdhXh8w2mej42b4kzL6Xrm
22QuK4+6/9+ZF7TpyoUyLKfmazwQhceJ76nbwcPaSSWutdHnDCkpYZcEHbf4NFAUjmFbfo1FbAkq
RWLtLqFctAG7nGIrFLW2sCopWqenZIDM3xOsI3IdgVOiAl2O2edpn9WF6jKRsmSihrSOAm2MOlnk
LYP83NRYcpIAUiGdF15bATXiZkjWZgHQcYSFYZsh5EtA0gYbr3lp1iHsoosq+pw9Oaxic58K66ex
8vVLYfAfGKE28s6h2fO0HHGHCRXR2ZnHK7s0VD321VLgP94YdKgYqhQuQ52OGy/qQzr/YnMmfdcl
OcDZNw0/xltKxJrWmAjcbb0XWk/xpvinKMDrdQDzHcxBTsHUkbiriBH9y7dojrlrf9xZZ3JVptW0
N/zreRydi+CyuvbDuU6AxjIMtlxDYW8owBd4COvhkVmoDvsCYEuAMEx+bsRUz/dW0sy53ey5igaf
n+BDW18tmNnvqF/uEU+wFPOA7Cx3kMXwf2K7NEjs2pM/ALk+XvFi6PDuyKGJ0y70Ap54U1EW72VN
mPQ7ejKIW4tpXvSG7kjY2b07+D7I5cmVek3YRjjYrGR9m2WXIAg3GXsx+yHmL84eYitKhp3XDVKL
PQPXs1TtSph0dSB+DHfjxfefNFeKrCg0ij46ROiTC3xWGZCpt0saqqq5ACF3JpaMqYV5kQVihzPN
O2/0lKjkE9CbHzRu7i9nxSS0vTJsIAEMpCNnfukZ58VXhUepvuH8sjuzVtUfGaCKnDZsNlvtGHH/
bdTkblnbOKV87V0hQk37oWjvygyJvyQyugwiKEytGFtn0nJWvHFuDUr6Xkfm2w8jI44QV25eiZSN
h8zwStlz+ZOczhSxraurewEjYFCilRyIG+fWR9WkFMh9Q2MiEAlsFFe9peN6ZknGeGgLfLZn0wBk
hqpDmB9z0FX7GeUJ27KN5A6ujcLcj8dvWvIaGPSRQ8+RsLSODUIlpc/Tzfq33CrNZgfxnIwCPchv
2ogQevZF5ccongFoPFl9f1im0dSmemKOtt1wfDsvP2v8JAa2P543k+e7sc3RjqRteiwGvXQyyIwP
qg2j1s3ILfBAz2n55LioMMF8xbEnQYOnaZeBUkKGT8uOaJagINSsud3Dy4YiWMRQGadE9Bgi3bMh
AV+eZc29GWvocuyXMU8L5z53NqsUZ/lGxHLEs9Iy3VGyVXdRcxa6Px6cSFuR0CcY+RtZiHeFdi10
+K5kAZ5FSnUEwuuPt+rFtDZgbdLiWa/mTaXSj+PM3aBLPxSs0Voq+iQdzlLuB4AQUjl0Bx7LErIW
m5CtT0qUP7thc0dbRhI808I+0e7x7r9ll9Xvk+M8BgodyqGyymnpVMejaLhgBAA2WrF+SWXM8/41
Chq95cuoBU1Ucm2IkdS0FOAxvKEd6e+bxhe1XcqJCLdbcs/PrUdOD02OAlzIF334QjzUVwInXPB7
XhbGbZNCJX8JMg6ov4g0Z8dJujUnezkpx3qc71PcArULK6WyhE4QZvLGhaM0KrZP6gjC+vP3m9+r
z91PIvqx2altt02OOq4lwzvokKzZN+5guemJkFJHssYwdXpkJMg9trxnZzWqEKxg68gMNqcLWEtL
KIgsAUzU1SiF0S9UTnzbBLLcT/X3wvaFS9tCLDTWUm6pqphg7qFZY21nto0ZMHIXPTQDRtnaWUr6
zEQvViViC7K12+KnfmaesqzJRAbQ3pjlZINJAw16uvlaXCbMFzUW0Hac9wApxDmMXgEihsVRmSGl
7xxFbjJYQ5JP3cN24+A2PQIDQH7k5JVLfyrdvEVkL4G7GhP+mG+wVRsI4wtT3F6YSBq/BrvvZ0HB
DloseOEA9BfjYNFYzgR+q6hySuyaZlsqdrwPAql9f87KG+voW/CkolUO5K3g6Y2hvdb6vY9pFfZg
2AticEVmu48p4PYX6lnfxe6CSZMAimmqi+32t6iDxuV8RPM2l1zR/UibnCPUrlA1KxujC83bh/6W
vVZSh2iLzklO3Rl9DByP0c7GqRb2jrQXl0frXW1eG/WN5nSPNYDrPqTvZN+PkbbnmlPKGKVOA2HK
oJduQD5gRTuMA0/QrE0SP6EM4aznHRL/dV8PSPGg8A6gd99xxNak4q9zfbGpKzwaGuIHVCmp0sMG
DAcIHbAhAziGzgKMpv8veoqjW/XsraeW8omqDF3QwjqAJ+eV5sc3sJgZXLxXALOEU/g6aKfpRlBN
GnjwjhI9eOsU52i6okjG2cOTMVwxca3xxeJvQy33JoqRcWdUJSjW8+XBEuko5G0XFypnouVUVZfp
TTEMFP0ytK1m8RXuXZ3XcfsU16eknfr4z0Jj7SMNmQ+K4NBfOTx2t18xAHETPI3jHLZkwparep/0
p9M2Y2SO+CnUgEF2UIxpYsG4C0mHZHkidWA0qpKC6YG24Cb45F0XDRRSklbwhjYn7aKzYV9DyS5S
6aFF1N+LqJ9TthvPNmbN8JY3pEZlyv7kc5FMESUy5cYbdwBn55Qy20Y4cf48BaVMnaF7Nszm/L93
XtnTQyDtamp2IOhJdME9Pm9Zuo8zIOlWwqMwMXaTm9tk+P7NcHtK5XD/GXJeydWdYd6MfnGTbAds
PqvYwC0G5Qtb5BizIHoo+G8tbZa0UoStUgeS2fSnb7XqzQrjgRqSj2U9V9kCkIh6oqRHczHHT+b7
ueMPv7pP959rANEunvHUDpDjc7XuaMDUnqsSztPmPFbK5maAM9SxYhLdBrG3TFWKq5UvyUXeYGvA
5qGujP15sEi9+why3dV6Gh+AiGCQVUDKCu8J7wsRH0yB29rO8t4v2QsaLwT6/Mz9m0ycXj+QGvBx
hw/GBgivAz2ngLNNwQlRQXoogUyTQw5vP49hve0kVAw5AThbzQqu+PvGV49n7/22EQNjbYlXtmQv
WuPkzoWrt3DL5KyEjNYDHeFJfsB8SwnfmGlr8A2PHW2+nFygmJT9c4vGKSYdK91idZ3H0+9+vj0v
pmWBJcRTX7HuYpe2doEgzdrEmSKogIuvG4ce/YA14hWomr+OylvVDvX2cHDc/DZC6Ib01QJqcOuw
vAnIgZ1t50+IaTwkp5IbkZXlEvC5jXp3yXCS0cefOjI3ACKJeLrGzwS4HYEPTPWM2Ta7JOP6Ow46
hbjckXY6S//M9c3bUcALCMLGt9pDHcGdC5ffy0ea3H/SOAkyXNozeojQ1cz9oka8H+vOeYQsz311
X38E+JDxLA3+f/gzUQDe4AE/jCsCRci+/r/vsHmQv0h7qmBdp62MZcOuZowmkMDuP1f3ZiE2wizi
vuCFo+9FV3xxh0oR60nm7No2iKRqcm74FzMNpzCfw7eZ58abumc5SPoJj9OD1jbX0neKBoRRJ1lv
trk3K0b5QCaiPgz83omsm+6Y+qT/cSkwn2dOCKTFp4RRPwSgdEd5HzMZRrPT1qXiBGdhqbRBGU1W
1tW8Xq0G6e0nLwLMyWJu7/kFJI6J6PJ1/xneVBtF0JklpXIm62ubOnNdvtLoMKxpT8/CjGYzV4wG
kNAlFOgHx25fpCj29dIvuGWVe5NE5jdjPmqjeL2u2wHhOdNabYKHwjl4txhd8/AKbO5DhPWYbv1y
MM35Y+Jmr5jELTP7wC5hEtPqfJq5CFXnX2UJKjgcQ1XZzhtoJKY4CRdezowR8Vdd+7Ftq5v/MDFr
2Gvl1KqBpttOPScYC61e7Tbw3ZWA4pyl1ejezct0qL1fBGwGouEXZs7HYuslrHTpR9Wvdt5ygRit
CnKMbL/BNLopZIO6Eh1nboF3UPYMPZKLg726aNmgn8scgR+lCMLepdnXZT8oMRiyjQsu+5eRkUto
ZszAEydDS1LQZmsVWigPlVOyDK1qcAKCP1xYCFsGwrtK5yo9BvsDWj7NWSr6YLSn2CQMcUhmoA46
hCTEJAqlacmR6Kg3UXr3t3x9+Ag9DGn0iD1DYGKp/aN/LcdS18hABroka6h1DdCpICTRWFRUNMAH
N1uFxlxAUG25p7q+GV/deae898Wnpb7PYxUwcO5nda/v/U/jcf0gmNB6lsNWWNtkFI4gctNOXxnp
HdwzAKhNSqGbcDwEuaPrRUNfCAs8FCQ1OwzNg7rv3EUKAckWPycjl53pZXVwApgRoFPJSR04byOB
aIhu7/XE2KmR6Do3QjVO4uxFqRtymjZRDuHLtJ75CmcchgXagDI1KnS296YGr/64sPsszuENLQ8G
dkqupCh4si5NvzxGg9OWoFGMm3zwc+LZDeCJ+wJD2/WEAr7qqbcKy1nNXaUnzvIfEqW8VNBQOar4
yMzrnk0GA3AYTo5IxQSNZkRaIg2E9zLwkp/mS3tC+bEHcuOcam1+7vNSvv9OEl/b1eMyNnYj8Asj
V7xiMVmJ+UhsVFuW3stn+Tl+iFD8gfME8LmE/gvhhD8UX1Q8LOyIAr4PfDoDV033rhu9S421B1Tw
0fRckS+ZUWL1vVEqKjz1hLWTk0OnOmOvDXQ4nmWPp8O0BjdfHt8tBgMt24TocqeWOlSPepR+eSW1
AXJ8IC+OnJ0LIGGTI1yIIQU8bA2YO8OTkO5QKCT+pcJT5CTiJFIfTA5KSmZJyNBM5OZxYafeoyW7
TYI4oPGSaucIgVAQbY0HL4GPm5RSjrFd9/b5Iii49pFngkkSvhE1nFnk7E/NmQHlHv63Q1Qa4wNs
S1HIPUoa7Gwbx8Hk9eHhfZQ1nbALN9iXTsYZVuMWNhTp+xk1BfIB3q0xGqUeZ528Xpej+NLJzSmN
BlghwApKBAnMqVdQPn4JuYrIDGhPpVTpbNWZzo6eIHxbJ+6bLv2X8k2HFD9imOs/NPs4Q+DMFEgO
/rOoxK59HIX+PHdUETVtWIGPXuu2t6F8DCrfZtr8KPY8HWVBN4g9QEC4nWnOVHLmwBWwaubCFhmy
LKhBJsHUDPFv8FeM3vQ9r+6qH48XNrnimQMG9lWKNg4SR4UQSBgg6Ucgu64CWu9G4GPCfHHhBoEx
+YqZmy9A85a4yolbZLQdwS6yCUotDeVewFcJRbFG9+VwaPNwY2yQe4ObgCH/JqWiMWWKCWLY7QH4
zolmBAqOXYmA0nab/C0y3u8sv4RRBYN2JMVyE/drGThzZaaKcIKyjLquAXNvrkygvaW9qB7NhZLg
rwB1mkiRs3iXNwHUibp32KQeTxkcpqGijT6Kh1nQPQPB5amoDjlau5OdZb8WleyDp1vlTSCy/5a4
ZcnwLeEq9AoDVc5K1cbAOCDIrcor+MPUAtyVXBEwZZIuWxyZ1/vqehjbiUBGW0OCfySZ2F7tOlhn
41UAK8ou22cO5FXQiwld4j/Le5hpSO9OU0C8YEHwZRrUXTfTEmxEsqu9h7764qLIyALLltCKhYbW
pUhYMPDOoXwyhOhfbFrJnzavnP+6PH3qNPyPJf6YBO6tE+5VQWZGWdXS4GD98muBJ75yzieP9ZPm
8N8J8JW8eb0upiSv/glYNIfzZYrARWjElMlnIJHfHhGDEYbdR9HQSw03WwCXgvjyGv9+lB4llQmU
JVJUQdMqOeroM65/RH4flF3IbThXbAb9S5gO9XXvMTFS4i+AxuVUf5bEXIt8dHCmMN/uxuhPVNPH
R89bumDilfy3ZL63PsfTo7SHXRhlK+SmjnxG3cb8s1A43MeybqUmqa1s6lUnWxAhCzhjnn7sHcNG
/DJardClghI7fwlhFiAUSQOqZkgxMy1dN+LG5DDXXVxrG4rOg6Yr/BMcj3bXK+DhI5TeBkqjrEwA
Iq4Qj0iV1TYznbz9XWVF3TCCjjS8wH8qJwhZ9vGPPHItd3EMzhZ3d5KFfrFMHD5xKxuCvP9WBi3+
ezSivPxqYBPMLBn8wZdaiqgrj9Re3GNO41cwUQQa0ZLHS3cR/x71x/g6v2wgghlqgVRvspsomjtI
jbBpYbrpgZ5Poh+TegXU9gkNBhXfZOuhqAOcEf19lyht1+0lpfmXDwU8lEsQBKRTpiECu2zPD3mS
dQZ0ZMSCzXqvXUuqhrSfeCKS4wwKa8Vrc6WjLD1l/Hxwu4CmkgbBBOuESi8NlNTy925465m7tTC3
ExgZsmh5zxBPLOcpPWUpKUa4UiOo4pONlrWrllp6Z2hIYly0j7oIkRYq82panFYnPlQlE4CSvmrx
lJWbgAQOWmjDuL5QX/9x550rgma5VSnRcLRCzevJZ5laESiHyiCOW+U6tAdMhQy+5cRzV8uhNeTc
fjtBMBIx8hnbqQYnotlKoBDx+xxDp2aosE8uwNvuid4cOBYeGH9ZUeNV01uG6osWICJBCdgDBSzD
HHKXwwQElm7LwzoAeRCXtF9fFTkiyUW7BHC71mp7S+nGsT/VY8LzCSSkRpOAo/tAvCywsBH9sYj1
LqWI/A9vmuJ2+tFsxQ4XRt+MYjRgZ1Ig5Hm+V4DuP6xWpa0I4YVelHtyuSasdz6UdjzFyXVtc8we
iKofJPN+/tU4ThBcmLi8EQ4IGrIMspUDbBxAglR/lZ/VE4JHAM/dEwkVj8Z7QV5FErViYk17eGE8
RL1FEBpBfVbZvrrKoUjTQ+4qMD7PToVfmXRndHrKIOriNt8pFp9PFF+t+qTN1RxZ+xFrMkMF5Ph8
XeixV5jMtkGpac/yHWvlRF53QrFaC9D03xePSgiBGibRAxcAHJxEf4Zpe8qUUwJZwR732FkJFozp
qx2BfL1/gTavc1R4QN+vLZMckqSjAushMNCVtdNDXMbVg4iFv2kgvQURAL156bu3KGyYZ/XDV3I/
FEwaf2wReOJ6u4DOFU0By7WD13dJnf3CoEs6uNV2evKVfKWemLTJq7eS23Kh30Hb8z172ltErgRB
p/pe8eujsDwJDIcXxmriuN7RUNNiBN4w3rHJXoA2Fr+sEkyVqlCIt8CzLmQEmFRbR88S+GmTx6NN
TdTxHPVTwZjAfPQ8Ohz0v3AqZ1wbKU+XdHZW6KvcI1vo1N7gCLvRhO7bquyTpCwgIbv1Xq8nfJ0r
4l+iMr8tCNcD5SP7XeELI9qxxhKNXMqaqWq+Hxp3s0ohLpaKUhZGRk46EnAojqMv5cdjM1WkzRZt
A0pc4v8+Ax9e5g9P4AxZtFvlzkA9XwWQpmhQo0Dh/8n89W+xb+VkxHjHy9gzouXeUluuLTgL2hAc
sNx7/99o6eE1iqOCnFB5wLK6JQNFqEJdUI5Shg447RKQ5cS7CG7SO69OWDfX6r4Z101za4A/lBIF
6er2SFAM7PyXDEF8nZ2wzrxbHh6o4mw8nKmm4oFtNdeOOFxdeMBMou6nBvNq2QGjsZHLHUCKui9d
ZfhbTpZGTS95q8s8ikVM/ikxfVUyPpeozgQpjdB16sl9Fcf16AAyHlZx4PMy86ML9gthYgPJv7Kg
ubQKfauxwPfd3hdFaXeqsGwt04huTVb6TXsc9v6tbdExAxmWtlWyUSKu4z8e7okqmaB3iZCNwR76
OWrwIWdTagWATo5bQTFJwFWHsc2z3fce5LQ+yH6V5t+TXpS1b7FQlOV/p732i0fUa5vAA3+qfKWc
csPKQyo8m5crYKxQvgDdnxgE039H3S6sbfrkeFN2cnyP78kQANj8LZ7Gwf5IE/iiTRquwjEbidj8
5dOaRXyjAgBK3PkB+pBUj4azVLXDvF491kcg9gmoS1XaOhBvHwdXYsrYtr8dpu+TfdVCKq0HmbaW
qNQyikv8arPNK9ivBp+4+3/z6UKD3sFLojoPQLafXXBrNxSZjtDDsKEfatOsmZevEgB/iN7yLLME
3eP96Ao2W55UKYQDiGX+I3W0T4qS/TS/9sFZy+jGK7W3gpIOqzWGVaVACKqMOzBYOL9Dw3w4h9We
9KGvuuZSIi6pxo1OFI9xq+V675UKVXuU+XCuqv7CAcGj9i71SDpoVz9zH4a42YcblX7UZJPxwvs7
C4/bSD+CTm0CTnwZIBw4YLMtfQuBKOFRIXBD5h0uK0GsG+BH4DiDv9YQwqH9sidB1+K5LnOSfjl/
xyghVWGvylQfpfPSjTmDDCXegyJUuMTNcqmPOlH1V+n7AH81FjiNfS8LwCfDd8tFw461YIyqmac0
PT/PcHYtauLzzkNrHsDtH8F20ZOxPDkk111Oqy8qGkyrmUNOrTTUo/5ufNROdxWlO2i1LW+ovsDx
KlkfrT3eNi66H5loTJqVt/fszZjbemBxJ6yQWqqZFDbNsLVewU+AWqladCaJVf0ZwZ9adHUTnu7N
jrnPXj2po3+U1nZElqq2flH4tUZU9vY0gbvyhsKDVRFRAcaho76wdUcVpS6BTyS2c9sEzpIZpXt8
j2+STwJhySvHOqufEztw9p6aTqkDI/g6gjPXmiU/67+FClXrjEOe+yvz1w7D+KJRXxPayISdw7zU
NqQTrJqFZi5bf2Nimu2xfGiaSsEoG05uE11JlUOPR5mQ825Ko1p9e0oUQRyPSn7VhyBkduUBuS22
8mC5bNY9Hwk4uJWpGZgusp/DUXmMAec3CElm3iFCtJqlPUl5r7f4aveevwNS4a2XkKEXcZXJZi3l
ktvlXLnSVl3uLHuvpeZNHI1Z7DhZL7WivmnrjW3LmyWiK6KioOwjrbExFY/nVCCTJ+oL3Mzkr4ji
2UT/50rPvcS0cjancgUHr8A5LOKXCt3Vmzi0d5qCID9MCGlMgzVCEzcbrPJFVi84d7nHH8tF8tiy
Ujna3TTfwEQp6dbAUBMPMEnAE4DS9ADJGP65FDOxhydHD0dkBFNjw8+2tVsNoDK6fEPuSn3L8I/w
sFa13S5M/tYwWSxeAQMn2XrNrEwqWGbHFRfF0UWX5k0YHYPZ3IAEK2Cilp23c43SZoi6Gttm+zxV
xoQVbL402i56905R92lS/u9tEHE/pk8vxjeeTYhKZbbUu6pYFNmNou64LF2hTvKoeN+jLHCaNt8V
TvMNjGpnypLGOjt/ZHxwrzoG3QP9U8jErIEYqy8W+8ozN7GXCBC/wooy8n4n8raHeOo+id8cr05l
hWdyPwu7lTs77GJXOjpmrS9+bHPB0abaCTuOCSy25TZ+n3WAv4WNrFewAiFx2s89RSKGX7hG9xeH
6cGoIArLz2Ee0gFV3PBZzNoAhmRQLZ5CG1BruSQ2UeTcdWEub53yzOuJK3D5q47bUHBVZOYel+KF
OrYhpRv4RNJUlMhEbZE13bkY8HYvlCxIDz6qxpg8TM2bClyTU18+2dq0OCGafP23OatCWeTlGYen
XQVfdc+5HvOWFEkYv2Rd1AtmF0cI0og3dnhzOaGT3CPR4Hyra9b7MP0FxwactIhlbxEbF1/sd8Vl
EBUCeJ/oEddVljd6/GzgddCh9zq9INc8gDD+r0T3PQiibyUHM23nrFd4biT2Cwdr54PZGHcadZgE
oUJSnUD2C+cFXvBVrORJntMoCbOCvm774zuzaz2kj8DG4lSzC75EEgZRU3X3wJXCKupnjVr2y7Z/
MjR77aJ5PQC2KgA7BoYWy2XcYDqrfvHRuB/+fzpZ75YlFFTgg3+uUUlJ2TwC7omtd+YPcZZR4+7a
v536QMy4qCV8vg11ch7eeEhBEdcevAhRN297aKy+atd/lPbAs9BkDO5Wx4raXB28RMDGH/i64ru5
BUsRFDxvK7dshKPyFIYuQ4GFFTAKFltQbwH/0/nu+I1wvseX1qtnyOeH8GifOqaG7ueF84lnY0LT
6/zfKETDABuvBFtjAsFB+6qMiFJ6AUXg4NNhKwwm+2xSqFCd/JzxkJ7YO9pY0C9WMKQDjWgoBePs
ceRDmTrn8Wme3EgJu021tOkiymYQWqqXKN6FN86lqsB2PF2l2AemcrphYrz9gR5hefbfNKS2O3Kq
1a7XWeXP2XFgg5ezrtBTcD6Qz9xtUc2RqSOBuOM91o2w0zvwb9EZufDcOhOorHx+v5HNPKjrlhQc
lldK5s6ZA8iB0j7qUIBi/aTc/J+kGhnPOHD3WpWk15XlWcI1B1S0Yeo2Vwu093a38eJgfSUBThaM
/n9wNhKxxjem4v3uCTDIrbV3aRaqDWk3j4vb2NwddDgwi9vT59eu58WkIWBYRhlQuyZ7WDLKEhWp
S6kZoom2+ra7Tu1xzyYl5qqvG9O3yw4Jk506SFbtED+XnBHyUqpIkRLwl/qsPS9IgRQk9sf1n2+R
lNMlNVWw+qZQhhfC7SqXp3gTK2DvL7BbvQeMDCt+qhIfwJy4mIRm/K0EEtBEMBoq66LqUFw7wDxD
D1OHoZ/3A3WJcsV4dgE3wyxeDYwCl4ZdkMzkpS51MNy1/J1UCALopOry27FIZaZsYbH4M3QuC22+
lZ23jH72HYgUdcUXkVv967HupbkeXwhe2tAHbvEoynHUvzxF5mqhV9a1BSjnqi+Ds9VQDYHjfVLi
9Il905fbXSLYO1D6/H/rD/BaL3t4HZpAjMv7lfYFZAZofoHSilwAL/E/cS7VP0Va2ZugxJDuJacY
6PFjHAecvelkr29EZHEAE+tyXvyjYeNeI4WxP4kyHEDXH0tkn8iWNG2COz2ZYyUrvXctI/dJTbyC
PU40TabpHLg2ZQz4gJhy72GzAg2T5UPFUgW0G/gx8iZVKkEdxyu83yLpL0+/YcvuMxuVaZT8tgzI
0/PteoNu1HCNWmcDEJ/KEswBguoKbANvTeZfrckh8ipmjwBHOgBVKElSesCq8DbKhFP7ycWxYUNC
DR7qa3iV/Va31ulssyllbEnNhSXBJKogUlGnwbq1YArbnc2xXlPlFruLTkXszFCdr/CTb87K6kTz
hldERRHys5wK/yah8aS5bLwnMTO74kadWMFa/YzK4I2qnlDXgU4COAidDpn4B7E5RVvPXeBbqPJj
Dko3fAi4o3QMEC9TYyJ8YcvEPA4ZRhCcCJkCQkPzdOGtquiVZpM7CUwxGbMvBpLVLZU5RQEoFbwv
rzbDzUce3EUbtCIHoLHR3/tUENZkASnCXg1WJMsS1QSsNIm4oradUIF9d1NQu25ltIygGaNxYrT5
Mvzb++4t8tk7COobh9GGqMqruC8AN8zkVzP1ckKxB8TUII2m4HZXVcTcF0FMPe5nXWnJJ9/ckFOv
QhLSvkEcwpUTpcKcGNq1gTM6ziAf8ptXVPgw8tqsE1ZjD6riacmke56vLx/ISGOKTPMv/OsKZaVJ
EfxsT16FgSFR5z3HxXD0ACVKfRuWn++EGcr7jEC3hoNQsBOlWXbo386xRfIMNw/1TowCrSW8YAD7
1N6EGwoSXbT3Sby02PIeXhxth7Jg+cefKUes1jlgLEneeWB7WuWak4LM2oWCHI+6vNeM9hmS0jC7
/q6oRM78mSpHQHcs7sMBLeeqTdLJMfjtlal7aWTSq9FyyH6Kwpl1uOjdGx6rytqLsEMtqggTELRN
/rG0oeiOatdT+6JXGwGQJgh4DRQE7ce0nEayI1ALKI8a8h68gZQ7SU417Q+g0WFTLM+cawQejyMT
Dwmb/HAr3sKDBZ9aO1szG/ocsVFGQiwG8cX1gebiQW9Ilayq9Bo+BO0svK5u1kPMjfJD1Cf8vnKJ
tvu/USfZXF83kZb8Rdl1TNi/USJDOk2zUp5WY756G8F0kqmcGS6LdUhXBhMm5n6TOMrEc5vupDOK
NVmsR0iyoWwXxjYcNoPVJvkhl2hAPsAJE/9H+3ABOqxNgnqZuKB732orBpOE62LDm+//7b/UyCWM
2gu1bIKZJHCRfGdFNehshVIVZW33SbzucSvl9fA0V3Aeo1vML5pta1vcMWdNR9SZxPswuB4KupW/
GvIaPpjAlD9clkyO993XRxZxpW9W8Yhar/x0ViVnftUNeayHrf2vmXmAWW9iXv6Jn/38DIoR5A2Y
DWEASU+spCDZUMothvuXW078WHfeSV5KRziLa9Tz77ZRIDJBbbRoJIbyKNdAAfO8+OUUlcgu+KId
x39Kxq9ddO9wU0ce8HEJb/cCYH/ldjGNxT/RWXMMS9C81r8XJqtYsOckcDc6ob4gpHVfu8WCnMuu
JKgjXVdswqByOHGedfjenwhKWk6Vb/TA9twVtvK4tNSpADbgcitnFvpSCrLN8R6qaYa3taSc248Q
VGeAk5Arhspld3qykXMaTkng1SI4sULup5V99q5ghzrgYKm6afKbBxbOhf+LI7D06uX80EO/aPOL
SMv6lUEEOiPtDOd34QOuqhOrmaYwXkIm/XMXqRWjPe+W9rOsw++iTNnH9efs1JHwW7lH791NKNR8
1Kd8tArpBOpNwimwPDXJgAz2EFXYXVsO7XRlmbCT1lKNC7r+JJQGNqIB5NGdpC5Dff8oPc6uitas
VjzOUO28jkDsEQ0ZQC7/WUGj6sTo8k4QMjhrkpULJCYtlMfapcpv0puNT9pRdv4ISItHm+SSbMeb
Idm3bmYoQ4bUQdmhRDSAAvCCcxrkSdSKnIOuYHj3hvd6z1ix2vZWfL3C/tcBkqr+NHoXEq4C5q0V
wjZWOMLSFLrbwAmRp6sYDP5uVUEEGd/9lp8nVvv7VNknTNF2AmTXJr6rzFGXRS/D9z8HqmvvqU2n
SXewSrmzNfPnGNS79ClIZm3oDal020BVNli/aPlhhzuKjNUouyAG5wEsYEX0BmwEU4vxq2utZq4R
KpgEr2vgo50dQ4irwC2qFQ0IZzibUX6AEEtfe0Ls/7ugCF/812gwStzyohjTcWM+W2d/FDQMqwx6
d0tdLjBjnTWUABFgTtBIDrsqOwl8+r8Di8TuP3Q8nduHT36xM0YE3PPhIIngkKjBM5CsMH7eedxM
72rLDYXmmU3/z2dx3UST+hD+g5HD31uW0qw89l/LCzwWYHEh7ovq5wVdj7DydDMj6OzBdTDseNIP
UoOwG8L8NpXsAdZDGv2SfGDAmTUe4ldWZO5J7KHdipSap2+4FbHl/MYKglaXbNUNVFV3HSWHr0qW
Wid91P7YwKKkamDHEerxXV4gIosJMjqiq3QgCpoKjzO8o71AitgOHJEDUTgg4VsGEU4Imq//EI0K
HRiXUkLIwpyvXUpKq5UTVjABNdecnn561HozCUlsa+qN6MMzOMgMYBaY8yGmURXzUubNZ1kA6mmt
DA85tZGGj/oaWb1ilvEzljv/27Mrbb25JP8eog2eDZyz/bTvKbVheXng7JSoi7ANI54FXd71hTBN
Vkdir7U/wG4HvSKE7QpKBS+Mjp1wLeAZ0avWPSaZELmXvMLquQW3WiQxAgW9/POPsLmf1dJR1zBH
me/FqxJTq+WkcskmtD8Cl1xMq5dwUm/FVNBO1BIX+3UYN47Q37pHl6tOGyQbKN4nz6jlHqw9lDtH
4yIkpJUk/pnTOK9D8i4TiqPeDDquQ1SoOfzA75PjaUlWRid8LlR4ALY6aJ7zXWu/ePEvgotUsYQb
kwCWzd//Hc7k99d1uCzXRpucuh9b2x7hL4HXdQVTBFnA1Su1KWIPbShUhc2NzHeDDRSWzSXYUzE3
7KJg+PkhumIgi0QkFkO+4SaKaZRUKf5DcUX3MiCdEizri/8IKZA+HUegSjRuqKgl5h1eJm0pqF2V
+AKvlZlXmTUSVgmkY4CBiK1zhOn8aPiyVNmVF0Hshu15Dzt/1lN6QyjETTdrYZSgnrTN6KDthlwq
Q3o2ltkjK0GHkT1uR4oMldjidKd/HNqcO4MFtJj5q8gUisl0gfkeshZJOVwYILJFQwm3j/ojxJmN
GNqgLKV+JpgfpAIooz6YUCY3dTwqgjmDGFejVTPhJ7vtUzWHgDGx8P7MSlCS7tmgnEE5Tt5+Lm6o
hJVZMDng87CsEKp2deEhDcDiY1SVVgZz5Vgl4Nw3IgdJaB2imdWYFwz9CG+c2SoKcuq/ZyjnETHO
YC+c/K3g2MxT2U0JKG03K8/hLZ4XtE3EokTmLqX3Jxp1eSdIFXOOEEqyKBHgmmrQ5JKrhSuThOJQ
vamdkVDlyOrXeCAo3/oziKqv96lnWlTqUHdZbEvxhsdDSB8R5NSqk2/upcJFwMd0lvbZP3CQL34W
NQRJ86DUvMnhfLIOIrzQH0MTwie3pBVY0+En1z1UaB3Ha9AGf9AZoK20b7HIiuIRtQP7+3tEOMSU
wH8lH5Ix334XncPStJeKtBjuMo4lxRXaxagY6+F8K2eqbTdSXP8X5iQZN/VFjfF+rX+vMBNV9teM
CojVwnV4aau2Qbm7X8mOFk5AEv+EwzLM6oQvrJyBsQ/7jtwxGWL9hrMjmr/CRRHwzRXpq8KFuOI6
OIl/ClQCUq4Nr3HP7dImM+M3pSz5SgJIS5mmO2mzpeAlEuB+QuRL7G+cjG/oB4OIGkut/R9j2Zhi
yMDGNBK4U7iAZUr0Okw2tsW0bSWRQ9Btb8tOplx2J4GSFRFnqcs1UubQknaxrHHnQmO+NBLUZWDO
t2JCwyl4k8aYYmp/Xr6FNOdYDoK+soWuc8Z3mjt4qKau7RTgrK1NS5bcp4xw4MKNt417NPYHMsId
to9pLwwV+hIULmmrPJdHV3fg/sq4ojXSirH35WU6Bg0iqIVpkMpRcs4sDW855tPLdJmmZepIhODn
Lo+BlsO8ZeKo5V23q78VvM26yxFxLW35DEFRM+t2CL3LFk27L27DhU0qBTBao5nm/cnYFi1MOXDu
VV0DALk6+VHxPKF0sJ08QV6/EsQHnVB3n3uLqrRvxuFaHunNaqSP5WN2fZP4QtrzGix3xSdPSxzq
+H2R9RXCB2OlT4Q1CluU5IfnqCXxIAjgwEquZL9EBnGx3MNWGh8YWJgnDyOQOc0uy6nl+OH1lXnD
SDSNKc4i28W3xW7Dl9c65+uba/MRvk3Nl9a2+CD8ZJB0+hEI6+FhUuOrzTTHfNnuTB6UJ4Rnexue
HxGWcjySXaJL7e7E0iJbbcO9ZATF4P9mfR7nngQE0JNPCaNxan7MkrbiyMOG4XaKEWfCx3GiMJRz
YHFp/t2883zXc+ccZ6C3mWRr515oNel5UdbKczxP8YzAJU7BpRtWB3Iw7pRAe/fhwxgPM71iTqQ2
IzgHYzXMRRnz1Ffjby3fNfkIn/Mvr2JQfjRvpe5C6lu4+AnNK9ss78BKDBEOwL/lowsQ3EX6URj9
Mlsl/EKAJOtEeM0q7GF5PLaUKuFBkg6hrmop17K6u0xY6CgNtw6DnIFMSwY5UYmSR97tuIQO5b10
LMu1WgL+SGUDB/Fnng42SzPQXPrdRahMiJD5lllhlsWtKSpviugNssTj/qe+wZ9yZE/9zTLsQxs3
w58InUY3E3Skek9Q9frYU/7g43ZWE5+ts5XhF+6VaiAvTOFVHp13pbQQcZRcvZhb0gUY4xMy4BIz
zS+l5mmokMaYmCCH9k5oALk0RYGUMLZTxMPSqwxAKINO5mqJMBdBWznzOiLGD/Ul/ICX8cGVOwPF
qdfoXRwkB5lLk9yw9MpP2j/zl7jK4yI/fNjcp45vhPtl3mjL8gKfwc5qqlMKPfodeSKXLovkhJKp
AJsvLJbaZdNHeW4y5ikdstfz5KRaxyXbrPGLnpSV15sp31AMDTRRrnql2ciChXd0y4ewf/XyAccj
vpCB0zJeqYSjgjzSaC3cM1q0+OotGy/y+kY/Sm1UmQzy+u2fHkllVWc1vHjiRdugD5VEtWALv/2M
F1/ySI7Xk+OpccKRKGiEk4lMfLYmRdSXIxs3roDFBsQkz6Cd2nos7KPJs9eoTURoYwNR9tn/dbeK
I3FD/KTMWO+nTzZofqRBNEfYphd5kcm6FlDsdWaaA1t8cY53BPQwgJ1i/8wuWLthbyZvA/6i1txt
rO1DRb0IWWN7RnMXDONSnOXaN2hE+WaNRijzd/gYK1itBF+dPdaTowX1/LwVEsJSEbhKlO3vjHhc
ftSLZQBOcylQSCkjxtO+RpRIRuBJ8Yofpy29hN50gKjHDxGezebnetCC/6Eo+qfF+eZnnqyMTnIS
4BXsLg9TrT2uhcwhjSF/u5EDFWFAC9Kife4QXnl+Vzn3M9TerSx9Ay1sr/ccTTrjYmPHptaKcKmM
vFHrR+G6+sX1vMQK7JWY453WzjOulACcMLV9sjL7Qq4GY0FM0IPtmYwXpmxc6V8fCbhLsfyHizsb
R9zJSudeqWEgBqJHUtISInX0M9+0A9gMwJ0mqh/uqUmJhiXtiorZuM4l1fBtDGAR2Mpo4jH93H1J
gPx0bGTYsUL/RdSOwOrcI12IUzSw+9DL1Y0mcGf3bg/pqjnUc2wgCUGjyanV8uo95yqq3Tk5gGBh
7jTVqLSj9P8enHwKGGr5g+mQAJedVC9WF8eN2eo+X3sb5NRRjNBWnw397f0M90YnP3esu7DZacQY
Ea/VXhwCcXvzc4d0zejFq0s1C6SmSCPZS/R7d3uXD1QUfSFMUHRvrjj2SVaAstJdNpihYu2iqh1e
l4fmOFtpSGEu6sADoodXj8ymgjbpFECEM9EODUB0ZB06fYaPkD2NRQ51oQ5YrWChnSX5p9kL6ym+
BrRM49KXBK+GaAlcPfPOCFTfkjG4grRFJsqxE0/hBmjBuMJySDWGsP6SvlkohwYEZtEMsRu/K4bX
jX11guCqvHweLPGGR1IJifyEoBg/ssfY4oKyR5exPzMEZS/fYvMrzWcDCfmUhhPW5ti7ABMsTSoU
MdWijFHkva3A/wPQ8CWmRQfjMh5O2kPgMG5PU/CWu74NTaIVMn6xqCvs48gjoK77qJzQUN28X7lY
+ud/iVsxshmHORNHcf+4BlqPjqAWj6aDL8Cf8Ec5yOH1xRSs9myH/wx//QBs6LZhNpceo68mUm0E
NCyfgHdfsfJz8TnWo6Eh8MJdMkM1bkNnnPEIDs0mmicLYwmaOtj24CTbOqrLU1jFAprIeIAFND0v
f1Hgaf2kyGO50cs9K94baa7ZvEbTnWWrVXGc/lGDb5uEdRaUlDdBN1EVoQx/et31SFF7QNcdEnNN
K/nv1iCYhfJy/ZK4lw9LoRAL5degpqLrFk8di4H9OeD/mCAYlK16Qk0os8rC0FWX1mPCxMElukJZ
TT63HBfvzec/r8vW0hPPDafaLZEuzHKvUJlucXiqMhwfFxUkMFiyv/gW7FuuIjDlEcBhSH9bTG3z
ezPb45WKZkco2e3T+jUxHTnuKFW94vjR3RuEQmN2aiwcpT+9SWkqdHcdZTCu6VMwzLdzuoxuzGIN
O0TI2W9ATMy3xXLo4W+pjUuFVvochTi0z3GJ1aASkoYAlCg4siPwrjT3nF46qPK0JjRWLBZiCcKd
jDeKZs94K+0zje/fEcTCaS275K61x7aXou5KefSTwOa6Dn77wsj+YgU9xn9uio+LDiIPbcNhmDSO
Kb6xooxGZL9hJsNI/8LUzoqBeh97BfT/Dtlo+8sHB+Fhp8r1QjHaHtb7uLgCV6KsZkB9eQuJ9yAL
5FkETIsUZmNbG41J0LhpxFxQ8E2aOX9xNsDJebA5P6uW2ZZaylflx+9emMh7Ja1MJE9Q99anmp8F
Et3Z85QtjfcMTqgsyKubILTfnhn0n1wX6wbJCTDCsAb4z3N6WL/ZuGRl4ZFVi4KSVgqJmS0q0elN
2pKDm8iiYZWQSsu1rd9T3YO3sjLlbelMQprVMnS9AM5sae8xJgnw159XgZezudivtwotLGqRhiYf
h5ygUuwWOotJvDJGIANntgujWF/IzJNGkRwVjOD0xfkbw2QoOg4QorR2eUJo9nPQXckjxpRUHPFL
uLNSr/FevUc5iV0kHw+H9CSrgd9VIARlm9mOonF8T/3Og05HHsQK702sDMoeGNzBZ1zd1lW3NZh8
u/CqXJ/bWP9VfWy5vFi8Vyb7aAywtRsP2kJOcNjDbMcATIVRy99M0a/uSjheazbW1xw0qc3NikbO
PX1fMNp58z8JkA01fn9SwxRdr2DSSM7LH4s2VAa+T7dXvyy11ndiaOAUmKABrmJJr87jDCtkS963
dMn+B1WavQMawMjB25Xw30I/FJiK2MZ0yGGmwDrdQkk+vwlqAeN+Ob/aPHzGnRXO0oQsuDyu4R/H
8zJrAIz2oVF3Vh613ViofZ5wSbnXS4lo6RzExbHCRCItTD+R2dYd21cUC9fBTQgBxCqHUsDcJK50
k4cV6/RNEU1p9vJOainljNRO9P1OUDPh/7b8ZSNcpNsSz7T5v0wBH7y3Xvha7tRUJ0hKqGPhI3ir
pgVofvvpuLAmUizfui5+cIECfh4xg54AF7ACCTLoK51q5EW8IynGfqNd8y2HGwLwASGqrYboTdRL
G9eojA2HaUe0TBQTKkKAg2x693LV4HK85kxy+x935v3FnIzGNhaUHLyMBli/YtYOVOLzXACYueY0
4eg+mBdEDjPadWL3jfA+s3nKNXMyVC6Bw039cSd5hXQqWrrynbimp6E4XpRE+qk+jYIvICw6ufpk
ITpsI3MvfJziE/F7ivVZ37LnSFuZn5F7gfm6zEBOVkGb1Kf5im+bxYHGoyMW7MP1VDUlvWKx4K1c
iO6KCTN0El9R+trnw7dyMlLhzqA3r9i8wzncAzoLDStRpORNknZCL46BCfDHW+pWaC4fTA3mpcCn
2HuqkjiLpoYYqyJYtEf6vzcKvt1YBgfwYKhrExzgTGlJ1Ckt79OzxCENmQFhGZM20os+89PXMQPh
sTPsz01sRbnwjyQX9LLL+/XF9IYqUbaHoXIEY8RfsYQ/9MeWXKqYWOCSaVZ7CN95ZBp+Y+mRbiRA
WvW4NNFpukRisScxWyhKdrc16KKjbMYLq9KANVGW7lH52GBr0Re+GCbC7wwL8oORoFlDUZgt/Spz
VPD2Az+2Ezmu3AiKjxnY7qSU7gB1sQ4rf2wQUJuT4iEs411/DzfAZP4mPq+S7O0OvBtU0b+YmCPL
Nr+X9MBNffCX/SzIyEhNiM1Hq2ZWnCW1je+AiBYIaBj/0vVOUaL72JCGfiBiK3w1o5TNQYk7Xjgl
cGPwFP2j4ZtzIbB7RONmaDCjPzauj1zlBbwlLcyDfEveOJ0hfcHKJJZ8VBCA99pTh1Qxtc9Z0rZn
ku82yqUygEb0liS6sqpa3NHlsQw3x8sNC56OZ5ba7Jv9PcU1jk8e3JFRb/2neMONpaWh6YJzA1pg
24MvsS2uswSMoHAClrSM0ja2NFftYgjP/eA/km1sXcZMY3t2oWun5mcDgV0zXIBRdVb4GQykJnWx
/EyF4Jv5HuX6ni1jaCaqqQtlXFLZY0cETTaLoXChkF131r16XQLmev7B9KaGbkoL8MdozMbc4xGM
4aWB/813ggGiDLuy2i754BsPMVjncv4NCEpElCCciU2sO7ypyFh5IU5osNToPjXrAdYudt88/aDD
/fzRCmrzdPwVbApAjQv0UKwPJ0SsR+xW+K823GyZoVpjrYyRFiyPYn5rzMmf7kxhdPNaJhIf+c6I
HK8ShfkpdqsXY3fhr37YGvhoTAPLZzwtwjYxxU/0A1QP9eHAskp6Boq9bMs8pQekV4J6ziK/3l9I
4JKvgXJ9tR6RbwCFM7JBXFj7ETGKZl4yzMS2i5Y6OjIx5jGpCENbptzzRFigeSEJOXMCFbfvImam
nFHySjMgNwZkAN67XL09f47uD64jpNVxtbA0zThlw0fVFoGOvHmwH4RlDXgVaOhNJuiSpb4LFGAc
yRtIHohB27kUvJF1JrHssewSvol/dwi3ifGQVG9P+riAWCG5p3XpHWIfoaq1H8Lcw6HLGF4zGbgQ
6XCMoz6e25rfZgRZNY8Fl+QlOJ5vi6XQKXMXghfMv9CrcTcJLj8vQhdaY3nwJ2MgQZgwRBE0eZvB
vwCsdvA2vSBnGw+kmVphcpZ8qEToT+VsEsFNzYeGZWQU1imXpdhvENpGtbrqD05cwFDxI21v8e2N
WThNhM7BKr8L50tIBuUsSGTvFm4C1tx7dNBF9qJtTWf0XmaHW0AtCQjVZtoo5nL0mu1WwWMgV+ev
xm6GLbeXDV3fU84j0aU4ln+zvIHmp3u/CJZ5R1sxb/QsUP2YecqKvuXJPidja/6vC7RMZnn8/9us
4Q97ShvI+ZSwV/kYoK0TiEz3mnyIZKrMECyKV8hcrVlv+VgWoIIRYgZP0rigt2zGf6AA3kSCiItV
yYNXssUn0t7qj6LN05d+HY4H1Dc3EXkO00sMqoesVvUaL4jiR4e14jGceH0RUy3XStPowsnrkTks
RV3YDrzc58NFxNd5tJAyLIG95+VXDIbe5VBslyuLSjMIR8TrzQUdS5xymoG8W1UV6S52eC+G4Rqn
ABhlotAzluy2g4G9Uv7Vyxp+RxluB8FziysI873T1DqXryd+SHbZyvxct48dvuNUyrZJhHKMLJ/w
40Qejiz1IV0sofoXoh6a/lNvYgh5YdmWOm/Zy/9H49Ozn9lHqyntEnxK48K1MNdKHKAsB2gbqKmU
rj04WQNXq8IcM8TW/y7R+xJ3NwjuRqbLsNjxtoRRkUir7kpeP85XLHC4WZn3rsnFVwGafgkh4Obz
Co237EKSZ+Xr6OMcpVamH3P2RzqVZDbpliJFPmgXjIaUfIsTjTbYdogEQpCaOU9Jnm1j0wrpyb6k
flxv4v0TMYI0WQspKAFS5HdgU7gya6eMcZvUEPHgIX0g/ny3CZc53knqPPgO/WxpwOFyOmrwuOX+
o/ZPSjFrD3M3H0HdGfLDOh1Err5AzxF7id1jqMxFLmfYqSdsuzXpgpstzhwMoh3NrHW40z8VOq05
5baGz6LE629rIv0NCPGJZr7MXx2NwI7bkTo1tmWG4HlzxY1OoPnyg5Ok4bRh7bmGD2ZIUhk4fWgU
M2+cTcM5U3sUIMTJVIEvX66eP1BMwXaMLck7hqClQeB9883wF/GZmcbDvBMSJtcXcnovQ3XnTLZt
TvwOeDGxyB9EBtK+UG3TZp7MDCAAwBNtwwfFfLUozVhViDhqp+oHZbAXKw0nsZJYYq5qfsVDDUOy
5aBQfexmH8SJ0RYFTnS64qw7P6UaNcHDkQm1NzU7EZglW/a2OlubtSRTUoTAyVTR7A9yP7PCQT5I
CE4kC0KZc/uTwUvswvoiDZPJgy01eKdAQWPv4LEA27azNVb5kIKogS7LOSw6Z+AZnTOVnS37aFSc
MgRAQhSR9y0xdBgIouXIyfqKAkrHAfiSqO/Ie9U2KAYsk2sxmbwPJPESztXhQBhuEhtpIwJCb+bZ
+K4UsBSLEUYRrsg+1DwkYPaUCeHz+e+dasgRmoKxAzKwBiH2Pf33dI4bAocb+6Zx1f5lb7W3IeMq
M65zd4raKPmHEDw+J2sd/WVnp8L7FHNCMHN1vCx0l4AZ4RobAFGeWx87DfnXB7tNuYp1Y2LH23o/
3/4vjzomrpanAGzcAFYzJ0X55WOi2TwJI0fk6xcXzs0EoWeqEF8y8/KYxjtKl9Mdmw7/Xj74ev+x
M2FKvK3L/2imTS7ibxKQjmOLfZvxVt2SpGAokIjfDm0LdwDtSZhe/4X4awss+qBmhKPp8n+Ui0Qg
os0WF4olKMuFXQB4hA5ETP5tvsR6TsCH8nUEngUMT3YDSQkL07AgTmOCuss2NEqEzJLVN7BcSJ2V
8nIlrIj/nAdKdq2q/mj9imx8Bq77aWBzbrCj4w1OY+Y4tTfK9F0HTFJNp8mN0rkq2/mKA3Dy3vDG
puTV9UORVMTnRFf6nkhLKqHLEI6KZhitDp7+Wk+UbokwO6csw3wdk5ve2J/6LqxOrLwF7LWlrl+E
tn+fPpOkJOdpqiLZFVHP5OzwCo0BvtGYiwx0OlB5qqJUtUOpt1VmEdwCaSW4Wf5Gm7il+w+vjfJu
tK3D7PDLkr+s6Yzbl/w3JPSdgbppdS6c7djuA9tk1dKsQv/pAThq/pXG5/+yb7q1INriJK0HQC05
5KNjOM2Bpf6arb9q8r+zAkpnoynVJ8N3/f1zONa+dwiYg/yVMgU4rWX8c6MKkgqBooiP827FzNEQ
SDe70kFYI7xrzyDLH6urPS9SvGoHVTZqxckPDWOSehnlS6jacODtvknx3a0TZ4Our35cf/mCb1IA
lhZgi/jhze8iHbhWuz7iFpg6tKvbrHHW7M5CCVI9q6NE1SlnEnqEkYFR86eoOtZtTJHY8A4RwMZP
1/nh2axW6L7DFbgv4ERVbizdjcPLQF+xgMcXFz5L+Z8NIfpdHFJyjcpfsMWPFeXLkW6INPEigeWu
M+Sey1JDAQcjZ77CYt7haU/YrBgvj/G+01U4Vbckgz5luzOjZgC5AT7c+QqSXUB8adoDRmsAjPy4
hO7LmFnooCilZzudro4/t1taMc4czPeh6ZzOtDNoRWO4UIn6H13ThmMjISLe62SNYhE360OoQ1pJ
e274CIfgV0nT88SYirxeGc9Cr3BrHSIF6uYYXZirzKFKqvn62Y1r1N3SyWIX+TSgVdu8uyFgWj+W
WayYSpaY72kzq5dDJGvAMivf9RswW7gnc/D736QalYHnBZZtkgo5tNEbsTlirTpJsWWFEc+inzAV
AydcWJYEEqZrNVkqBaGSdKUnLOy4i/noq4wzfibZk7PW85EGooNpsE0fdkHqUwpu4dtNtmLYY9Kg
bQWMFPAOU0i9CJs2NJbU1r7GK5bnFt2x6Do2itbknHO6MahChelXAT8ZoMgkXy15X6HaTadW41bm
39mLi3vKanFjMh6DdrgVto355Xmi2iTwXX9yEdFpRputaf2dICgeSw94V2SkmcGOz+/wvWxliBFj
9W0fM4tLc16drfvPMteJf0wZWpgLgcLaS4RdQbBcqvktFNPhzckKF/kaMocfzY4BVLxyN7Oapf8l
EU8XpQuEuv9YIk1JUmYwueYkIJcVhEZ+vVl6FGMG0qNQBZu7+FAsd5aBOLhcCCfsI4Lpu3T6XiaB
4hXUcnRbE2UVupVCrrufTmeki98q+sQgm3oU5Il6DJETqbIQgGKLS85R0LJlIWEkenUDlnKdrcow
bU+rEMrXBlE5EN1/zLeK1RVx8eEqBndVYN4dGcFTNyy6nuexM44cUAUROLYWJRb/4bG0niET8i3Z
gi1oEn0AET2wcfIgH3SarWYzrJs5uSum0NYAOHFnLsyvA4XWTt0f8ZdU+2UW/TDfATrC+y6ZNqtt
L774nU+X7JrOtL5/D1Rgh4HruJ+2WmujeuQiqre9+/EQVdXG4LQu0oFeClpfDEhF01k5cr4FCxOQ
+K0dejHIBHWk7TerqAmiqxAw1N68vgup/jMh0dOwRLYe8N02ABBMBZFgKVXoVUY+XCSysMyTfMh0
+5+SRObCoraSN4azuacMjrMeArkhNBo/h59pW7kaovHyarYMaXkISURfS4cpAeGaJYTF7ShDs/Pk
8masyedMwWtlv7+M/188OEuCmP4mEZLEXOOrWmy3DEPqBj1dQFO/uuPfB87Su/TlCoxfvKCU1trO
rnEfkhjLX2xEwHsKhrqwJac0V908/gB9zCavQRG0Z3PjRFSZNrpgOkiP13YgmHAufsU1EvWfMT+G
NUSsp1p1CqMEHVcYow9BL8GyRgVpS0yZxU7H1Y1EV20mQX1dU6UpaiNVmm8SvQjG23OWfBdiceRD
3Kxj4+wqLYVdEQTW8mtzXh6DgfAvPJefXloO0jZnoae/u33eA9OTtP1r2VMU6coUUJNDzQW/qcd+
qf96UGPfRx8NCF8ZxnGi9RSM2iqIyixsBZyqrcGudIo3jSfX2iUl/RLBLsRk3peyU9b73Aq0hkG5
5t3irIP9q5m9H946tEOLRR+CsjZPDxguLYJfxkc7C7EPkFJo4vW3pNblKdH+FIfVI4JgwF8VebO9
59BRMpSi+ObKiXou9QxM4oFsWetsGY4WLxRHNtmEvhjY+TSCRFmD5g7/Kj95ATUmt5LnCRJU7q1M
XukMbbVcy9ntP87o9TVZ8VsxRkd80ReXwQUpM3+yWEjLtka8Sk4RNKaKMoDs4D3Dv2nTLDCADmxW
PVtG8feSi9Ye+L8TZWX6PL8Zq7kSLcx/3vfU/tsgQ2GIVvfJt9GryiIFxUCSFcK7GzJAm9B+fJBq
64snvmIkxwFdXwAsq37mjfmOqgZvV1KOkMqtIpBTo3bVTCEkJVurXEZwchcr4fU5efbMNgCR6AlY
Z7kupHBcE7qOc7e1oexv4HyrtX1GA39w4u6R7PCZjRYHQA8o10tILhd3OR2rlX2I19k2tBrhT4Oc
Qi9MUmzsKeG7nD0FjIQaUIPiufatFFOtCLioWB/k5uerYycEfwtNqYNQcNCI9KJE3+ZfznF+z2Yi
gUkIg7uhsGCT0qxMhygfaDGrax7QstUvkSsyFDdosO/b/FYQeWFt4ZIVZ3i9icx1f2Nsg/28QONg
ySLCi/Bv273xwAZD8Ib2PxWKb+hPLarpjwwstRsdEHAuszk6xJR60OxscYZ+ihNRvstJyDQqJvVO
o97vWxATLFZNUZRtbB3i19hf4lubQXq3rH72DPJX/R27yYCvOWqUXc7AS5xGhVEepIzalCWF3HBP
21fJeg9cBZxPDfeEajK5oWfAB3VlrFLQMCDoq9V2tnpzhDmO7fDLonkQSdz8GaypkOF5CapAmev2
sG1m+pqugAHdgw/75HKdmI48Vo8G1Schq9QxbJHJrsP0RJK47ELpw5R/VbT3xVcU9O+yfipoCSd8
lcGPgeOQ+ocqoc9bgtZqVFkxs2B69rg5t+b8YAGayusv6BJgESOAL4PYhrJlNNuH/J2ie3ZKjiy/
nyle2TE3lAYuP154ZJtTL3Xq8i3R6aEKvGy9LEZFgNvbHee6jBIyTrjQahFCQ0eEcLaAcf0OVBFX
pa71Lr1unVeNxUeCGLlVB7+JKpfd5I8TXilYh+mziKsYPHWf5hll07/MhGno22xyJBxr5AH4DsMh
xsv5FBYTGsehMFkdKDAcFXmEg6LbxpOfzoxlb+2UAWyyM6zYXp0m5u3VpAYzkwMm5vUiKw48ivqR
poXZKYpu4iALW0r1kNX74S0coMnaIxwRw5OHUtCv/+owHRsEaxpb5C3A5ZaFtVxm0n94AYvP7+cc
69WrpoU1CRAc4SuyJtefjDOrreAizVSlfi71dSqbo+X6fVKYOXAs47BDcgO8F5LkYlg0JhnyzDPr
HGzPmyKaQIrWDaaYcqLNU0g2xU0FKNAEYHelqqzkjPLV3iO6JG3od1WGksOxp+RYRCOfB1l8wJEn
InNPjrCA2yjBL1DNiJJ8t9jbFcc53ZV+IW78H1JJTIC+nDnjexWum3kJe0IOKZqJsa6g4MuW/9jp
a1VXQpV/Ns9xbXuuxuRmeqWoIqdtyR41yuTKLH9X/oMz71dmNAtCACz+sazmdD0dMkgyP2YOhDwL
aGBPXnf2PeNLY3fgX91QXbFETfSB+60QP2C0d4B4DAeYeFpqei/ciJxkWWbXAqmYHlXnQNgzo6zQ
0biwUyEJQTWJF8ygZNtyEaSaxpFi1T6Kq5sfthj+F7g/hs15KrtHxB9lXzab6W/gE7J0SAIMJP83
3D0OdqXyF8TnMax0E1/MJY8cIP88jfcc1STcHrFxD1Ck51lTBH/NE/s2/mEGKkFPQuUCvPSN6gm5
BVeHRE0aiEqgCEmF5xtf9pAoV87D/S32s54oykxCmOeriDdoHHy8jtDNsnDCdyWK01jNXKKxd8NT
0ALJl3aXzvPoGppR+YClnCoZC/mIS+C1BCRuM5i78WF1hYh617M9baF3NK3ZrbJTzwJKp0zQHUy0
3S4LmeNTOEktWBax762gewUuCjBzYwU+DwDeoOkTe0TlXTyVATbXDZ4sSx0rUNlur+1aEHXvLweR
rVKPmYmV54TG915gUv0YNsqjuS/yvohDOOcIKNv7A2eNNhvBCVbFKWeez+LKeGEh3BCSfeySziCu
F9rc8NZw0in0JzeyGZE3lpo4YUdTEYij+byfzz90Mm5ciO2u2CJfmlEGBWFi3QhUwFllQ44ZZkIb
dUp9OyesksJfcUUimmQJf6xX2pCih5N2bNSLh8ma2SESGkxa1ZsN9jDPSEC7UxRkvB1PMBK3UI9D
UCwBKM3V/NIEjoDjI2IzP0M+Qhs61WGjtpuPsy8OJa3k4WLVAkaIe0c18BQdAxPHJsulQlpk/nza
J9eWGW3AVUKD/mAYqjJzWwsQqrE6uT0Pwqf2rQp9LiY/f3YSE3j9fUgNfnvxU5ybd4RjiJ+IFJ1p
z4QKn7xrDAG3WesThoMcIe3o8lDnKuZW9qR550wskPMDYJatBVB+cU8uCfK1IipXXGDKUj/ze8Mb
HwLsoEwTgOfYY6hKbZYpDru/5Gxb2a1agNvXBESmMdygiPBI0v7JZFTk53US7peeHEJwRfbyVDTh
K/zsKBWEeykKg1Ay6gWFPagNNf5N4u2PNyENp6VUKUI0Z4fIuv0bUPVT9SYDHwj3lVAuCW4jMkHZ
jAMcjvtCNdQnBjrJkUO/iayEeNXEkOxgTDYwvs1m81eMwH5ZVPgNYyfH395zYfo++jjMKeCpax8Y
dk1X58v7dzopwnQg9wAGjHd8yCvWguQh2wAfSRyxhMeqjmj21mKLzlPdMXBkEzyUJv1bSWgjDTka
hIj3lze2ayM0twlef6053uZ13IqTAfjcPMLf9IVF219JHi+LPdCNDeKUtM1mdDW8aZiMEQY7zkKO
c1j7vPQVOdUzLgo6bUJwpkJ4tpwLR8VmUc3ZXF/U6D+3UOxM2BdYM/K7m/u6oQzWVkQHfCBdj6lD
xFDO9ib6I+EHwsa7pslZPKJLrbWH0aNZqcwjCOQjGvzQGm6PeYo/hWZjLuMeurBT//0YvEbArzdw
CbK6ypGMicGog1LyA1qA0u+YC5bdgg/5233ECkc8Mqd+uLOzXUcV/yEFnQ013x+wGUiqnodWsBTz
J6QQgV1iPGVBVxwO2jFD4NpuTdhmixVbbDeUM5TXFmFbxFnQqkMMgunKr6YNMNcGZx3oHMp1vAEN
FM6rIOOG7f2fkxPmvDTgx7KHFvl4l7RYgsxrtreofFGPc2MucCE0bBr/2frAOhmx0BLvVKp8KClU
8qM35rNRURaxmBoekGpNhy8sKCy/cMnLbt/Ji0vd1JF/IJG3yibc4HrmnIc8xlDiiS/z00GtdjeS
SeGuvNCEIIewDwXYr5VLd/iWyZY2NK/HbIT3DCawUARQmOBmMqQJw1gtqADpDdbviaH/L8sIjkSW
Ndb3ub3gHEJ4QKgJG8d6Cf4EaAA1Fn2JAiVfTmoSemJezMCP8qnUR8YCYS37W+7KxAbUZXI0yIGO
15xcYoNO4rYBBVg2ypzBC94fLYxasi/aCF/sCYPE3ZX2ron8dxiU71APirCMeUbWWyQ/dU7zZp8M
+Q28yT+27juwZaeKWPBtQNSc6HPLAKw2v5sohMtvF+ua+qYu2R3Xlw4rRLi9o1nV7Se8bCsy9JOH
H9u3YNvmbykCs+cwy6yKmJeevto+8L43PysjtC2JeRLEdb1TsVVBGndSfIxaqhG7ln9GivMTJZ0U
rWYO89ixd6psiXMctpQGhpGjV75ApkcKGzBnBSsWrVntDFJtQIE0HqVsszbmhChplsS+8dl2m2wi
RpLLaD7kC0Fy4eghuvjOwqsGzM4ssYxNzRX+ijGNtTb1XZaz2j/bubBg1AJXDpkSNxeE4QDlFJfB
TVSdVHpdvB/GsENrS3aRZoC9AaagQrsL9cOyWfWVeMumb6qA9whnLNC9WqKRjGJlVQ6pm3pFaRW8
pJWc0z/GLNgK9iA0X+bCClsfcDKvTfkKZ7LDC0zoNMI0r0Lz+90Naf9idL4LndT3rYGau46QGBWW
RSrpRjIi+p1dWGc25YYwvhK67JAIV7mVCb44pYmEBBj94o81f72SaL7jOUybnhEbAGcm3ogK40Tf
ZUWkbVA9t7VzeMZx/kiBgBeQOTionnL8yYMIDjhaffEuOh8Dni8eyPcfwbqKPC6uCOXKysWNGHaz
zqjgTLs+1hw5BU5ZaagBWue94FO+NYPE7EHy2xj54J8XStueVRPFAr6Nrglst89c2JzEa1CF4Dui
QEQbMXqDtIniHhwvd84lKREhBt+/gUP4SCs58RdKnz9jSucoeHoTk/+Yo92zkh5C5P2+2bPwUAzf
vqhJoZpw3C/2Zyy5mqxfnLE8eJQ4Xeyw8j6ZdXtqkWWAvkyhVp3qgEA8sdIhSSzrn99NJvC0+EJt
BRI7oc3mp/InIkZHhihK1+JK1EYXmVPVgYTK+8g51Pc+kHNp7qUVR5la0o5oz5rYaqPzPSonQHG1
DBk3VB7RQplEY1tYDSwLOikUqwgaHlgzssBkCGN0UFGF8qeaqMt5jsi65r2Z6VllTofCzFryccbn
YISNzTU/g+lWV3teIEgrunfRZZ+XTS8Tnpnb8CryyYGIAcbO9xgNJOnwmMHfC7C3BRWL/nrBsfHn
kZMcdIkEuthKYExUNQHt97uaB07lZTN2k3BcYNmQ0sLySXOb6fE3adbVQlq5fHAHlaoXctZLNwRP
EG1yHx6xmG55I2rHRbwO9Xs6kNHrxXW4LjfNuVd8ZBLRElZY6tPwCRjfCH8hzNG8YZWQsFSSoN07
s644BZ0m1R4WpC56vqHsNxCDAMXUyB9b+59WAVmTeP9IC3XyIkNVebgAPM9dOyM/jFs7UxRMuTmr
0Heyd5ZISece2W8FbTnq34BZHEuwCjLdhO5Olw5efFQxcKfBUgucIWU7wwUuq1CD5NUaotl6JDcR
90nWYk5MiRnfS/f6f8vZzSt57u5L5F5jOHcizBpepzWoKYizShWzXqiutkYq9EjdlTKjubMW+MAX
XBopRFxNvES32stVccfx3LyiuIial/vXDr4LWITRjLNkgVqb1+IABM2E5OvrWRYyGmPfTwmEiW3c
W5c7jYydr2VgMnUD0SuosXTNr1dMTcS+CFCOyvdbk1RMrVLvvwLQ0+liwlMt3fU2pEkRmLbfhG9s
KLH20yvbZEi9rkkbujqTytptsYsr/8KmTbDKjpovbWq3Sdlij47s37z9b5FP9EPOmFvRtDAtVYeq
IcWH893uJ1HyjQsGkDvB7fWQ0ZnGvtkQe65psRmvuxb+5yzeYoy8F1YHwwCdEXqueo1tzis0ZruI
CYrKYXsnH+FwgLzARMSLA44xDR0rWMlo8NGAIFl4alBhXAD3gWznVGxE38Xwbd3ypi915Oh3MUQ5
h3EB+mUb1XXWCqxK0dhvH4JY4CBdVWOE02ixN2RMOg/J38mla/cVfeHUYYrJuamHC5dVcMQe0BZU
ioer7qPzETOGOiy6Cm2TrxEolp8SaaD3+z5aHoJ3zKKUk73PdrwzrD5vfB/ls07OD3oXPhmuxU3T
szJr3YtFU0tJ8wJfJMyzDZMODXmK5ITO3H9lJkDi6wZAnkgmWeyzXwtpIK3eheBgAESSIAndaIuG
pbQOCsLlSZk00vI0ReYz1oyl/DdS69tWgMFJPynXMNu+0geTFRnfwFvThI/A57ZfzRQeW9KJmknu
cj6q3lG+VRp9K4lQUiXc/Uc61RMabePkjldnR9dV85wXC5oTTrDLY8ir9dNvY/fIi8zqnVRGaBbE
uW68S83iVP4hV8iCes5QN247iV+FO03lU6R8MxsxnCCxjjXY1zuMr+goH/ZYDaAU7BrsVAgj67xK
vr6p+nHSfZTtjt2kw3vcB18DToWByvKmwcZWanl3tM6EeFkZCFeEcly6INSZSZLiIB5IWkCS9LDj
dRLymHQFuEY/qk7VzsG+NCheCUZ12NLb3ohNfA30Sk16WvyXOFc5Y2wSZs7VOKtx4gEsOY8N0T5W
wr0zTbhDHkoUpzimg9CsMtQQMXC1g6rxjE5w61nkkBs/F0dJ/Qb9GYN5gawxMz4B4LhKMaonA/1E
1xlmTi4s7Q9MiRqJmh9FxIsjBJnat8mGNVPKnLTmbR6AraLZZkGqehqewfELHml74YNVzWKpEYPf
qTcWn/bFWk7BJXRZX1ecRyz+67tgV7gLnvTNRn3OX5vjTwCsuUFYDtMDCCeQFfYPeiN7roYW1mIX
IC59jrLGQkTljBRxPMR/G2kGoWqiI6Qc85+MgXvJalEcP4TSZUc5eZeVbbHmVez+5V5YC+lsAGKR
xil4BX3/+XO6fh/JOxabuJqBmvo3opN3eiCgyUBnQt3qeGBLwHTb7izqpu7UeUGYeqcqVtSI7Epl
iYI4JrKPujEzw0h3NOd5ANRyn3NwerfLgTWlMXSD+1rbNCiwLi1Vz54dHZMB0QAr13rIkZR75P3k
mC50KvPTyS+S95lXpFCcYY7mJYoEI0xCyjTBiZBTT6rF6mo6fbI+kXVxRmyRA0IqiZFkj9sZx1x5
Wg5TerCfuTcRLPhh8V9/kTP4B/vfWrvnIyZswUVwD59Iv4uN/0fW+olZS2ctunQIK+AT7vYM2MEu
AxCe3IR5FZxe6MI7L6REQ0bqa/I4v+eOAQPO0jE4vON1jIlrj3ouKx618OqKeXDn8HUE/l31JB16
VWnV5ZpJVj8HcquaGtzwTrq886Cf7h4Lb+9lwXclLa9nsZtTvD9R1dG2bcHNAFXdGDG47BpmRyDC
0Ya9wsNGQ6NFKRY/BbKr2dgdRG4ysekcVSL1XT1C43FLWTt7CkmJ5ZL4Z7dgR1kn5mKbBSOSXdLU
GvsQuszFSCEuHy96qfJF7WausvXk6m+TQjoR74sJY3I0aRVHAgwbGukfyFnmonYz5HKFkK3Royj9
t/o4WJ6Dd76atDKwBvgG2yjzURnKMja0CgySvFFi9g0+Wiw8G0svmAGp8+4Vr6Hz+c/KVWtHJzDG
XaEGUk5YXOl1PctOulRTYzcIMoMWtPuW4dCGrwftfxwap9i6U+uxnfs/fbVuekv6EU5tZL6NUH78
3XCKBHt7effxBsDkXKXQaiPP4WUrJsHD2uNH3Seh86bXIXAnF4MPnsYeP4EL2bdbiLlHtZEFR02+
i+g9aU0OdoRJ5nBO+kOHN6g/BDcNxC+YieYQweuaaUEWX85jJlbzsi5pT0Ix0ohiD9RJSbVSC2RA
qG8nv3jttzN0flZrbj7XrSbeLZ/KbRozIhgscLbS+Ikmws7XKiV0sit/oi80TNLarA4fOW7h7mZ7
AJaqkoZfK5S5MCc206AFb1qoiSp717mzYLuAqAR5kae09xodRfTYglPKF6FNMf4qXNNzRMATeLCg
/U1UnhXoct4BfWJ13AxljmX/IrRjmI9wnpegp/LFHtyG3EzJ4+6pWHb2yyiUJt7y+c5IVh2/fnv6
32Otww0reJGXtpaWc0joqBYBS4ARd3U9/nAZZin3/juf99D+a2tIQmtapXRU8mcVsmUhZzhmz93o
ujDB1K8Yd6/XMT3xjee0qsIoZf3mAbkBY6vsSx5Sv9UYegPRIt9cIPx75LQ0I3iyoITWztq6yNUK
HJY2ZYtuZkQqkpg/ZOSCeCLtNXbfwNq1L9A4gr1vFvX4Ww8z1dyC+aBdTAuIuFPxOXqXQpyFVEHe
63r8NwPs1GtRLUZJh2QB/SbjXPCxWd8wsorKtIY3PzNl7frcM2S3S5GM2ZJXK1HKVNJBDofxam9H
oa+BSCTW5Fa8D51+55JXIfGeATEblVJPV5y8wl+FwMjPe7YcsCJHMxlAT8RaWu3JfdKE5WZzXPH1
p/EYg8TkeKautjQkzJbUk3RXGH+AJfpEigkqbE1EHyX6cHAYOqjY5x5R7RFV0lYPPXsIPuLexxdz
D3BxB4DsUnPGLPPkATadHgXan/doSPtnPtguPvVTmj030tYPgRPzQhGYMpxXGsTFqfPLOtIzrgH9
a2TfOtmNrpnWrlaYH3Kd+xG0fPH4H1OuYCvmT316AAIyKy1DA+Hh9gOvgygG67u8AOJrFOjKCtkp
UGRviTq7dy1D5G6AWm6S+72TslW4DfFdNVl2v4VmZYAessogTYj7R8ANcgxGI73wwexUtU1Cs1/Y
nuhu97it4u73qQMidya4tSJhGw58pRpiR2RvIUFUbUaEbgFOl47z2Itk3HklnKabNpmORvby2Mrz
rM7qmbpkv1e+6k33Nn26aX1sBTVHb7GOypBgvD/8XGrKp9U9S4B8+DD4+WJODdvv7sC1/0ek4I6e
1dTpj9jpF4LWzvLVmsu7YtIpHXntUSIg1eukS1khPw4ve7KlSnlonJMQonkvOiIrWcTw3BESxczF
gKcs2b9vYrCKNbUeSFxCXPKqm5SG6a5rG31VnY1rs3lMQj40bEgBdMCMps+XloejvJXhiBZvGPuX
zyGnUfjDpmOY70xozErVPc4QeSfzCc5rLrT6zdCQpp8wgQ/hdR0E8ZCKpFqDzP/y8M9Wylq+QPJy
UuiVTBSXM5iM0LCZi3nRmt/QlJ2vQ81KjpYWQGIdf/Yh5gkx+ouguQUHjDfVDunvQAAmS16LXRh+
H1wZPqQU6crvw4b9Z9f5pIctcIw+GBGDGmdrRv3wKQWuIptLkJchqFdWlVPQJ9CmychsjSditYC4
Tz9ta6ZSrPfffVNv5lCfpouvBE8tvbtOmDVeUb1/nD6+ebXGwZS3axPYmdFLZxf6WU0p1PNHn8Ou
OYSFW+5XbJoHaq9UmS1b49PuTFhSQFys80qh4PSGLJu0SbkGUFrzSw5aGnTvfFTooSx4u4mmokdn
2Qa3ntgCS6JX6uY/VoyXnZmdNMM3r2dvwxUztS8gsPC+rY876t/FSjqTWwgM0b3+xJ5lLLN6KY7k
BWE8QSlzhOyGdpVWNtYaFOp9ZqFdQ9Skg/DMf4/ORJuqiBUFL7xA+wGxQoGU8DgYSOca7o9VDbdr
FoIQE1r4kJxZDu7nEjyU8HwD3U6N5hF/wX1wKF6jh1wvkM8EHR45WbmpqqoDBG4nrnzwiojQ1dxl
QkqAnS5t1e185ETr7y2adMD0MMdz6wnXZLkayeLeQ7DoHCegTZgt1xzmuPhvakOggdBQaJRPxIWa
puIHxGpYn5HaCqL95QkgfI3vCLyMpu0An5l3Ht3p1kcaBOj9JoP/TZV4j6u4wovlmgiX+CQ6kI5d
oGZHLS8RaAzoMcDvJ3pRufjZP2sV+gKAydBHwE2MZOaioRU2ddhgCoWlel+77htvvX9traps2MLY
XjK+biFzFFlGGyCJH2oLYOrRTi//3C1LRjMElGY4OnffxEuSKeeyifVtuJpjbU239sMkV9CVGrix
ubpU9S4FKTKal6wOkYSH6Y1f+ZA4YDrUwOViQythgDWpB9E+EELsiIsVIamHaDLUPHx5k4yAF9by
dKnbfhgNFm4owYGRA6pgRUHRizzDHP0xhM1f70CQlXzcIqYeRwsve3F3HBEUcEw1vkI52xXCKLpX
umWt+/ZccPTlh0HjsfO3Pm5V+oEqLZI+XbohGwZwyVJiGo+/8sSJyOAQdnpI1R5sqgxKSvNXVHMu
GleXTWsuqslYz48LE5Z/Hl96dWdgMeEO8J9Zz35V0PhbmQra/1Zzr0VJ9fFCoVZUWsxwtb7YGGbm
Vc7Dw5GYQU8vaEWx28BfW4YWqNNL69+NtUOdSlOclGL0N8OiNRAJXHllcxFkNrKW556fjH3oARI0
Q5BWH8IjpQOrZTyGANFR10l/JitoAIGcqfUcxMFFVfWuPSb+m3qvwwQrngoeUlGSJhhXEKkZ1CNz
cIyW2rKWaGXvuzlxif4ONGxYmVLV50skGz9MrBCO2xqyruAk3lTBXu68I5T/iuS2D+uADXgv+Y+g
qFoAPlP7RnC7sQyseqiWyXbCdIwNtdfrmHX6Wo4UQkTSQ6uLTSJd9dRBDT0/Cw3/k3eebzzLSOTl
s+RamOCI+NslNFF656VfSMVLE1HyfUC6t2JfYzUzC2Jbix6qBpiATSH5bc7+lj0cPnkwDGob2KPG
jdElgyNF7M+7elPbD6lNMmCIjHYUW5PvawSvja/bikZkWvo22lBfjs0GdPfCqbVCYgC4sFbPmTWt
hlrwt2rgsFt9Zs3mMiNy/wPz6EG2wOCli6fvJwTQ/oAlCERTRMEEXMIDvZXPUIp5ZL36c7zix2SK
s19sgymk9zXDbETVVtVbyYFivenGgOy8aFoFknnHtYvyn6Uxp56XcAx0g2y5XcfBYVMqMpidN4cK
ncZbreyn3KIdNwUI6JV2eq7xLi1TwbQcU24kFIpJhl1IYlC3a/j0fmLKFgZ71rjrckipocqquHVI
2lOKiBScPlHfzIBn+XLU1mpUInbNU5ePwY4rjLDYcF0kUpynOYIEnWmtcoslYHPy1orYV1lLW5q8
bwvlIsk5e8KyV3F2pQzTgSJ/U4CTmeNflb6zECmqa/BO7VOk4D7xzx7rd3sRk0VevBNVIk78/8b1
Q5O8gRAX9/HD6/luFtmW+mga2VaT1QR02qfOkp2AF8Owu8CJMXFnTbq43leBmMSrnKrdBRqjztUc
x7fBoKIBO2xrVEzAr7cqpwYhkiuqewbtVoQeX7CZbt3gKRo9nZKVBORd1tcxOaEwTb05vv0kTqof
FE+MEquVcDT9wJ+uAc/8+lExxADkjRBfXyLVX3w7qnjj5Aj1jYqiH6AaCRXfLNyh11rN0zMh83hj
Q+oFoFzLToRMjFVVDjS0wRXixMrZrvSGrWg6qDCNTObE/QexVR2ZMoVSbQ/+2RtSP4vTMJHBJmc4
j6eUWbOOEXuZRVexVJpJyhjk9dmuGXKkBH9bX/phlhQCwSZgXuk7BH8Km84qULn+8PkAooBJoPaE
qTfPjSu4Kx6zfXns1j8UZXVGBK4ZGrb6vvQUKvArQCd+JsttlIRN5EK4K3DhNPJiDzynt1YbZJMW
QMEwTN+ETnVu6BTOZJw1eSHAQgUxFQWVEJOJb/8TXAMrzSjxF42YpaLzpRRIdfkcBrD0IwWPjyrQ
aKk1jXvl5/y9ITf1xOdN/Y2R+mIt/fTQGr5Z3irXmx6FZVh5vN6h+Ce1eayj4dzrcmAqf4ssjZy0
/jCmHMBcJeqglXX7wcZZxuJitn5+U3uR41ykQEFk5Wznf2k7L8klc5DCGdobe/+XiqTUjg1RL427
GR7x1nb+gHfsr6RCp6yXYtUK0ARsJ6co9VfDngn9FiCynYR5sSBz+fCJzGRqONr7Ae4ZjLFQAIgO
7bPp1M3Bi1oOQlP13st70AgtXM7DJqA5UlMjXT9+kYuagiSWaYMW58UZ2B5fcsQCAifmeb8tV2wG
kVTgW5vfXhXMc/dysMiadiDAEwnQgVqY2nfyx1r7I7arGaFQ+BFwBNrxXazCi6XCy9+PSAYNnZOD
cmo5dOOBXVvkBZpnfEMLhkFv9QU70a99XMH+qmBYAlRcZQxp5YpkFvdjx31ekogyiF3tws9U02iW
WL06b/OSS1fbvNLdU6P2jBrRHMj0lRnJOj8GK4iCLGSQEjTplVUXY39Yzu25Pzf64I4L620rtMRX
mwKH6Yeyzt9x3ge0RR1OyWMJ9ixhHNzeqX7TG2vFCwH5gC+Al4vxpD7wJhRYRAuq+RP0+4kLNnDF
nkweRe+QPIoJhX4fyFTw7Zg50gCojFdLG5AYtniE5PME5aM6KxrQdjcK1n1y3duO5eZ5dXzhWVCI
tKlfyrM/+2Os4FmbPOcg/CU9EhMNvwpnAnuatGCx/d4m5vMvlD0yQIfc1jIhFyZgWVpiLT3Pw8Bo
ZmJAVzcXl0cKpyLW1/DS92oy/5qzH21Tw8hyEyrXlZjyDOdEEV/ESGwyHQ+a17UEWAz3iIbiZqlf
8yjciT00n6HY7LM/inhEVFA4h5CXFqldlKa/W7UsculDNIEJJbvL1Uuh+gCEOvm4DbSta4023PJy
mPEsupjRDJROiZKScWDrDKMV0GCi8s+R4PbnuvuT8X7qDQLSAyh0v2sdzufO0IRlmDUaYiHlgzZ1
9P2+/EaRhTgRsCYo4osGGiWi6LFlt9hEMM+xShCtGdnaULL94c7PKorC/ci0mq0NpIymRNdER7mj
vr1Rlb+yeWiZ6jCXCMphMRKw3mUkLLEzGgya+hMqXkq0R0+6whEa7JVHXIaOGt53i72wxz9yxgwM
BrXDZi5NskNrb7Vi9bgtYi7dXObcqxx40Y5eaeydVJWdnlWOrUjL0/zpJ38+xMPEmJn5r8IjwGtM
kPX7NLpRUvTU1v5NmScMWj4P2nyQkpstQw3MLIOFFNM4RcgsqAZnFTWlEmRmEZFdFUFRMvR0ytpm
6pygG8d5iEF5o11IOLCwKyzWWODQ0JA5xXkk27TbgRT6j/zJ7lSRqYSQd+6xtpFwRcWrWHCoi/J6
M3kh6roCu4JlFgTTa6MZW6zKfUWfNHQ9Oc3MZggRGQh8LvKsnwMkyD7uhdIn8SnaaDR/kAkAFAxV
S4FiKltOnG8QHUqVwNdhxQswzOerasFapLZ5e4wHFsxGbDQDrTTXtKCrRFOhkOIer9avzfXc6fok
wKQeXJh6Cgy6mGF89V9OnIQs+Yb32TP/mLWaGaFIgXKC8fjIpxeziFjsUCkOBhOZcYS6HuFh0EQT
nAzMC1JBSIyutNXrSIVscpUqbmRlKa0IvDyLCenBdCwQAkDmKb2IAXfZwVO6gjNR7mY73slJX4Gp
jJhzZEBLhqc5PMVcHjuqiOt44NlI2Sff69YIUc548LO5oEANOU99IepFYSmXk32kPGi1BUkto/uf
459Dommc8zWlF5tA6+ZFLTE3ASvxDWKOYq7T19e/Z+PN37f+IG9moCta6EMA74D/5J0WT58LWEE4
0O2NVb7AM3uO8rAARuGq85/+9S2Ap1qJZKxCV1vqvKyVuuyDEqGhjlHdg3hVJ+exOCvKfWduJBRp
espAym7vdcjjs/QQ96DueaUh7Zcvnd5138FY6V/S5wqurZdqBXS5hzQJLo4RkF02k0Ucv3sGwUDB
HOnsQjbtwv5wSLHs1bZjgdl3NooMEceN1xp2vpaCiJxqDxG7RGOA6TX0MDV6SzXlX1NZ4jU/80Jo
bCgmo3xftoaRxI9aV2COh1h/57KkS4My/nqTp6w7f9ii9XSG7Vuj5d16UeyvWsgXDl2vxKQQH2n3
Vy44L2jqVDgSlL8YVHZi6WLopvWTD+CXXgC6kPSsW5cQmKi4wXGOqda6FWC+rqUw+Udz/AFlIbHi
VTAXdfdWVMn1XglJ5m2GJ4aFcXKKmJTkH/NBYW0rHGO/x2c1gJnpm+N2oRfHpY135sUFIsEpoigs
KW95j88jqCZnw+RabmaiTkguKwhoTQAmyBSLCliSAiVt2TA+rCxZUgiqxhfqBNa0RbRIVM9R42Ah
aHb0V5MrkIHxu79MpMDY4Ib9z2MNjGB+PCctbjI9HXtBNhoa/acJK7cjf6oC0a2V1T0weyOipuqi
AAzzIc4WfyOyhG0rCUHhaUFvvd7ohBWqQeHgkIeDZmgIRimoC7SshfNFQxp92ii8JEcIJRVRbOIE
wIeAr6kUe8UICuVCxbskHFXROJwkYa2xP7dTOSe4K3sZFtRNUv+a9Mg3iYfpNqnkurOKWAOfIYmo
6weBo7dmBzvjuNEnwwUfCVXTGz5s77lA/TgVdigXo2lobvI3884ipjzNVoDt8ObSgVnxg6xIKIPU
0w5KQmIYI3KZtN6mkO3zTcJAv86lB7+5o8H25yIzA7IxJJ2u9/MJZHVnNks20sMWbHYacQo6Bosf
Nl/R6WqnFEOotrqyOJYqjnEBSjib582MpadmfhmpsawGq+BrNM9lXQlPwYl6zTdbXvaAXOqm7xPq
onDHydCTnBLfF+uvgy3XpK1Wens2IqbAvsXq0urdF8+57GJZU7Q0hjOpls1DG18AChK6qValxYYv
M8lkdzXlQuzClhMydHieM60wIJvQuFfBbfX61xUVh7k4aKz77avzzKVW3ZXAaR02ajgINI4U4BY5
BxkT4QrVo1smNZxl9O0YbGgerBOCWS8aCaAWJTo7jR2EGMrsp8MpanBUX5kxB3K0q4tW4Enxesr7
iRcO/2QHSb8e7KMS8WtldLkgxDafd9XemAlIdFCcywm1RjflyIYIwbgejl6PGIi4C99ijgPr8/yC
3Nhy5s9FWeh5BcUMXsJaXDbTcCvqpvCwJwEuITh2AGJJHMAL5RgVG1hR19/AD6q0itmAOIaQmsPB
fPV96gVvXHJwmV+3i6awUYDlPMrAxdZDu9b/EHkmidInc4TZ/ysF2duOe25qWLm8sTwaxzA+spPS
hvsNpqtlpYygaaSKT385aKyoFIsYKy7IdSeSdR/2C5q4E7ovkTYeO8Ph+LZOZTazpxTp6OBrulwO
KLsq8qI1vDlFmGVQH1becRmZfNx+CluYG58YgDM5pzP3nDQlUomrc8JZI+yMOIMDaMM7wtb2044S
O4Rq3sJFNRyVoLh6j86cNDV22JUqLuuDifBXO6Z7Pve8i9itRrendtgfGEGTda6hXfvCb+da4cwl
A6G3HuZe3vNj4vAFFgpNKshHFDkJMYuLNSWe7LdfP2Eq38QpX/jL8RvFyw6g1hPBr2GQ8CKSMeg0
9TLZZ72qxZBGcH6+umgt1heDntPbJL+zOZM33hb4s6XPZIy66VDwLl2qkbzDpx1LI7A7LrGjeI+P
S4wHYDO+LcmGIg5+tzIiF7T36N+9WXjF++h7KfHUk8EyiX5hbfkR4DwSUetkfxDjpX7S7BZpxSCN
OP+TA0MVukE8Jne9cYGd6eyrAjqrR5ASk8Ky7FzQsIdX/2VLh7hL9xomM53rgeUoI+ekPl0QrHWT
7kcVLmzKQ40e3SjGwE20gcGjinDWY1HHsCS72APwgwOrgj2wUcHPFWpu6H8bd7eQAFjFK90YNqVv
pB2CkBs2FdT3/qGnZtiLKg2etWpbdJml1V7Zf23e7KukrC+66tZLxDoAaDbD4Rbp+ThvKTUmnPim
gF82+iHV48AD2EJ1aSaCOCpmMqM/ISy9cmjAukEPfhqbDQkbGUDwCkj7O1EaVmLgDUQ/l0D7Tv9m
Vu/dFmzgbEP4VWSZSKlLdEyPKdWMnJDoewwd4H9urZshVk4q2okZwHZR5J0ly5sn9yT7tcPVzrSL
7gckujc8Cz+1F727xQKIEMmAK1h76phtLcDgvyH8FhnBCNs1sXYSlPDw9iZJcuvPscC7v3ucQelW
yQI2aCy97Dk4/7lLo+BGF15yIaUmvkvnUVMsEjLJwJbQN+/QrzxkoyB+G6cfoR+mYujj4/6P/XF7
hBLFlD2VwxRyfbjlTqBuG2Nw5cZDVof7b9V6XaPmgoDPmgFAkT8LjRKVLoSbXDJu9empRTipQZ10
d0XiX01sWj+LgRbZ7k/T9qp/drxNWSCIRMjuSDx01izMBigu46+ViEG9t/xh3ph7dJU9ikkDcjrI
g8HtfY/nQIQDIt5EfciKv2jj4alaoqH96DDnGEGqd/dLaesELT0KNdweHE6ex7kGxNBgNb/EwTl2
AAGj17Mbt7X7zoF/Kb0CHZtTB15ogyZpzvlvKCmIO8uJ0yH/xJyUJ7LIcWtkRYAEbJ26b3HJwXb3
xsta9C8/VSiMz1NYm3uvH1bYRZRcfWpJqFrNo10co3cw0PxMMm/SqeXN49f66bUrcaMkpWPQ+Xtv
yOj8qMX3MX/Iz1JMwF3DQSbz0bCsZxJulf48FbaaqEQvdG+5/KpiPV7/BLWghI28qXzC9dfn067u
3nRVe/lH0e0OnxI125NSGYzFZ2l/P9tELzcO9ScAELWF4JpAn7jCRLlCsxIVjwLUF+VC6vNgXj9P
qIquhAtVPayJbwICoy167LrFCHO55RCX0UhPp+2qz85+QEJs+rmwgnRA68jngCSDTAj0SqSW30l+
S32N44LvK+AP/Miv0cf5hpiGM2V2iKvAnf79vDCaiiz6rUk+mnOqX9xaWg7Ys1+87n/QvYvZycxt
DqSR5SFEFSAOUNTlwPbv5S4cydmc8sVyaaAeXQWAoK5obDKARGrVS0Ow0F+OdiWDC5/yIE+oIjuy
y0uHy8mtzPuzFOaSMj+rZGiQ9fvcd9AFNMdupPuoUjYOHudBqhiEo+7ow/XLJHe7DD868sYtC6YK
VFmL/kPdQxfrvlQ51n/1fuemmlXbvxx9mG8oQkSakHfKlOXs6b+E6CWRB+uhEwPpWANIGZjzcU3S
ij8kSviWSeKHKXOVS9GPaFXbCFFa9/pXySVQxG6ILazwHCYRbdSG4wCjQI1C8jRrxOjC69/0/Svo
p37ABXGuzWWvqZl14rsmySALvmI1ZGiD+McHid9AIH3VBxvYlEGsvAZaVlGeghtCbIu3Nv0EfChy
dDHQ9JLq5P8c61dbSXR5r1jLuoha5pwOnjJ4Mmpp9WyAt+gLAxGOtDL2rVhueqb6kfhtEp9F7yyi
g9In32sxaBKfalRGSD8HVs13NshzwjhYAZhMozjWq4l6vEk8aX/ZnCCEdsB3m4jPBrCrZqobhg0k
jyHXZ8XKrgCncbwDJQ0PL7JH9ODp3xyG53UfprCQ055sgqFhKAOM7/OsO5eJUbNPnakOzZU/Ghub
YQd3JMmEdDEuG1fDgqYFW/bAm8PTTq7mlEcmfLhauz2xUSLPQ6SrJYYXPgNwuJMDdzOp94iP4zs0
oGrsqnT1J+oRe8Eab7BHAOv2RLi3E+vy1VI91mN4HHduZdbm3Lg519oCveFPzWJdiX0//YpnJfbs
ihNaWdLyucXoUTQsZ4Ooyrlxp42PgTbtM2MDe90StBBPF4ouBnGrcvqggjRBusH/liAJz6/2o8eb
uxF1uKNyE8gNFk1IRRNAKl7lUOnbAwgnMf3ISrlhN2HFMcCYFIaxOev0iYTmUwGiYN8dqJOnvzis
wfD15FrZEgOjfAsoEARiMxz0atQPgMBV0kiW9JsktS93ENqtlwX14BbGFFCHvuqZjDfyfC9btM5l
ywFLt0KFapicCRuahhnmyeoIf7STjkGi2L+9/ZmD6B8KcjGQmGVi9SXSdRaWL6wPoUZofmb0JGWQ
9ngOxKrLyFwVq1uciiKaD7XwCx9xLOiErzSnHeH3q86vYh41zaO8Pf1koUTcoXtHZhVjAo89n6qG
o3qIvuCzMNDD8q2afQLVWG96tVNGfeaJSu+erm0YxpzEab2pMlszdhvo1jAdOOnh8SiT9aK6NY0y
k0ngLIw8GyR7/coC7jy7k88V0OORFyKq+f6xY8mwkj3nIaxlbRlQPiFxL1afq/ic/zn6l4UrQk7K
76NhqKn1TiSFhV+2QOtBXuawlLNycMUmih0G/BoaOp3KtCaE/rbceCPeNKZe13ex0Fwwvw4Ka2X3
BIXR+hp1SZ8ERPXqjFfjA50/FMHEMfAhsX1cqnjLS/zYqBkTFihp4I0sToVKgHgnxsUQXe5w8h6h
dWqJxWMkAXDa5pKShgGHj40dCpv2Xl/0TroYkIhhKqk1a0PrT2goeT1bc8SdHgOTkt48slCXVROo
UX8ABL3y5EejT533aZK9Z78sfLKRAAcLlTh+5vM83IL/MeKGLtjyG5Zlhj7V2iLfWHrK/eHeEVK/
LHCcWlvNmH2FwIBN9vNvKCPihYYQyPOKz+5KgvzUu2HEDVrwOUSXOCQy9ue2rXlPGU4ukI2q3Tst
YqJwPpFrRAubaBmDqxFKCWVmjWAOOIKMkaVIr48fv6TF9CNag0Rcjxfp+YaMqjCFV8crOuKIZbF3
dR3S2iwePfhW4I6ZhxmCdLcWuqc8zIkrtXE6LmfGx2Co0CWnfOhZ3Mipr3cOVzk2WbDVf1s0abDU
6SYeC9siG9iXS5o31oeQmTDJUf73YYP1442hDO7/p2oHcRG4KtAYouokVPFN9ZAUFVbIQjWufGUy
l03zHDplmvfR61yONyHPpPkQ/aCZ3hEMJDfKDPj9yMh6/DyDoDOdinj7grjW4y2xcMGQLjXwD/lc
XeUfHuHpWEhUkJ23vLsdhp51HpUkjixBkzcD4ELqIbrNnz3/Lr3dIRrSzSR7dUQVwMXRkIbBeeuM
r9WuJNiup/vCkFbc2/uOKimPDWAmkQd5xs7yd4Rd0qZL+BLKqE/EhgJjOq4KGkMegpL18lOLcflO
l1DkEBKacP/PnA/VnC3mHDRGvKK65psrgIvt2MTKqaCG66YzAW1WFGR9oLMakcrNovHYR79BYCkV
2x55tD4Qa62/O8vP3ZLuu1ffu8U73tRxnfn9nN6F1ARgELCLWHXFSWCqsx0TNkNx07mhiRFRt9Zh
aAICAEr8A3vILq8PzeZFvfKK+ZIVTA5rW0xkYbTQb1S9ytikZZsItrkCmBhHxN3ag20pBxx2inFq
fVsclCpwNct/jaHve2xUzN5Sdf54+Rkzu42Bj8HXUrdA0FwdsEOqMPxLqWgSevOnHG0Fk+rvnNFc
cW3GCdWn4bBWaA8SWUkBH7x6sr3pSL1FMvWJnAZpuQwDseeWy6oRvDhzEKa0rmwHESWxCtcoR3D9
5B0OX8KO8MCInqr4h2WJC2VauTmJf52LkQ0QhrRDatOHOtvbWj60KjteCCOgu1mYW53A1sdZVq5F
fc44Ptn3t9cDoJBkA/QPHOLu2/9UlRvGJZGpv6iO5hJp2NkUpaHVPGbXRbSAAzInrBAoWWJzLTVJ
03esh9PtmFCX3eiD+s3WGbQcnEvVECKsvOGmoVetFSaXzIYC2WTFa43KBvUAPHeqsyYv8BvGpHSN
05C7SQYhx8xJ5Yxyy3VhxjpM1J5TTt2w0XN8xo/eK+dcJeofg0h00vjSHlYpMQ4sQ2F3440m4qpQ
iIRxThMhhExC3VNDKg1cXYPWv4Ss5gT+xLfj11CTVdtmv1iqaV3N/zS42NlQANvVfJ4vNFmRqMUH
bpqo5TxHZPJOJwWsOft8ACLqob5bAhwjMlUw8skNOU0fdxLc3bA8RFj+aygg5rSHs9hiLXoKTGYm
OiHK0WDSjCRgBJOMPENPpOYqN2LxBFJ3qqwgKikxoD66Sx9Sv/6ZZp94t0ThrdySN2c/DjFP6yBR
v6kNci4bwz5PyMZrbkzD6F+6FXVGYuCngovhLlV4bogHzC5lFGzDdihtbk6TolmEPaVAZg86vI6o
4CLBzDD6sXhIX73FmBC3TQ4qYCedav1pyQUDyyIyWhAZZsTVQjI1p3/Cy3wy1ZX0vsvSfUcEaAXA
lbcBGDYeEZ2gcY6Tm7Q2zfmolL0ICnttV97ry4VrW8LpyYo+wlr3eu5rOft+VnzJEIbe+7IgyVxN
bX7VHoOLTjDJ/O/g+48aVUJOxdtXbm5pjVE/QKMORlrtfNw1CZHJvxsgGOgdlitnK5iON1rZX6Ta
EHhrhY/mESiZUMSKfMvxuQMT1yyIbnj6RLIoGL0jY0J3xp7j11o/L8OOGo2WCS2u6N51g/Folo1/
3g76Yx9Ux5CB0QIRbvhNyQl6k2Plym/WhmoaCxN+XQ6UkIFBmTBgG7L8GSH8fc19f0rISA34Wdck
30tkNRrMEsV7PW/rZkHU4MQ4OWFVcA3Hy0PKE8gbk4wpktrX6mcaIpvPJgy5urVw3tMN27vxJU+V
3oEV3K7BGfWtXi0SIM2smmf64tSa0hQRd//nQ3BHGhI0ymZrX9D2xevKyQMoxAxLIt74p/HL22la
NcKDRSrT+NKK+VNFLQrf7Wl3dk5C+I6E5dIXa4RsZKADShh5k9XMwny7M0FYv8vkReVYYylyjSWn
QVVk9V3fY74m8Q0oH8H4MDem3Bxl1d06EaFg1NI/R7Kq17GtGIdB03Nq84hrz/ibidYDeCCXVYvO
/RgELVxuQPjg5DKUbenG29ZyHWlbLgWg19XV+hqtBeE0a0FJS06Xr1LUAN77XjptMfb4TZ0FU+fE
9yiP/SaO5ATh/n8wWkxXZJCSi3Jxie0/FQOlsUgyvpYzTI7CcvXziEFEMn+WProWwYbVkDJbLSj9
F8DAMIU1wl6KnmsQCatVjT33BS//hWfDgA71ARlHmDo6HWE+5hbSjBQhUKn7KQhndCR/R2ikVBIZ
v+6Y6sG7OGiGBC+rz8CDdNLm6/8PGnLruPwMMDjYMQwFvnRv0vQv1+KiOWxRxSth8PqCKjwCQUg+
4PW8PVNhI2pG6FEW7TG7XJzU4ZWp3vAeDX3SdrJZHhFxn6+xwDvWpyz1SsdfPqqGqNNsmx88KYvi
9hZDwf1cN/Mex0QEzufP2PFKKu2jLqLTVyVSMiGLQYTJvb0P+MPImL1zFuWC7D0Ny9E/PeP2fYPk
Bfsgf7Qvi9UvC+wQJ4QYDcfbB+3zKbmA5fc+ac/EEUDXW/E+w7jWT5fVIATjI7krw0F+IJJsC3kf
M+VlPh48zdl2r1hW25svN34aXyCl2kI6HsYQDbUSV5oyC0jfbbiza2xMzfNCMwlLKpvwL7BJgJEJ
OxI/a8f3ndGETulsRdXRAQh5qRlO0UcW6EFixo3NNUQ68/CL6bj41Kfjz/aZ7hjkyPKyXrVCMsXh
K6M/tVfJB/q/Kaf5tiGSAzBJD6t4TbYcDoPTomBZ8Fnngwfy9CkjkwoesxYjaqOOta3m1rTsmzec
4RA4JRXWpkyACGWrTzHvMyRHUo1AW2jNRdGMjg6Yte3TyFoGC4BRS2Omzw1zJ46Hr9WSyzPU7jGU
laD9CKkUyI5dO61pGICE3yMdYa0XDWJIYCTwtquFVoQXbqIP+cMahw+cP9UeO6+P8Mi3kyNu4S2y
zDg2XE3j8gU4LpQ1X31G6+66rL11krBFRbnGAsuVxolmJdkCvCin7kr1MPyZbNwaNN3u8SkKgYrW
ZhSW44cI6GE895iueIYf6fWv3QxeOfY2K4HAG8a0YeaVms7w16Ifufe2OUaDaYSsFmmqDRVnM2ts
1StPkL3Z+LnEm0Sazb/1qt6OfvcAKDwJwpbudbwkCIsRELrAlWMzmOdWSkjIzlR74YYsZf2mm1Rf
rwmp3c72uadJ96DGHAAcrSdT+ylvEsNKZFKCr4HTf25e09zfW4NOykTskOyrbQOyxsPR3mjsgNu5
VTH7vKF58mEodWIoAYLsxFkvbKuQFhfKLVkjiyGHd8N3w3l9upHHm1esWP4aKYJMWH7V1NFpi8ot
PqzSjCbcxqoOASd9ZbROtVBpvqjV66g4Nspf+gcTQxVfQ4Hz4Q2HoCr12xdK9C8qttrD3mS3GPpH
Pzb8pPzBIADyzkj7gQ/YSMZ+LzioyR/PTIljcAnDbsM9Iq2ZTTtDFaNVfuU3T5nJCdw1Q6gHAHyQ
n3XIi+Kk5HMc6QK3CgSo1v7KJQ45IeP2c+pqb5ihyzt6xaEzLIgjtyJWibgPbG3la4r2XzV72d4R
UhSK709RIJO1EUAw/KeiRzQUAKCw7mFZKOHRVeeRbtXh94Mx8Quanfpr7SqbuLPTg+am08Jz+djM
/dwMxRIkNQIwjXxUVXbAKuWMnZtm3uobQN7R2bCAqV6Xzt1TZJFr9vh8qBGIcDHSlNTm2C/3pczU
8X21bho2sqLX7gbpymDZjrWyeQDtsZpSVPI6qF5oxtlM1fk8Sk/PiEsxqx8JzCIv1L+mID52ZDHH
bSrVE7eV4oj6jfa9IEo+aWBhh+i997iElzNzky/2PbSdeLBjIBoa65mT6bRIMI4/yVrXnZ2sn8cZ
unYMyjWXn7i8pTMJdHKUKmeWvuWTeolrZ0Yb99woYqXL1OuCTKIGoB7WGp6G4BkO6fceZtKk/Wyd
Kulselx0GPKPZPhzW4oEQQ2IyVO8FH9bamFxEWtCcIbZVaKONcS2myy8K70VGxbhE7wibb55DqQE
97sE2AA9jB/FKt/AIR7q+9LxfJbNAhgvO4cnvd7cEwzN64NZSiQairXfjxCjVAmvwBOV78vCaiUz
VHxyX8l1JfLET2D2WGsFwCV+YWlOIy1xltSgdkZM9LIZ15qw5jMXFH0ZXIrKJQwtLWNPMlP0TYOk
jw7ov+s7z5OLj74IKLpsTPM7nMJuk01n0AzJhGOZXmlNYyX3997hHSAih1NdyoiSNHc9dA4L796k
aevYVGrBT6OclF6wl1H7W4l/M92hPSIrQjFCY3ecYdjtKKegUlyNeeW0plFway/zkY7jzExX8LLq
tH26xSm+vUS97sXahMELVVh87y1bZ/jaup5GB12R0tvLpT6V/WwvFnBkkL8stJ0YOuNI4lLtGl/l
xt/kCisBPIlsIjw3yJ79UJ6GbBzKKq9i/Eialmxpp3JHBr588vifwuIj2eOUsAlxhzOutk10/Kyd
+v/mvjGgLAmn2qy7MMgiwIMO9jt73LPa6d5quqxnzWzQX83lWqQIM4qOiYq4DijpVwXtoEcgzIWb
M0vE1inkbLvWJrgxqSRWgAJJQTHHDNOC9X+RAGXKmWgymoTOwijcDUhjej0dE5/Cm0X9vGWcDkA6
YnLpqjiiWLliQczvZMZWMgTerdpfHEDBlRsQhsGzl7NdUgzEnDQ32XllOcxYeZhW3g0maHe3bUB5
z0Y2NPCaawLxHYjutsnWZgF3jm4V6gOGGgLkUH8uIxqDVWUQfosAvGRMbVFc+I8AFQOiYsBadazT
sDa73xKYvhdSNh/KbetpLepoEE9+xlaEqPPHRPWqnQy75Z/W7FgHY/ZhZXrLMA9HEMBa744ufE9c
+w+Nlm8nGoeXc+SItqIc1bhuSnYkra/qowdeGuAKB3SRz6l+RnA17/LUpU3u8neVrrkrpCbUGC+p
GaKm7dY7VlOXsJazOHn4RbNYp1fvO4CGXG0sJy4ghOKQFOraU35L1Ow5HyQjatYDqm88h8OxKrdu
fE9gWFAPawaUqPZVvvRXtv3RkTbJlQIbg8I3jiWXdZLtYfJF3Byw8z8j4KPDNcPaqNOPoAkj7StE
yScotPz3UQuhu1Mj14XRtxy9BFwuWIk5+IfReMGoNMtTbhtR8tashXqqwgtX6nNGda9OH7oodBTv
rawdJMY07rnFinCGcHyJPIyBK00RdWVOQlcogiLgivmyUwrKT+XVHXPolPLWvSC7c0scPwr7BpMy
YPQpYIYYts0iM13WO4bEkbckynZ5HoXh+JRxt2Nh5/oKz6x8RePnt4JGhtRKwxIMhxVNBfgNZHio
Av2WLgbV2MW/f0wDrNhkILrk2PP66B+xdsxkxxP8dKwiHtgZu4VCnZax7rLGyaQ9yUUtuYOUMoWQ
Jh5B5tH+U4GUmTG5nv+kQR1HTsWtGmeFNndQMlPf8B3xGNw1mMvdJJPfoAqAe5w3/yquTIG+OE04
8Seo6HWomfbFTyUszRVkx1+Db9mrjr2m5ZlyVKouQplQvMe1BxoD5O4Y9c2eGu5N02WT6nyCNXdm
Uq3OcqUh3G2G/YlVNEiXao8QV+AZhtdWjgPg8jHuvzGIU3qVJI/UMe3a6ew3E2Enw2/rZQyfPfBy
pulz0SEtG46RjWkS0YNQn4rDNxIAHvOX7SxZLwdhmaWZzqN2vIsYmymVYusmWz1k7gAgaWhbkR2I
q+v8m7jQiDqrRQxunwQtXqnL1Q8UVxdIADlRdiY9uC5BXxBcw/wehVZZtvaBQzDiu4M5DmhN1awx
XBamQ0R/HF+JIEDfZMZcPyyrIsK5e1WstcwpYgFho95Fd4QGyUQhMFW+11IHmNn7oDCFt5eDQRBp
rwwLO7puaKUnBv0fHmIuherNktCGdMSTNRUK6iX+EsFUQ9KhGjzWZ2VogtWJG34TL8zGCjmNYtaH
bc1ZcnNhC9c7TJ+2+AaQj1sn7Ac+2ITuNSfUfWh7NmB8fJIBUA0+xrYGf4k3AGupm3nSegTPjVy8
tlTdXblJn8JxlwwKhdAbo9wrTBHfKd+Nd+G82WzhY7zObJeYHIfJOUCgcA3bUGLvinsfU26byvp0
A2UUp1NARWYwIyI6wHi5mVcAw8FzuZrrsJW4+zrKMGJp49I+qd6gm+LWDxiNNHNn18CD6KVukp3A
MvgumgDKzDwVArJrn87dhq+GZEqooylQYBkvL+kWpVdZtq6hh/RMHInkOAAcrtNMM/3HCPKGLOtM
fgw08LnNOn94Rr4uS98fvARzaXEmkQ36OGNgiBhdDfuyJaNWIuC4vxn7TWTlDpaPbVXJhOqMFR3J
O3Sl7aoW/0/UtUZ3BHUEbCGXFa8j+TBkc7oac+5K0ImvGARDRFiI6vdIundIRgFCOkNOjP71rvFo
aS9zbLRcMx0Bvlg7e1AdrDSeRkMObeuhJSK1K6Cl3TrewkL+cPxFsUm5CwFwaGVJaBi5JWHJT3eu
9UiIk9GOlQW2eRmP4fSmd+eC+v8Bit50VKCUfRLj4TN1Cn7dHWPj4+QZiaYqJK9eus2PGZ8f504W
UAWx8Z6vcURVlCHebTDJtzRGlGowxvLVoIxCkWM6KZD/d+pQsr04LFNGXgo396i15FGw8JhNgVWL
gQGQ+PdRWcMx55E3DXh512iSCDKCoQ/+t5sI0V2k9tCwm132Zz/kTGe8+31SDbm5WR0qVWA1uDBf
P3ewjaHxzWOoVz7lMpNZbSM3uX7+tUxS2kuITja+kW93aKR0ciQtaoie1eJTuddM6E5RWXPDkYzF
iRtZ5dfQzV2cw8RTOXvdBp3TOqA462i1oVMm7FSRGgK65clMFsNFnIonRfkZBOIfWd6TRD9+Y+Gn
Z/SrtJarAjShpAv639FXtIA8KNaajTCNzIJ1DUEmykHoSgdyEpPJUD4b7fzrUD1EiUXUZoPvpGw8
Mp8BjPfjd78A8FBW7NCYDSoTfLhVC1m8oK0K9qJ8M8mc5Zuieww5BZJsrg5/S2ZvV9st9EB1hXmx
wkE8k+YpBIcXoyTkvTfI3ECNnb2AtHDbyAZr/cqBuf8ppocBizSKWEUv+4O/ZipPB4JJo2G6VCL6
bDafVNQROM4foUNIHSGJx09LkkPSuuzlz/Eho5iFLGRTIptuQvUDHcXQKaWzTbBeD8ALQTcul8au
X6GhFyO17ttvPHJTtKAomhXNN1HB1d3nW21YideQu7/UUYY9lV5SRbXdOosJqHXr43bp/9BUpMZV
pdfdNThynLSVmkKrIvOgIiJvEdYnZOcYVNFD0A93V88Xzk8uaTD0siFjWoPumuwIHzWRJtKbJ8gc
xFeOLBBn73SzWD8b9llF5JINXF64rFskWSTti8L4QzFbCAI3FfKDNSVKnCuaRCqTczcou3Azx/k6
/ntLg8oktIjgINVlqwskcKIvPTAvkXHFJOkUbIq3pyPjzwxo5niWhuexe5MrUZBKqaQi8sUYQokD
vlH2siR88vUYa2PoQ4Bub7h5VLOyqF3QGgdl3xr7TVnmpFBBZezR7NHRQSciDLpLsVK04NpgpCce
rHXlmp3aQUQn4PAJv1s1KSWfeo66br+NbaN4n/zAsVRz17SOUfI/fO8IsYUleX/jVo+7N3K0R+cf
cdXUK9H9sqbYe3kJUTSaoZkh3JQ8y+boDsDBHFnRr3bKMhAfZT1Ziu6EMb3NaJ4CHXyx42/qBr4L
XHOsykSN0ztv2VOHVwmLdmp5R3YpNGDrPXQKi6/KYzMjTP2LQ5AXGPkex6QZ0yaz74B0IV39eDwq
ruLDpnmK9NU3it6sby9F3mvHNknd4HWgtWUDgItask4ZIkEL+fI2Jdxhd+vubGisjve5k5G1i1Ci
3naxSh5oitD0sVuNYVrzsHBFN2uh9hIJejHY/boKkSFF/7HJWDcdeUmFQ6TYA6G7MLDao1SUrbwv
Mlbo2t2jNmzz2i865Ar8vtOKjkhsIKMAVd1iBsYxlT4el8t3z+CkSCayFdN7s37W5jCHHEREWao+
trssqA+XS0cDs3lmAruj6T4Aqd/VsrKAE7bLEQmQZEBvkPJ0amywDomzQ5j8iJA6xGiGsidYYZXJ
MPUDAVqCYNYQKtHHKQVFifzB8yfF+76K2DF2JN3jLvT+z8QQX14J+bdiRBlTRvChvX3QBHJnCmUg
cZAvHAEDcBMdzsFRC1cjTZzkZFVzxNrBQNAC8cJxq1RsiMUNjldlW301xRhuMItwWFfDvJW4suEN
HNCrfezY0yWZofv+DGS7Flq5K3LivtBPWlJd0R2VPrBmZysv+awdqSzsSYz4DaPfWNOFyx5rbted
yyd1qc7BrmIxssCnvkMXCVMbfr19NHG4uRZ7X2aZmd/V1x5ogx6tfnysrVIRvMRsCC1woiNNfEqG
zWU6/6y+RcN+gVJEjJaprZndYgQKLeGiJWFtgNmWOhTR7LtiZb9mlN86g3lLeWLium4HP+qy0W8X
50WCGQLodaJSlzVZXx9LwzOK++srsT4oU5DIvbavIJPK3fbjb8jpPBowXAW9AtSnJKI1HPZHYdfY
7EQxaxfwIwTK6ujL7ZUMog4pyVtiTTyn76mifwIYBEEUZKw/zF3y6Xb304cid6LJdH24J9BrttbT
Cae6xbIXaXJJCyOVz5sjJJV8sq8rAh1KbnjmEnwb+78y01lqq8xh/f4zOOeyy8MueOakOYnsDpg8
5lysdSCudmJzC1A7O3aCM78K1a2cXbQ7umvxzQeZaaBwj6JWFa+bp/UjhvVugzk57f2qdeHgQtUS
fFe/Y9npQlEjKgfZzup+kM/Of5m7LZlfen9Jh06wqQmh9Jh70NKaMu+C68r97smg1ZeYc2T80r/7
2ESasec8RjorkFezYyRGsWni0+nVcB3u5To63eHanIMtMQ7QsGohwzfQzM9ee3nhWGZlzGK4TAP3
XxqjSqyulFmRsKf+7fhyV1tyudL6r3ED0Z+C/6/rdl2HrHMGRlY8AYUbI8EIfa4Y6Fn0ih/hVyQ2
AqOlx6dz1nVcsUQV/B8t1uMl/15lU7NpM2CC05NZfkMFdHeZh4Q3hhm2yr+7RMMRrsgJiBW3BTmu
C7HKi5VxkQNr0IJzubP7R+0I6Zwk/UUyy58ZQBm5Z3v5GqsCBTEUQQKGkXqQdsDy9y4JdofWdy/S
bMphRgFwLpW0rwG7eJWr6m1JDt42ZXreq5BYNEcPTvea/9KaaetAssIb5W8wb8JtPrRHeN5ClWHc
ixIjSimBwpfDSXv0BYsrtNYK4Q40XCDQNKw8clXBffdCzw8mP1do1cxXj8O1n1RHwYH+M1ND70iB
UwSMdIxM/PexvS/VYCQh6Ov1xCSMNVo8tPBy9EEIKH5QgBjkvuCUxR/Xc42WeajqYs7XLs0m1H8/
rIBTLPfFr6LStlmKaCfAENSFV0CPrbDg2cCanTJBtyx3KequgcGTsCao9+nBI+Ix7EFKST2Bl6Rc
KlfAyLbo27aBQXY1Daz0fqpHmgKEMhDUdVMYD45M5vbwpg3p5xngRX2QwPjFQhmaZBkGCEVc+yio
bUrnYmn0BxbxXjJDebR9qtGWG8hGsQTs7miybjp3Lj//8OvVqVYyzHV0M4GF8W1eUlZl8MJN31CR
bsn8uDYiaQWa/bKcSoon5IDMd7VdR5AvoWGQPIGLLJGyQyI9MxAs9/7SH1aB/WxgDJBYfdqHPG7I
TaJ3nKN1r0GjJpI3/c4/CPR4tOXL2bSzSdJUPsf5mpJ/0Bi2lHHAq5wuOYranb4jy+Dcn5YFLB1C
NRUAb8eKL+xtFbr1mUtGv/LDCAt+aNKyp8inxBJtPD/NIywuFI78CFg0XWI7pJ1kheX5Inp2KugP
ue5cY36FnP2rzDC53csMOc07a5rVIZSBZSqiyHoFdAreOZ1XHOM6a9dmhmp2rE037OmEc+mZlWMV
FwRCpawhQtpgocRg4w4xjUVyCGhOaw2UCXKqpUKwSNO0Uq6EAuJ2bvCYZIl2DejvZNnTFDGwal7r
tIza8oMpRX/bHVevo7XAHtKPoaG+npdZcQPXziGCSmJQhOAEBbRJzQqb47m2Ho7wSvpdVFUOZblF
tIdcI5oK3VvKlK+Wjk2za6VN9DY1z44lIRc2Yruftbwd/FEqeVbs8kxHv4UeDLjtoW2i4P+QMYwK
FEpiCrgbN9hIsTcj3W93h2JeiTvF0VkQGaU6rGI5mIDgHgIhRY3hIRi7o0P6dKZYW8hi9pmPcn/3
AxORJK9TimWB9d5+4xca9OqtDVNHDbROoYYp1hk1InavpwMURDYyxQ47zowZ+JguNsRI1zra2SRQ
IklxMolg26frGFcVt6ifTp+O5tbxKJ8K7GvMzKkmm/d0uYKJ818nFsDZCmztCdZLDtQ2s12ouQCN
PNQEK0O54p20c3ZVCsnrFFPA5vPk1zLhty69J/V5GrRR2ww8YGQjPGSMAP5ZiCRqqws5okuuA1yx
yNiBvzozKBGnQAOKJW6DnJlXAOi+V3zZ2cuzQ6SAsLzs2xp8uefKu/JoW8RaiXwl3y18K4P6aVJO
RWahN/iZ50Uyzzxs130ziYZWdu82YXwFuXIOfDmWLrn9jsjBTlLwz1ZhCq+0Aabn+9pkERrBRjkj
vI9RqqKC0EwHPbP1YinFFEkWaI38+zl+y9pSQKO0/nPIWihi/7GB3b6vdftC06BeyAaiYL+LRyek
hZdfTJPPgaITL9hPGNFaXNMbsu2K3xiVIb6mTHck35eRqJudmWSW7XgflqvLCcsBdgeePR65WiFR
uhr455Zlsl4Vbrmku3qkJ+gUxBn0ER2QEtnPezu0kjGQj+kjpnJ/6zewBXAmoC/Fm67zbZ6mqxbE
nOgsTNraPkLqNoEcwcM6kiMQGu38fwtTXgZo1wdpVzT2aSlLyB9KoilwkrkVTsSl3ekkVe10UjEv
+sI6su29jdPMQ/8kzaKsTGspWdNA5P+yDq/lecIX0VteWxUDNn6XuAYeNYosIz1CRuLHfGZBZTno
CjXsHMffVh+GNR1s3T3sKgbSNAAJ+5z3xCsZ7HdSJ+prXtYwG1yu30nuvwpiAYw/InJdPMgeHQTE
Uq6WC1zmveuGLOuuMDzg/zXbm729YBLHTM+oUxeKJUimIRoNRNOVFJvE3nKACo+cJ3iP9KNr1p+M
zVyI1yEBYkPTTmjv7sTI59t74ejqwQdEYp+hUFfwr7mztewBMtYSFjq+UITuxPPJoQ7/033029Cn
M+UJm/Vn3atUvik701GKtca5+BRmXGySWdi2dJw8xabeK6JCh8rUk2Nzk+PSlDSdIat9CoTlt7Qt
tACNvNjCwxaaQSWItK0DWmdtlwOCDW664fwuzhSxwPlR3IZ0Y16wmhd9/yWQHq7c1vkLXza5HmXk
UBNAjqbbCmIqqYGFw/qBtlfkP7MCVpevwj1GJh3DwN9Sp7HWfq7Z/luubzU5NsB1EtpjEwziQEJL
kHtSm2G5zPdsZkBIjLZZn+4d7lfFo9xVo0F/2zIOKXzzF5ERR/NeWJNforAUo2g+FNJIZkWuAAcK
hlNPuyNVioBvYcOelwxjyl2pzu7BVpEK3kFyeNhK7k8vu2JfLm8TpSDri0zag1MuoiQuLx1GLU53
hkTtmfZKYRfzBlW/4DpR1E2HLRfZdV3oYcMKsK7+X1t1I2cy3OH1tANk0XiJ47t3jiMjXx7gVEfE
uwUCTNOiOcFTqq5gJXzSsKKU79JVCVtkUD5/tvO2z5QNWVdwN84a1K5PO5ZkQ6IePOUb/n6BtS8I
JQFDTVhEitYyYYohnscoBS2hHEVLR/btZ7R26VQOkN40aEn1esHtw7Ec6rxrR+KTXEn4w/9MrGiE
ctFcWbQ1rNzqU3M4WA3njH2sEYf8z2VOP37B6l07FZldo/wqwcDNnR1M4QwFLM2mngxWFqtfLNTQ
Ry9xqfkm2AYiPrmw0hM9hXsBp4pNg5j1ttmLkthFvSHEt23OwI9ECqKReKsXLwqoZQQqOO43x8A1
x1xRl6yaM97BrOwnZlAqV9HIEKcbMWrW81IE2MiBQxeqYdMSYbCB6Z3CJMqFVXJoZ23VNJ80rJ7y
fbeqIVClyB4QIJIbqprFwimTmjlkRc+dkeWMQ6OEeqo1a2ryLtzZOzFdIs7gew0UgvMr5Nfo+MPY
2g7csk8uIs3sjdlTEvGIK7OZ/jpTtblfuGPnd9NdNKEY527bP6lKH/TpqUW26pzsAUlWz/+OeHjK
JOysGBRdG0m00207E4I14FbZri4HSO6wQ8oeY+2kWiMfYoHTAppIBrKsYPoPCnwHn60C6Ncj7Kr+
jhOU3sBS8AsK73RGzEqOUSWsOURY2mdZlBgbE8VX34/wfdjeHjlsem0fw+VK6q0M0N1Ha2cfsGl8
n/667wNykn1UconwrdV098sjoyOBNpy8vEzQG5j+uroPZP3R3IqYOo70bXLpjRJUx8GOgWHP8cko
wuRwd3MtwwpNCKQR+DQ92FXy3ecZsuoBrEzm4uX3F1OOFBrDQhXmbDngsXdjGhww0XcZrps5gBXk
AkAYvVnQSd4pPbSwS7rNqK9HQoaMb6dB7nkMeshVmyvqVntehpSjKhT8Bg41r2sOkyg2c5qPvHFp
/i3daxqgM8IPyebkuZ6wFkGZKM5UmyHB9b/VnxnhK9CRz+YEw56zxz3pZjqSSDOKgLSraqpJOPBi
e5Q6QaajSsWs69J5XCs51KkbhMtweZhMR3TW3G5NJvx+a7vUGTLjJqlhIWi5S3BuRD10yaUv3SgQ
OzTfuS4j+RJryeal0n6D5Y9v5KTTZxC/bD+r7dHjKunrcyx+b26tCnB+DL5zdqSaYG9mZHMw9ttN
yRhTr/9QsrkXvLy4ZE+s0mnPSTrZ9YxA7ryZxaIY6BuU/XeYDuFRQBJO4zDpV3FIlizB9n6oj0fL
0hw6QZdOPrIB4Oi6kT+hINtM8B5OFhb4CKBtErFt6XbrlNlo/5qiqIhKiYBMst1PMGOCCL+r9icv
WmGE4Kg6qUo2A+TE41oN41Z1EkLG004qzDvCc2r8hhDQaDpGZans9kf/VX1zxWq4wjGTmfQlSXqS
D9VCrSxF1xg1ZVA55skhkqpejN7OgacFsHqV7tJPeHNrr0odjfosBElokKADfU/w4k4UKYk4uHnV
OkmET7vsQjHeFtuMx8KDvbgVlh4UVAOIc08eFlI+9lPhXYOx6rVmkGPYLh1LsG9KtQ1kLyrZPplQ
VoitEC50xXdjZFs0UPeXATcqAoUlfvAT2MTUuSF34EzsYHkeqDozT3EFnRO4ZlS+5UtVCRVedTjx
Kok5BaU2QP9qdwdK1dUr/Yy9t9PJ7FhskUmeaNQXt9JMfY4ONduFIYEk749ewD1qHhyi2TVik895
QR6cos5cHu6C8Z6El3OzShsprmqfT1g7GE8LRQYLAawf904he5ixwdKvhgSf7md08eQjHRh6Plp/
MJT5+U3+QoJ+bRoTIbwnSTUjXCtVo2DxBjLJ++dZMyLACrGLRvrU7WzhztJckPDT2EjXYgreSGYj
oW7jsYLvGoz8TIOLlC9GdkFJDDSXXBJ3TQz9MkBDRaOUhpEJPTfmc2Qiso7krNK0vmA4izLt5+A0
Dv12Bve6qMR8A6HWw/WRGhH3ffHf1II7uHatYErnaDktiH0TlqcxMUuCABhgubPgowgq3cYRZSmX
PeFDFoy9jkeMOYAhLGsH1PXuAtnRI/XkUXDbyh811VOoF70FaaskeDr28DK+6X7JisxChWPNMkY1
dZEJZxqRBrGRZBLxDHzhD+/9p0b8m+6Wnv/mCdMSVdbNuAWvBoLkl8b0Y+9DK5ug5JdAkGz2+s8r
nB1udCcSXEEmMS6PJpD2RUl6SgHOOpdwbdfzWhTNbq0qTQvGY90qDJqqWLNdBCxxdhe659hqs5nr
Q95czsRGTJ0mmJfWeYeSeqURdDvmMRGRvOQwn0Un3VDv2lz0EnDkBnNd3gS4bYfelPeibXzI33wP
dMCUZabYn+wG9XfIE6pGPhNfBiDwd8czQGfMVvrrMRImsFvqQQ+Xz1klYxGjnUG51SopFO3UHKj5
B6Nz+xxgdcYLIur+0YavHfd8TnhQOZuIisWN8Fh3RWHdghikN+r7A5Vf0pV0x8UTUl724PYdLwnT
pjKngbZ1zASPtnGV6IvXWEp3/6ddIwsYC+f++jMnJf9UISrkJdEAph70FOHTUqV2+djnjTMyDfGa
zeYd8HUhtKnQOWJUd2Nom/MgI/1SMNtYZV0QupxSQ22MwfJjpQWEGnYTs0CLo+3rLeLFC5B1UtKd
DIHUmviM+U6I7l5DuRsXZ973S3tlVka8Ia0hfrh9YNq4Axq/0s48Mi6cL5VxJ8l8Tuw0JuRnb5wb
6LAj1SlnaD7iA6louBjjpH+nktCUMyX07uJw4JqNUsKuLgYF7s1lFAE/jc4K/rNpAFzhVsXj/eE0
voRKFn0qptk/hB8fgtym+7s9dP6H5i4pl4aDpchxs9V/iT+/g5IuVcO3oq8rEaaFlN1Ch86dzr+l
vChNMPBq2IB3lm19aEhs+3BRl4/eiSQpaoq9R3g+ZTZJuTI6ShCS1V+lJLGOAtojo6+Cobo6rH51
vAIU5uN1tgYnEI6+cGXz0d0r5lSkAOhPrq1y3ZTwJxd4+1B/2ap3oMy2Io0P5Ek+84ymbYx/W6Kv
YujqLVjLWVAI3wl0uZJXlzsVw3/zQLx+XdBMIzsxz/052thMn1UDP/robocEzezDApiJTFDMclbX
iBSi1Aoki/ut7DMjBAVTb5Ejc2K/X1B+1NbIjum6BG/68uSE2G1RZoj3Loowh5vuWRWitIMXBjRk
lPj6/Sj5u3C4j6aXB48hCJqdfWasHgGdDtj81kPXyKcEBQMKEqGRbodLEODplTnIYCGuRAqlR1Xc
gmVkxgRdUebJGV+JVuIRmPv16+V3qZk+etrO22NHpGjuqZBv40V/dA9RXzOif6T59uBcmqkRGftA
rYgvDrkdamLsLf1YhfM3nKU9JcLtYtrQVGcHihMhPr3Vly/8Us6CEkhg8INbCi5Xy6K2q+YDT6PE
7Y0fZ10ydHnKvH3QMtKRb0muh7UtLauWyhNaNyxQ4Ft6K3ODqTQdiFi1k/KJQqbkaraddbHHRBWu
PMWrHlIunn7Hv9Ee0AfXHKESX2ei1zY7taJ3UpmMACJW0GWqtZnZwkHJgax0ffUeN5nJp8LIBkXh
PPMbJuq1dorZxQc3ksi+Rd6V6/Mi/9OFh48jTR27MoaViqjsS+9XwqjII0Btr52Ehpc/VK3Xl+uJ
EJfgubw2Eoq/VZTA1iQ1EYOWWOkeBzNf3GpScjKtzi07o1v17qQ6B/LCwnnLBHeZPuv/X3p9Bf+6
sJNPjDHTwUsXSIyR4bpNj1TiHbc2RDkRt4RYdsrzOsT1CbIzC/M3MgoJ388sOxpWLs7ex3v2QMA5
5NQs1tG4ysnRibNaaZ1Hge6UD5Z9KsAycp0hZ2mmWp/arO6Qe8OO+zJ6TLKAjkEW8gdrQavaYkPb
hzGmpXFFmuiedHt3xnYVZnofz3unYdT2LJ+CyW26n9qb3y7xedcH7ByKsBDqq9JEGT5cGYclMe0d
73b3peGFgW1cTFC9dPBCEpRQ8+IRuPS92dgXNMJWXyQIbs3sTgVoO6l/uSuCKQ/bJ9pUZXQCKkUa
F2uSu2377QJTWISHYWMawLqJ1pT5gWl3/ZNUXZAeYyQbdHJZvgvuYChENcq3sz/cig8EP24R8rY1
4WBwm+U4QlUnvHsgtoVRGYqLLpqYcsXlz/99u4sfKPlfy3mJx4iV7CSGk8Kj0pSg/3tW9299Sd2j
upJunZ7QH5P/rCF2ZMra6Fbc2JTznlDAGlaHN2wol17rOj3cGdI7XXbQi60uwUBqjJwayoim/ZBa
22Nl7UXnWJYqMdWmH01Tnn7olt/bQDf1AOj/QNrIrRba1ABUmzxQ7WShX1/lPxnNd1003FKe3hT4
ZNRMoWqYV78fHRnsU9T/JS3JUveUZU65rrud6OYCYudR5wNuTMc0BmnvYZ+nYywUtSWLkTZlQ/cX
gj0bEU1+AlpTuBxCHOYdOPRz2zJahi7IWRg3Bj9ofivVsOtPKKP2sqjqMLu2z9YhuResNe5JgsRp
LopVzosNgrIUhoY61gh3ku8z/4mP9yPy3snkiuqxFmrpIShzIV4jhH7nDH0c6iVVfTkJ3KVs/hQO
OOo5ddi8t//xZP/KPcS2LHGOlp78+n7XRgi29aCFtfkprPuG9qnk7qd7qC2M/VExHq/0rVxoJnh3
muthODmGJJVaXt4iGZz19hj4Ut0RMTtyAGHTnX9kEAhrUkTfMJ+b/Pu7bMHEszHt/ptDmSAtTgiN
PKQt+jTQaWpA9qmz34NiCx82hwWoN4NW5VYDWkH/wbYcux4zEwZYczEtEZnPjUz3TxQaRdEe+EfV
yRssQVVazvKJj55R2z5/twtw0cmDAjkrR4YectuenBsO4Yh7lcGtoThMmH/jr5AtHj5HkbkBNI49
3je/tZkh48ZH39kySH5EmLv1fmyXHwK7dhgPrfieG/zPJXISUqUadpPR+kAedxDo5dnuHKGghcPp
2Mw7FdvhpTdhN7JblYOCN6krZtZ0rzvWgiuvdcpqLrM2oW3gHBhjL/yc0Y1EEG+5/JGmF5y7YJsH
tclktWYtZh6PyrDX2eWCSxx6aLrKZQn6ZbTbnRlr8bNMimuXTUw6YFdA4YoBPlLKLWDY98kzkFhK
/e2I8LmnfKV9i7gQ/N7jLGI33UrG7YJZnRh6iG88GZOL7BJRcYccC1zV8AGYNMz7CSWhLoRkQL74
itk0TYAGFbGatB5gVqEIjF/HxNpUXC0+07yrRpYQolFnopT4annfxujVITydjNI63Qk+C2QCYP/l
DV/+q9M34aXBJToAhqvMHxoq+02wK48DO627kjwXpGpMfRgerWIzrVOpcVZFP3fqwt3WbIJ906Mj
wKpX4r1reAqMyZwcau4TimETh1L9DF75gz40mudbVQUCR5eCPYizl2Vp9nCNus9uy7lU+F9WAw+u
Ax07NzpjFNtFHIkyNygommCfOHhjvPA5QYde+w6H05jxgDjqe3uHfh2YNExcUb+lkphB/AKD8o03
zNkTTMFWnskBEJru2gqWx6i1sC7zcxLgqXg8uqv2vWU0uYYFJHzDwdqIu1k73Ls2z8ENMpLbM5vJ
KVtOSpTdhFu2UIl5MwnS+czrsuJjltjfxXT26mChJ3lgEyg83t6C4T+ToNCgmUszF/gztsiBecOr
+UPp2oVUhWkS2gGjnv6D2QjX2kK+lSbgt7s1IvoVnf2VYAceid0o8G8m2zK8kGlSqy0uVFzEy5O6
rZTXuqbPnf269SRp0QKX8wnWw9OH75N72XDnzOJAAqlNZrfnfs0q9u0jQfQPNIDHwZ2u+mlEbOzn
tmEBZExvkh3/2aMYUjsLuNlCJ9nDZNiNjNFAGWxDmcf05qNvUEfe0MblxgMOcBIK5XDdGGvm9GDz
p1jHUzd8jc9aVVN4cqcy57o6WwDNyt4Zdd/jNd5EYtjlWh4Z/o+LjotQU7TspkmkW9AUiKQ+Jijp
YPjv5rNnLP5aYUbJtpjqK2ItAwo7TSrLOSkmTmImwvX/hF9G5qSG3ZZXtgJvZMD2XuhIqvH3Ek8P
Mtuj990XHlt4aQRPMO0yp+m0GA0cfGCOns/dOGxTqHalFL8CM48kFbbkngYsthH2lRVTUt858vul
GqXXZzyjYGOjbUO27YK5cDh2Fh2nZ7U+qFRmS6s70sQlsZDVDQjbSvqpCwVp5/aBlctmvT47DoP0
w4CSNSzOxHaUJoxkJN0bg/lMcw9qHfryqHrqAQb5PFlvNIolXgQU3iywgiGyJQ6bm1V1d6DGpxrL
YzxIhB7qcjkMtw4N4xkqQEBU676EuFfU5yuh8bWNtLQV/sWt7wuPRUSG0nzk1OiDDUIwSfu70K2Y
Owy1VuVv0jjDAwUTlLsXgjQbJ1co67NquFrzBAFii8Yqx4L2eALlCt589pARN+oiQN/JfuTi83He
BlOhVkn0SjeAjgpqBC+Epum63PtAiBkaaSBk4ykf6OQtEoKelBNxV46dfcw0rH2sVY7YKjrDzIEj
CPTaJUxNjA/Aq936DtK9pk5rOFwNfBT2pjtW93g8tzsJ12dS655L6aQF29PaUZVqsq6pMUCueuoC
dt5yBE5NRlnhvifvXkipNMjNb2FDeP901Vd6CmJRH3MqfRX1vBvs43BwQhss59SG6EXy/b/I+Chv
Sq2mqpPHBqCA724eZsch4meo2KLhsnUO/NKEZItbCL21kh0OKhUXNQqSjNKEZ69RjVyNCtde1wki
QBe/McNn8dOD5eLVybPO2MTt5WgqIjQdGGLQJzUhNzeaN9I5635VBhuUYPrVNvSmFsxFMJ3vSTQ8
59X13JPAontYjQhWBvQfuF+WRsN6bX/lmzQSu6rCBrWi4Cj4g42qmJku9KTDBTj8V8lOrKGdZcVc
hOklM5lnnjsQfxSCBolK1nLH7XyBPt5bPUWZj6mfoq37PI+7Oc0TVwf57yWkgeBsGgx7Mygju2M1
yPwtakpdoH0YtTcwj3sCmMVTFaZmNrgIT/I5RmEnIuPt9KrTO/SLMjsOcsBxLcDOCEZJ+W3m5SIu
R2Ya6DyyO//KisZnAd9OWirkw3cB7q7Pfpx1W9XmAnUSiNc8SiUyOn9OJkDB/fug1akdVaNH4urr
pV2hMSBvBKaSC8GWdf2RJ/a19gSGQwl5fl3rEdc57qtY9ZSx5Tpj7Q7FWoKCUqDpNdS2lPPpknQ2
tbvj5lekCRsyx4d7c4rWleKSj4TJI//ol0QiyRlKK1e+resIAJfzOnMAP0PZSe8HqxmKx/H3YX3c
AopVg2LTwpxayJ2PC1mKWvY8B59oLFUu/KfZj8cVVHpXCFJsaUtq0y+nBh6JZFsGZCbxtgbWn6+D
D+HTcvnBXSZFSrlmxtBg3SMXSZA+hK2zADSq5qAzbG2n/KCiTjDfGJJFrCge7TeEH1A/PbJHmACD
GGPfthBXvzcaf7iwCY0mATL3S7q479cFisyx6jE6iTwV/Kt7sLwbjgg5n+N+dkK8N2KFnMAF43KW
PDp1XE4TiJfAk1FqQHlahqs3nhg01g8lnUvqXr0ah6lIJuqp17GkUBrdHk68FYccTVTW7UIlLq48
dwJ2+Jt8hnlmQ0ywRtn5x2WtVVmG25lLQM31EeJ+NXZSwCEvIswOjfQ9nORm7cXBDdFqkreoms9l
V5bq8sCrJkJ1QlxA/UfW1gdJhGjyO33IEErHImC1Iq8jQbh1axryMDlgA0OIdM4703y3oJjPHuOE
m5hX1bRN0r5Or9zJWVyrrDvUAyKepXYE82ts4PBrNrF704PRWd5au2nWXnjDAowR6cXL8npw87ct
jpS0EbVOYGp0CLB9dVJLnhSh/bqkgzaYmdb1Cn1eT0z0e/doIbYG5JEv8MfOk5Yw+qPugUvv9loB
a32qFtWbpVGTWcHTRm/VU7YomMKHh+rLMFDhViihzRXgOw26oKG60t7zN6amLNNyjbzX7FTmGUQz
qmVBBYNNtZBMl3+wu/B1oJ5QYyXXbtYzK+a9ZncJ4rW4Lh0cx7gBIDz5Dy137rh5cOuDMg6YNFSk
j5v55Gsna4jEO3DLASUQV6tFJ8/Z+4EL6sim8d4N/QPRcCk+YLomrdzDYdOc6+ukuyWWNoS4in32
7fh83ERpIz+7qg0/iDwrIV6mD/jR1wgX9rea/Zr2sF5TX5daxIpjXu7pGKG1xQ177Vj/Fdykq5ja
N98v2qUfUxhpjUsaA1O2Oe2m2jRfQkoVlZmzRxqw1R3/MwcIQLl2Euz41GOrC1OsXVbEP85G1DyQ
RG9KdSRMJmerZLDGYHwMdVxBVWj7dLVdvRH//VD64S5//5b9pvOWGQiuemaOyIc/gUXXB09VS+Q6
tboVy+0M8GdS0j0UdU9KRHmOmrHqs2AT7X7HMO0bwQF4OGRLh4JPDxK4bDaYA9da00ajY5NiPNJg
UvZKpoXiEOPP+ZgMuG7VhiuwR7/2B0Q6Q79W9OaQo3GDKa99aaxdPh91t2phCqeF6pxEk3dDfU+0
maxRvhNNs502107//RM2pkE09thaeO/Pn2TlXMgZHHoCAa6xy6cs5iu+9gWWkCIjo1JoEdW8007p
bweuP+m6tvfM8WMt61CHQx43un/OYKis1kTSNc4lh+Jeu+OjoGbuPq77N3z3/6wPQM+XW6/juv7r
nAuGmwmASN5HNOvosR0iignPd47f9H6XgDZQ9ZM+PzwnCnRFSbTuMN13herY6jtL8AUi2x4zqVjq
VcsGXPTFHh/Q4egKcArvJDZkyUEUe72RxesON9N4H7DAmHfitnqcKY/OjHG/1vozpwqhZ4L5FTnv
l2BMR+wmNkqusPj8OfYuyUSyPuhVRCpCwGeFCdpxxA9Sv1cLC110Nr1zhKERyTKBHHuhGVZtGPip
dK6LuB3c7JX+VUslyaHDU/b4BIq/NmBHZHwUDsJntPXHEuvc0pxNe9LycEsZjoJm5UbuQr1TbLTT
oXSXgiew9awZ5RjB2nxUR1aET8v3N9SOtN+jv9Ig5hkAqeqoOh4JmcayGHIp4ye+2k0Sq3Cvv1xP
y1Px1X18VXmr6IaFB9f9IZJPkoHx7nKBltdgWnlNTkKEfVKDGXFovvxsy1PvX9dQI5pELA5gh2SO
vm6caUra1P7AbtEmTfx5ONMsteGbvB7L2mg5fqMUfjGV/qzhEgfsUQZAyTRtA8XJwGF8wFlJfuUu
4SvWp9am7TPehRSQmTPP8g9/w0Q7BMU3x5M+4VNnx8qMZo2SMrIghi7DkHCMh+dBlzT0qyEc2PJG
Ii8I2RN3JMEzMrDk7nl7zOVVVWPK+pCgatd+HTxND+rjrgqnP5y7eKoq6s0cvlP6dMYftwMT4Ila
PHol3THYJBLzttr3R4XLvjuRoCgsWwLRD32CuldGna5f2CppMdQLL5Df5uJSKC1AkWiLMB8YJwFI
6c5Qh7XlFTvVTzEx6RFQdvX2rhvDG/aeJsfwUnlEGHlNUqnMNm/CC39VF08eN3Zd40Q3l0v0UALc
cUm1oodFdk53XvHmWvhGzhIWWUuk6KEJ60kTluclJC+nV/04slUNfzJgtAen7Xqfblqz4q4I+BTl
EXF7V3e3eDJuloIpKL8FIDJkJOyLegPbq1lHG5TlN9fKJyVAeqCIHaeKzhJHoE7i4n4aP9emrrAg
ZGoZV/SDK9xU6SOXVbN1DRm9icXjlRlWyQSCv2A66HUpLH/b+iPjXJEz5NkG2t0j8Xx/2BJjzpJf
jjl3NXsZ5kDnwiN4k/qJ4rnxMjUhS4JDxZ4rCdrJxM+NlM+lAjgRrSWbfZYe99akRGpLdx0V3iHX
r5UUN8e5UMH3/s01ZbVUR/ZMHOBh7g+UGcClfQpW0dYufHpXufX6WzHBy2sppky6w4ihYYYMHGHZ
AuzVS/ReDsLHYsJioYf/Sz1n3AV+AdZ6DAZh/A3/4gnN5zkpXpqnt40XrEwAW33WADCuNnmt71vb
cspuK/kvRrQp66far+XpgrhwA1tY6ii+rhTpy+KTBtJqsm1xH+Fney9gXf5JLluGGYQnkQmKJqAn
80taW1uS1uODTlHlKnGMG3ZVPypwGuF59DSTgkrPpBV50TaJ2Pktpzj1LGChtMSOiAPHEIuxxSfv
cLuY/BaPMN2gH7EToHsyF5Ed5OTVVOfN0Bfzpn94gcKIr/P7Q+RbCmaUKnhkEEn6Nu0QXQfJ6sQb
AeKqHquwMAp4fYMiQif1Cc2r4qeNxq8WO/2w5Yq7PZIKSdeQgPmwX4Fo2pJZYmzmDXDRrSIPdjAb
zCTQmZ823MWkaPv8FasPQsvMWXDrNsVh5Zt0Q6SYp3JpduPqmlOtadMRBJUN0QiCuCIk/vnyXO9g
X4NUfFYro+9wpgcN4g1RrMk9RqFpIfid4umtrcyEyKzlObEbLCClwnZm3mAhfFwdIoVdsrQE5671
shJ4CWJ/hPK1KXw+Bvm/eB8hTNfJ/oEXPJguk6w9CLGIuhXO9uhjfwrbgAaV5Re5yctiQ6R2XaRh
jCpueTQKCBZvChMvvqUYeYxxTJSRZWCfit369HJArbAvO5iJKLDlBLlXjhNkBd9eBz6D3jS/1mfm
frV/dmdkzNgxKwakQrILI5iB6WZfDUv4yeIK/QWWHCTy8oCGEKAnRpzgw3UgVMnm/QYvODVCdjfo
UJMnArVqRyb0ticx/23o3Jndd/m82dxnWBx7wMkhRfE8I28gaQesZLXTiVyEOhvVlPip2VupvFuY
BZu3bQDAGIEKF/8uXSBRhIDQ8GQEavWiAIC2xHp534rv7NkZJoPAHsKm1Aa/PBiwnp+QxCVv3OHn
v4TZut8d5rMX2hTFHPBPsMfb5FL75KmE0CyvMO6DF+cwzM2lCa5KEiTNyrR+Ck7kvoAlYVK37zdq
srelcqd1cpPaPekSpKPt4kqXCHGrPfU6wZSKbUCZ9SpsWyyBRPgMs3QG4VpP3y+k1CBiOTowQzli
rScUFscZKzmpbMFPdT8Sc3rCZQx4wXX9GTrLj8arjKNlvIp0eVvI+Go95npy1YfwOIPYVnoEwiXO
HTyVBzjs4YxHV7fgDLCzbg6Ld1gtiueB92T8t+df0IYtbS2gRBVR/ObVdFLan5IvduVs4xwebfu6
Mge8qRyNVKrXoR0XbvaJKqQoC8qZan3sg9qx2YqlCKLQVbJbvzoEWx8oNqzh47lU8h2LLECLYS1O
i5WQ0Q1L3thK4J6Ja52ZYLHKygdlMjplJqqQiOlRS1C91ovtbfaEzeVi7u+JSrXZX2i44JTIUgmd
ULYMF2HYlTcEcLGC3z6qNO6AmpJFLtCcXWcdQDCdwlGIRpjuwGcMfMoCBPqWfSl4D73Cp0aDqS7r
vdDGYHcI4oc1rdClUB6jxk+/moqDlfw3jFiT2aie5dKEMVywNpxd6OJ+ikrP3pahtxCFnR0Vmpow
iK/j9B3W6aJIAcXazfXEBXS5DSDKHDxqWPm1Ny/0tGDlrBFj1J3xZqRQFkj1NLCiajHV9PGLYGOd
0JcXvIHGpSoFu4Ycc3Yb6FoeQahvWLVfpTSo4HqfBfFUniZXjlXv4tBFpkLRu/5/1+imR+GY5eRn
4RF0DKlex5PvvdMPhPQLzzh534tg5t7PT6TSwgpm2JKDpTJKeDX41z7D+DohZik4OIeZuW9yB2d2
k5bnaqZzcKxQwPlLLaCk1yJZGRdZTYJ9zQCZrl0QSIJX4qPgzDqgck2fdu0tpJc3nWiy51ktAejr
DOQHJkb2qGrTmfq2tH28a+8+1++5HCL72NAR28fugjaj7w1thmVGqCm9pky8PgooPtJjgXCMLL8d
4lbcOVkxpyeHOn1kBnjTjJMaVo8EvTDIUZCCedRuEvLX2hEqGjPyV6g/Y8lu+gSz0ft31Ya+CBFj
xUPp0ThVP6HsStN2HiUm1tkZghHAWZEEpquielhA7szqEzusChyOM7B5Mt3GNopG7R0vR4cFMjd+
UAcq+f7qAyupEzYbDXn70WyyOjxbuUdgbEwjjhGyWaJAkDX/iJCiwrHEYK17G6WWC8hdLLcOufE5
HaUThmYouDy6C1aZ4mcTrqMOc4qDs3UNWP/52GDEI/x2R+/Slz/TDpRuYtMkm3FervEQNL94TPxZ
guew94JPH9zKUmwE2JgVoWWCVGWf5ykD1BxSTc7PKdI5gQMCQs6lVc/P6/bLb3sim46IzFKCJsH7
qzJAKq9IL3c/YIBpWhSvGMjNivdl7EnD/1Xk0qUA6JYkwUve8VXj5+TRNnu1jAL26iSCdquXnkJo
ngrZdactPFZjnLVY7A/k24zoP8lmnJf0Y5KX1OxmGxRL1MKjjrg3nOZYMUthS0hoT7UP9lFqqaWq
8g86DJYAqR4tQnG1xULA828+o79oenE3SxlNd+fVBi1l7Kd97d5NWGYubFgGMFCRjHhvGNiK9zyL
QgzljQOqy2IoAY+h0yt1osVSlu0S+saGKpxSQXtRIdc3S96Wzk2YmzXRZxdhvcCZ1CPNVcP1+GcE
UmY50Vp7pyOsIbMLRCM71HqDU4WiRodMJ4crix4Q1jar6mgFJ6xRgNiK7xxlPliTsHGTyGe6SEmv
pRlW+Ga5q6A7JOrF7T8qE41fgtwpCoZAGAzC/myMBTjjL8I0bap6nvIOE3t70CMhxwkDMY1XFML8
q6rlrp8T1TrDGlN3R0qCFhZwiACc0lF5XEOO5x7gb/mBnXGrkCMmQQDT5BG8WL5vITo1dpUXyJZ+
6SSq1KYN+ZRsRbZv6YmDVKDoqVolxdeXtnLkNkfWkT2WoaY7OyW2PTD/JyUygP7HXIWrXtwH34Oe
Hr2rPm9e7xV/CyjokfsPUcV9rWymCTAOlzezMdABXRTiIDe5nqLy6U9yHdBh78ljbnbpSbyZ4Q2n
bF1i2aEhZ0pQEk5WuVsxcFFCRXFuqk5aMr4E0qq5Xzanrdx2PdPHOjZIP+3VR9WqRWawidXFeSal
kkVFYu65GJ4XYe8myiA2yvi9lp3ycPUOhD2RNlO0F/XDPKpB+UMKx1oS42lFiaOY2PG8/I3c8R6r
V7M0NvYWYWtSJB1bXdXqVpbK/C33TR+sm+rM1J7xN4+LIL9pmYcAEv1/oTu4DstTQoQ10M7lcGTz
2OjvKiUqk5Zaf25AiPsZHDdh2ovxYLKe+E+zxtKiq5ipWrYarfJHa/3phBlZVmFVtsO4a9xwAHQK
98wvXVeBrSq/c0A/ZMkLmnrWejgIBcwCcaD/RWSk11LTs4jce58gpD35dVRXgpCVkeJnqVr1MlkE
WrrRoG8Nd1p959H+eb+zKi9MvXy3zXxWjYkmBBE98gekbO6iAdGqErwLpJY7V1gtynVj/su/5tWc
+tPa1ET6CUXZpGfAwEEzh1suUQKV+El4q1AMesUPWCdVt8hViPQ48PjfUgvvnUJNIWSIZUgKCEtx
v3UyLTeM5H2/TEVtJ3LfVY84EST6zihPP/Xfbuu9P5zG4wkDsdkcTt7jItIiW8lRqXhJr36Yt03k
Nb4q0SU2N3M5ALPQkCw6APHvXlM0Td5RD0dJCtsfE+3yz4FzGeuNNld0Rsi8nRHaIImOWIbhcx4n
qirN157OR72OwClJthJ3MJxfWKnPO4Rq8fQKaK1hEVv1aJjvb/J2PDqpFluDTtS6vkb30KJ1pMZA
FJtNzgzgHpzaNrZPSNlU8w5V4Tnf6IXlgddr8zlCEV300DaqqgVdSvXc76uGN+OQs8fKBrNzXHWt
VV7udUxsDCQRkCkPiKFTNGHRVsofTCb18lMJrl3ozAc9q88v2Xd9po4V7F7RAmuG8hrAPC3Z3rTJ
aM+CKIUMiSSc+bzBzcMkrp4At5R7CrQTNy6J6X8FM6obTdFSNWqivocLZVfikGw3nda4mClyvg07
UChtcXW5/7aMBY55tYpfIK9OjgNrPLy2awXgaq0AHq71dINc4YmC2m+heISFmRxxWdX5yOc1FGem
K5+2PJvd16CM2Vk6oFlIVdJAHuAQn+C3KAft8+jr5b0oH9zM/Fgn18DP036lGQpsejOD7Nf5HZCV
yvOcf8IOIHyUjR2fN54qdJlCyLOWYsgL4e14z8JxBdUGYpuRzgCXsebWHcaoRB/FOYxEcCECd5ub
4ONM34ZGMA5eHxNg6Xe0R5rL0Yy66JWwYyFKp4KbomaiLRnZjEUV44rIWtND9c/LxtykGMJexdcm
edy0ykLZKKF1tzkrrDYyeILo3hJVB/RW3FQVAjJUbMTH1KpC477pl+u0GdCqYVt4MRsUIs7L/IR4
o10iiyFm+rT78yBH+xjkQWGNOAqmLZRpK2e5Hb9RKxi6PWsLkYJH2/hmlj2H9u+gNiUkFkaVESVC
37AXlExgmG6r5XrIrn6svcu+XTv43vRQBEJXUKnY/uhBO7tMmyiBerQ1drkwa0gWUBijLqFydrZO
7i3FlQnascYg1wm07OY676Jn33wJ9T11ollpSglNxY6ODwlIVt4efZSG+VZDX64ffeeVozEYRFh5
VRrTB2czWLfU3nljRBmlm9Y6zovLGq6WoV+Kf2X9UiSr2PJAGtNxQOPM3l3z0IfgcD1OUGlubpMb
jmu7TbyO4yQMvacvTzw8iXVmjMzE0b7lA1uNIuYEGTCxN/kwGg/5LXauDr7+72w3mGJfhfsZSt1T
tZpclb6Yt9lF5gkJHhr+cu9MJUmbYUI4834tQKs8aKNCJA9WFajpK53ODZY4ncu05fmfQvJvLhW5
GRCqnau0W1HnDm9SOlM03/AVSU4s7tMNndMRVZdtsjsvQgQ+9eQqUWFkF7py9UvNJhOKSeA7CHfr
2J+h+2kcoNbV3HexooKwd+7z+0SsF/IzTf0gsWTf7O8pjGtFkDUtx95NMLAqlmk9mm9Vriqxsdl8
LEm6J/70Yzh0DHTgzUAC83rZjoh4uL1Je7H0M9Be5BL/FOx9L1S5mQ9aXEzcz4vX/BbQxv+1F3PL
UG8QfcrEQiLfJjOfi9cjbcD16H7KlfNpHTQUOxcQroQwGH5V3/EH6jdoPBd3QgO6auUWq2bc+r0x
+3E8SGP1cyhetIAy7uwq5WJSXHmVL+9UtTP43gZxkKV6Uko76OuVOs7ux4kt0cueF34huWbW2KBh
0+/OiZNY1mUKKNxmCy0TN1DV6aOWkcDI2AGnX5TvPsJh8AWS55P7S9cfe1E6i/xjSjlebBtolAKF
rFEmNvV0bSL/km3vnxL5O51eaVXSKFBFx5m9cna8Jmh3iEAW3SvQ0oTvy6z1xHnAocl0KnB4A49F
x0fQlEZqtjTriO3jodclJFaBu21v7gMQ8wx0EnySdq2Q1av15M8OeZbBKnMHGrmD7KnkphHhFTLH
5QkvPs9AzREVWxCcLeo+lhuOVYVXVySlaiJHFHckXChhjOz0RH30tye1SLpWJ2S+5yjd8zRuEwJG
RDMxOSfwfKcxs6TI+jtx7mrXLAhnXWUL0A4YGVq17g1qZrL7udBkO4jFd3WX+nv70M2nLuXwihVD
C5R0bD96cXHVbZrKTLJSbBZdQYtsVI2s6QfM0sxisR+oYvIZO8MWuJfc1T9TMjr4GIZMTK71QcKm
bFAmEc7BXmKLTXzfjt/MywQ+iMhxRJ/nFubUwnmQ6d9SB8dLC7HAp6eUgijl8SIuxs1mTQ6um/sk
E63JSilF5lUVctzY4mWiZPcZjXPQciZweBR5YSm1bvgscStE4WYD9xpPfXQoVhWiyXVBLLwyZVA4
ZlDanc2hr/lpDvPJGHZ/8fFLmk/w81CJgMl7GDnaxnNWTe/TS0T7GYUlYJOAxVdZ498qJBsdEegC
wJ2q8XlQ7mpLB6estSQP7iRdqJt0JZpj+JBRxPITKlFKN5LaoPN/bsmg1vNcZJjoVw67XtZQ82dn
SlD1I16CqWOZfVKuxuYM/IlRdUQIktR300uiqPuZR1CT3AnF9pGGCYVDu3WXDQUIOPP7pKb7jX8T
X8E4nucKKvaJP6I29JhV1mhXod9uYCYm9X7kKwT2/NJgqu26BROlxuN4TeS44+UsYkd6+S5w1e91
L8pDmlIWIVRlEydZCDzOHguPPyCieCDhe9ycdUJXsAkFbXSfxVVX/QfqE1hzbaVIzpnkHVMS7OLO
lxUNKB/AuRE24o/Urfagazu0CzGFTOXRrLxDq0FK+TarHQKlsCXQK94FQAtNBs95ShN5dzazVr6W
gxS/b8f4wvO1x9n781A5wPdsv6BiuoahuEz+MfJltl3vrCT0un24ame/ZnHrb3t8sskSxh9sA/h4
RElyq3PfV4p7b//jdzyWUMtBn949Hn4Nle10Jm61M7umoVHFb5/Ii4wh4/cNx3b/Lzfln0we59HO
mwRDdJ9uCRfNZynBhjylselcJCUQo8BINm1Nd0h42TM+Eg22fbUGO777ixmiPzJyYvlgJ3eUQrn7
G+C8szEWByqwMnxvcF0/NUN5RsvGek2Iww+/oNUPj6T5jpA67caz+eMn2H7qQPJUsUtRyS7QcQHI
uYpVC3ddXe7l1VNZnT38wSxMozgoKamx2yaxUyBq9i1ESflsUkf8K3Zgfkvj7qluadE2ROKRSoU4
HcYBQjFxh0WK9A9oMcWTmMMMa4O28dYNL31EEkdZp4swX+BVjk/jS7/exuQ+1yuE/9XrAoEZL2q1
fXGxL+JXpjESjUOqM/3oif1hVpV4AsEG/mEL1Y9EpC6egqWyIQHLwDkYK8FAjXSFdMx3nCNcEEEm
9b9j1gzglB2n+4Ri0BfAhVclC4KDmv/e/dbinIEmELwbPbEmPxZkWzcl6gRUj8aXDHy3PVuFc071
mebRUi+fRltnKijG0u1xb/YJnP+BrATvXXCK0FyfbumItiPMB5pjx1aev7VPMSXkki3CvKdwf+Ke
5/fYDnLORJGiaBqMBuaBdRk7NgW6kynvfjFvyBOyxbgNVw4wAeOo7J1x57E8t4XJTt0CXIkby8vM
2rbytQDssPnSMSEhz9dSYvKbw8SKzTwNaoaYSgqX0IkkgBaOkSVDsSWbrTuy/33KNOKeqIktQdPJ
/xnTVJzBiAStPn1m8+G3Jyrx8LydQotNw3kt16un/p7tIzq1W7fw0v1/fENiIKcCPn/B1VZ2Xm+c
++R/n/RZRsuv3Da2Ro3aPzpyB1PF3zZ6kQCCpOvjxjI2uQsZc1dKshXtk9857rDKfO5Jlt1OXHxS
vMrXOFbsR4QKviRnClMdS/wyE8PFAmVBINNyP5baISBEufQhXUFR43bKy+nL43sJ+4nEuVp1fKZy
/0vIPamBCMbJSEPXuoGj9vyBZ4kq13wWbZfLpOayvGSxYS6Tsq3mCJQ5+SQzuvmncNtuOG4y6Epa
uoAKIJzF1gcN2y4sfhcxJ+IwekNP+CUr+XHxv8s+y4p0N2ec1kgGeXqmoY6nrMq3I8pXUsMESdIy
6r1poLcb6c7FTxSzxyGnHpdwfzkkNJM5eUJIqaVPiJzHaF+RKAqbF00krbluY+2o1kbqpJZhQRM9
hGWiHEKv92zGXp+75YLA5vJBYkGE9hN9a0csKZHYfLYqT0xZGLlNRhNclzq9HOZmdEGPoO5RVgiy
Ji2lagTri9m4iXBixwr3LVU2I+4nHNCa9uoJtS+MpSxIm9TuaEuwmIiUFIUdxOkikpSvE1NPbLpg
613K0h9uorIXK9a6LyHhFczlJMjdB5KsjufRbydyWxSvEI4Wp6/3P8aOblq54wGgcZ+kvkpY7Zuz
7btzhbhDn6BWQdzDHgZ2esq/IDqtRugNmFQ1UGnZxYaD4B3HLoUhBDq895fvxIlhqyKHZlKiLE7l
sjIw+J5rYld6Wzf6NC2IZMPTNgF0M01w9gtMYEEBw4tiMbflXnbWgYUO3DvkhAzfu7078hmy2+W+
MvO2EO56OB+dDyEvYtNiXtN/r+2hL42VsekdXEFWg6wG1pJxzlNVtcFiCp2in3qrtgoTBPPFDp6n
RFdmXe1C3DKRCmFIqpPwNNPgV0GsVlXWDsM2XJO4C3D1fQvyrRU+mS0M/lQlnNwf2k/SXJGzpSsf
FkLEincfj2gSymmQ6/gjw6Mo2gQnUBAXqnSthmAl8aBMGoJDn3iieA+lqj6PUQA7Cxm1oehvVsub
jaOJuUkxzmRww/N1zrbCCCmPCimG/3hMe5rD2FCUDGYEBGW+oimwFsYa0XwurZqLDG8ostyHvGsj
10ni+My68oFtCy//yzRCa4OG1mwcAvhtLZqAXUj3fKRISN94aPzJTk5GrmF7o2tl1OSzYFOwwV9e
gE9TeOtGdlAb+SSbuURnBAJRK/rJ9v3TFkYbqhb/wAHZiGoGop1pYIHN3RHd6UzPWXax52bA61r9
SaL0XOeCAjWAXwyBXRiexGCtG1gUwNK3996A0rmYzReuKlCswSJO16tZoNuHOmdnanP/9h/sacd0
jx/7UDohll0TEQHwD+STPN4etvdCqVawU7ChfFwab23WDSadW5M3+c0VF9AOg7HDnatvCEbDaJhU
YUEC/s9pYPKQKPHRyqr8eu45mPtgdU8zWE6peZY4Gea9oAiKWNXksstVpdDMf+9OvipfW9CJgjMq
ASqlexqe/yWnXbBJYmh73WEFrLjl9ARRw2wp0KBh6gHlT8zF1qdAB+o0xMEIygeCvzwgDqBtZZqZ
EzSj50xbDVp1B4KnFuQMVHIFTwqaz809f7dxw2nH8qMYmWkcRKLlMMZx/wSiTPwm4y9vssaBb7JT
4d7XN6mhecrE2Gjbx3U9Uol8vDONq0ozgntueBAEztxAU+V8JFbEO8PO4Avv6Ca6ciCgH7mJ7y1b
nlcsZdX3YdYE3GgL0tRc15nrXfWslBK5r0A8g8GqFkTo9VJrejuw7HeCqW5CDUarlIl+GUNJZRCB
NvkM5w0b3CtXjuGPLT0YFysAhE/ypm4i44pbIJNALiU7scRnOar/ojYjTXT5FxglZMTgRdZNoIVF
a/DOkuldjf4reGAOgBxY2gKVegcecbRi28JLIha+Li5mDtnAf0ivslJBEeN5GZGTTdPxOOfu8ibr
8EhZp627B1JvMCIxc9IuwKlttoK1UZSMCSfo6WWiVDXjG0JJsXcQ4BAHZ2sowK3R+V0+vG2sM4vA
rsW2lH1soS7fNUQNS2rTtNx1b0FxEFisWXRNtC4SV+s+V4iz40MIEtLFN2fxxM5+IQWvi5rEr5Lr
t41D+eVg4UFb24HlTv4a7CgLh0pHTunvjmpyIgT20JcAKw3OH2cMAY+FOx1/DUNnWYpqLiuXUUj3
P04TbCGMSkp2OW7OKd5i/KvxiJlTEmJy70Ss1Apun29AJ51cZ9axpM8OXIa0z+fAFw4TWCIfdYOD
Ik96iEGuc0BM85RLvH0k4uZC4z03Ktrkuvu2lVZxcR7QUZqLESbBf8OC2OLGbcdTIM2hxS0rUz+C
IF79HUsgXwfuaN5yLuiRNRVFAL330PkBqTQT3hlyD0N8s9vvsiJDBg379Hg/N0dwWa16mobPVQ32
x5YXA2d/dn2PWNVL4QsmsFqFdOORNAzkUkLLaaZ9edBq4PF8PgUGs58P465N7EcwMhsk83R8gfFe
VTkV0XgucilxeieIdiVyvORJGwDsUJ39XRpXYMajelAgQXMPFy95lfinjx8N0mU4Frr/qT7UMvcc
qx6S1Q7cLOV+UiesMKDGdPJ6prGs4TJx5kyd8Y4CX3iesv1MeS9z1l6qYH8zkQcUnrmXznwjLBpG
xN2ivRZWYBCojz8mg3ddiQFrSic7Hshq2SdSH5LnMguc0bMW4WcgBBbwG6F8iAZiMqFU1RwklYZq
iZr4mRbcFcHI8yv6IOD2ZyI1o7lLkAC0bNKNuXDPbDFzcp7ePSP3vTUB5YlrY8i9Ngv/XiX0/zYj
3dEUz+yR3NrMSnk2P5DgivF1JOQ7LooWDnBcJsKeJNdSxy4qqarqMz2nop14+2QnrhorSEQF9sqN
1Qh2WNL/WU7nF5GF1Dp0nPbzLu1pNehgZqf1vQhhmjoJu3hOtfpYU4IoE52inWQmRzEKAXtKDhrA
/QQQg2u6XETeQjHhKqaUWmlHW7RXCe2FzBRbRYde1pzCOeRzEwgKFxXa+lTFGF+uWfLadIl2IpHk
Aw8J2cx8n+F8uHKxtbsKnrTEpDlhHZJUdaR7ofqdjss9MnNRfsj6HtuZTILVAiCCztu4Z6xui27M
/0BtbhXtqdFx0d24CS69GTxvSE9KwJ6QdaURG/REhkag74cZSHq6Y67yz82qGGwKwWPZAfAoLWMR
iSMlpMxYrOYurTyTmVQRXzi6dOMZ+FtGH7WPt/z8X4vhz5pWkc5pbAHU9ppvz9GA0ZRRZNdUKUFe
hluVGoa0v2jNE2Bx6Qdd5fEZRI5EwmNgmkaxp5U/+ysJxJ+hCxw0okYbRuil2a6FwDcC2IWnRDK+
dv5cMo55qAUDvjvJ2X17jED6OL8qNgpBwum9VqqMeG/2ilulrI/1wXI3oh+SMQKdnaJFoZpNKpmQ
IkaDQa6TH7fiClWj32mni3xOdzZxRfYMe4+rkSa7BhGivh7AKrwlv4yx+wACM2qDEMm6bjnXbvkD
X4HMZ1WWCoWg9M0KnLV7bwhmWmVPqrILY2sKkEaIfDS4TdQoWg+Wo+ecKl2GXfekIgJPWmBS6QFP
8wG3rg5Ok8YXMbscxySkwKLaIG1hT42w+cUscJhVBRfcFEDAM3ifZwklC9pDMx0yNlngCHrwncyH
Cxtuw+dj1luKoF2hCKl7gNF4XQ5mioWzkiUd25H7xF/Ul1hKVtqjiFDBjrHgaCOMsuX5EXiCZaUB
dJowm0uu3lMZsZcCKEuKqhy/x662Hj0Rk+IdbP109aTKjhMdrPp1Rs7emGqGK4VDi2d89IqxfJlx
5oZETuZCPIv406tW2a+35e2ZSJONXNKd79vcfpYzu+7C5/x6b71fYkGLGL9/nloxd9kppYTFT6P6
3PCf6AfDyynEORB6z3tosECv/lQKgQXTklIsWGUsIsUi1xlC5tqK0ykA+84M1E0mzJuMKndqQFC7
3q9HtLdR9Y01IS1RRJyQvmaH971iKrnZPOi1Rbasw9K5LdqPb75ldRRcOKs/Y+Sq7RA+jtkGnZ8O
GQFJ71FzHnQ0RiYwMz2NgpKXov4Lc11/hkRxmTaoPvvZaRLZdjyRxPwk1FXH2yDcMqiunLXVRKZw
vyjc/H6p8VoCiD33OQJSKYfTGSyDKmWGTlL2XYH/NJNW/qzapEpKFeDFuxJH3oaFbZyEk34LG/MO
QBW3Ba+YI32Mq2f+VvANSw0KN7O7UM8/lJwRSDkNZOSuJ7Vocs0XJjmZI+a2gf+QJpsOuENxsstQ
K995yGydkLR2/4V6GLrm88eqlbhQKqZaqcK1j2t3LrMrKAMcgbMw1Gc93REE4IqXIBUzgfy7w94s
IayK+6k1JOBZPI1+6+UHiMmPk6wt365ftSyMiwqGc3XJfL1gjaU6RCLcpQgMKVcL9i/vSCmB4xhn
sQU6rvZrAD2hZJ9o8mAfmyXrXeFSB1G8qadVWwwR7S3jUWRyW3600yXKOnk2OxlwbmokucJDdFHZ
/9iFG8UED4gnzD5wmjAqGtVaH1LVOpng3wp9d2nfJBLoCvYBDRMy8ChhwM05GaUkaYRhll7k3XCV
UUOsz7llBBAq3kVjaIEzZBjMhDCu3uwgx7RLsk8bDw4cH6x9rzEeKNJmxqaTZXdX5vT7qBNsbNOS
84aF270yhlYiH5AandX4hy2sC0AhWwvNPlJCTN+vNlog9fw+iIKeUCuETRRC1DZwVgS7AtQRsGeP
g53eW1tvzrgbJIIvbnJ4L+fAFFRKQmFtkI/TLfTGObmMp5ceaWzW1YBeuHHKJMDDYP3iTy1tR6yU
smxDli7TPeP1UF8w4B5/F+aLpLctNbQdF2DbfYbzEx5zIQI7N534vTHDHi5t2SRGXInkb/yHa0b9
AMVGY3mZtv8U6ppg3WgB6wIv4bNIrPHZ8W1+z8fE0qJ+Bci7JX4ETPzvRMOKqGYRtQTbXRXDkTs+
iQgUsv8A8a9Armv2vWtXZ1veSh7gOk3Cju7lDqw/ajqqfC7FMaPR1ALcgz5tK14iHuMghuEsNEfZ
5YO2DGLZpxj84Q2aSssFZf+GyBqxpySNLDmJElPnattx4g9uHv5bFQcqdiQKlju6YL51+Nbc9d/Q
0Kns6Q129GH3VbIe4qnNZbdmaamVWRUGlRrijExJ/Q7vYJRJs9ft7B76YffqiqGFZXz4MDjz9Ks7
pT8HnofMIdt6JtkmHhmO19fuejMgBOot/8MyA3mIP5wImA/0x/uprB+N13QQU+svnsp7gqzgAcu4
dm+zxqDSuBW9g3QsxLYB6jltDHW5W6ccZtZtKD8xLt9TEHyib5O4E6bcf4B2B85BXo+APt8JQMg4
DNh3oFBUbYrqAI6K9o//4+0i6roSrGA9XbFGDNmYVVGAc96D7343H3WCD04t+bUe9agf7x6CipVt
+vmjCNh1dVPML7+vRltk15HYaCdgqFUXcIsR0fnc/R1qZu2pEhDt+yxTT9o0dUn2gb4/frpTVrNb
tb+QxZRKjo2OhndxKmI30O73cnkUErvWqST/xIfU7pdNt4iIb8U5xrKbjVzec35Rbjxar0lR4Eiy
mS6OMNSZQ78Gm5SFSw7hKd04/VJX7YIxC7/hTdXuM1UH68AaOEWQN093K+bQqI/dQX/XfSvHoOks
xyHt7mzdmCTTuTYmWJZqUvJlxb6DNs8D/VIr+sEdE1DucNdxCK1trcyXcf0khzM9fEtDHMCeYhfl
JwgRkzw8sa/tFFTrPtzJ2/8BWkwhFM2fd3uvT5fbZ1uxwR15Q5rzzNpr/cWuIKp3FqPtc3W8rsyt
8GUyRDHlF+edjehJEGEb1vAFsSRSkPb+Zk82C2INi3VGYJQTx1ypnSu5LiYjWFTQ0VFORbUFgcqY
9fElKfXfvZVrMjdIVnwiN3rzFozuN2Bp3+EEzlXbSnmWHwTch9qEebKEYqNqmLpAB98wU439bncX
YhIjVH8VkMgFrX72S3kp5N6Xf4wBxkCy8SI+Cwl/pyvbPuT0T/zGLa1IbpN+UYjGozjj/n0yRHqU
+valjpm30MADV0KXYSviBP0GOivzAI+xeuaOGfOoyC4eQl7C7sQcvhjhXtxkLPKALqOzBV5g8WbC
hQnoQot/sE1VtJbNYRyGjVKnQ7wGWlIHjR5U0+QgNPOV57Yhn6ym01kswY5FDhL53Wl1nbteV4Nx
ggF+xnL8u42P8u9c1Uo6IxL17rd3SITkwv/xQ0fOOqb9KAgsnklJwf4yScvwMS6HCoXh+pHY40f3
wW2ceRAWD9EJ81haNkql9pP8Vn8QpSlIdNY4tV6VYIBwUy7Nww/7pZCQP9cdK0qJIRhmroo0WPMl
RV8xL+IRcvnY3PltkXs9g1Fj6jbw77SGyHHOoKFJXFjn6KkT6/Ov4ZU8lYVICFLyVj1DoUlJcfH+
HW6m2a/fp/DsmMO5Us1vmK4x97fPfjsdb15Ir2ZJYR2CbrStxjUahMrU96lBs6alyzFDRu4ju2dX
nefE575AzpGZxkai9FouFAI8mjgINH27l4wcBb4HuzkdixR9cblLniCQcN4sJFxNXSRSStYTaAPY
SKMfViV704hwkounPan2Ix5Aup1xZsTJbXNuoVXuManfb/mWTEQ3VfWEhh4wVtve6JzB1TxUeKba
LBmyLpiS9Qo/E2Zq9sGNQzAlaJIGSvtsJqi/d6J0p8pzGMGhYFIMDZl8HHGbDSjO6rRTC+s65Ijw
VmUvX1+n4K/5w29eEdeABmIileSzHjHL0Xe+V8FCuftpkVyb3V1AC/YpnGaTT8jF1S0yF9QyzTA8
FwiQaN1H93+9Lhc3uBteR1ZG5koGFU+FYe+Wa/zE4JSn3IGxnOs0oaa8PIIMM6BzPvbeQVPeh8w0
M0ZKNvq91+jodJQkQyp5Kw7rs+D48HANM0KhdnR/Q8lNlsiYWcmRbpSLttZQ1Y1wYdxrotwa5hOA
XxAH1LQyKG7JBXKLVrb6bgL/hL0rSs8DYWx6dVNRa40myAbzZZXZQ9FEN6ABN9pckb77Y3LUFCkR
mTcFtU307mesDYnX22vKu2Azhj91htyfy3Kk9yz3hLbqB1V++RlVZmXlNaENenxB4n/0hD3NwFJT
5lxVNfTLgP1PVsDtynU+PaSA15ATcM8v8Tz9XhKMXKXX/qGi9fkzGs/5WrtkgVeN75FvaJYHVO/W
Bb33lbshjgKAgsheWq06RhWpTy2jlsXRpVaknOSNKc1UkGCAjpwmS4NAsD6HpdlAGeRKxGDOMbmL
QKgXBjh1+xZC633q6S1rpgv2Vp+0v0piayCdYVKtejz8FIYkd/ucQqB7k8DdYpIN51HGGJdGcd5n
La6YW/fLcL0MGA43uqcuEIPqfWJ4uEnS4sbeCRdlu4Q4CGo3YYR0YABAkAuYkdyYKgAOIEAF1Pqp
velK7TiiNpWad+SjNCKpMp43Vzg1vXmmJTwfsOLkx8vtcxOcwo30yhS3O4MIB8+xD0ABgIgGigZv
JXI0t6fe2JFsknHbXHgy/BhqSYFibWbgBsdpclIVmxwzGplSHu30xYDhRa+a5k6+UJtb9HyLxD1v
odtw9lnEOZexS7uXej7gt2cEi+TCfRuDcXbmWZY2vq9ACfB6Kb5RSWjNB+66zAWKNM+B8/4hv3ln
hIbG+RUMxuH4RWJXZWGShYl6kcKMPEKQGayVmGP77MYIG7ObjyatNmH2nZHPZu5cyjpmIwem3BrK
4fXKy4fxmSAg3fqNDOW33GaPaLltus/KmjyMw7bnOQDqILshws5eUtoY8nibchZsggy6A/OokKgu
dt4E23xWTEQAoHA0YY2ZXkxJDNGlBB9m6t71+FqGquqQ2GzAscQ4K1GCnMMdXbpp/4Q4n293NG/b
IcUtMdvIf3nbL5dbgoIEDcOrb+IfVCh1uADuGeAAE/Hi8U6AC0O7zqARFFtYQ2MgwqAAropR7Cm3
r8qo/clP1iBiwsWE7AT+FJszO6qXEKM4E4BFk4ZkRMsxNkZIsrfqVukQ1X2L02S8WnimmI9C/Wj2
dF0TA3qFiR8WnMQdldqNonbIBpNpBjcMKmIlzTrbzmWoEXrAPO4Ta1eq18Cku3AoHyrD5IKrEdCJ
LhlQCB65ROhD58+0wl0Oi6C26nkM7QkBhCUw2k4c4iUEu3eROMEPfLqxtjpe764sR6W/154y4LE2
iQ8wgm+7w/ElzkiboA/uIMS5iOdrQWRlfdjh+cojF+IaIDbWuP78EETQEXWPDQQ+9zlmhr0hzg4N
ENBCfMmwrXWuyADE6JAL6penRumqKchsZBQZSnunP8zxn4kBse5KEk7Fz2OSS7i958jK3nBu1oJJ
Pu6g8iT9PQtzTHa3R4hgJwArf1k3iIQKoYn3gWjnMyFzPGKjUWs2HN6P6d2wtT3iLxcO51HdBr/S
GPoOFquZaIp6nHz+9IdwdYNBbQhAIkJDiTi2vwAlkTxdo5Rn8EE+GpLJrUnFuqrrE5XylOML82Vi
2KUGoPdM6BUOPMX+A8jesyDI7yZWP5jt7HTJd1xgM5v4EoocNyGybfzBVCd+UbRZ91BEjnP2SKfK
ZYuxpZ+8J7zNs0nmmCHV31KdL8CSVxNzXlknzL/vIbnuch1HEeg+xQXS0MrE0y8/cCttRsX4mP2x
HUoL01Izi3twZqVKH0XeZZ4FTKRhhKYT/kAEk0OUrIUgSCI0aSYmEmbjf1S0fV9Sx+NVatBiXvWC
jPa+c7JTuu28fHqoaumDJ/mxV71CHxOjN/eQu/vgYs3jb0Z1ikV1n1hxhgk5vf52OnMqpiXZvYwU
xJNRhhXwdTQRy5wcqm5t5Vl6nf6+gvPtyXTNurx9SS6iuYlb65RJNStynRVEiPwj+b3TL3kZ5M0g
b3c3emFkLJOabCvOIdpSLlSTJnqdHnkLwagyuXtBUJe339aumPBnsStemk/orL2xCnqN7NpN1XlC
FbrdWHvHQ41j3xlh4d/Jy3ue+qDDsBQj2iy1RjkrL/MOtvt0JwobpsEjGT6zs3ypmwDvJCX++3Ey
17oclP2w4gxcz4hEeBP2IHEJKbBQbXRYa+x3Xnf9XFsbcPylyKLof6GUBxRH0o0nPri+mBYfZQlO
ndqnurAGToOGucVzeDgCtjF/mROMKVd4w31pM5+yrsCEcJTYFcLm/hxrFJO4BUkPX/W+uBykNsDR
kpJgdrUMN1A8yaQcmKk+17oQcARWmTDOm/EfGz+nDVrnSnYf5uPE8bhR+9v9sAsDVWBNWDMRB9MB
uaQ62qW8jkIv1ItkBmT9nQdQDNM1X4OrJh6L91QvYwaPUnmYsvl00eqAmk0iw9VdoanOxsq5BlhF
Cp0x2U5ZSy2E2pQfGMMNPRyp5tXmf+ppU46gAhgLG3GW1eMBdudJ5Oq84/TU+Y1m3oYQrH6BZf94
ne3ufAKUhHc0r0cJN5MHPMk7nTo0rtoUTN5AtbKSsVXYYAKYPlA3Ok32w2LANPtvUl/klfp3I2rp
zsV+MXt4PZ5nPVixWvtyq3W5rCJ+Xe5iMd3wsD29B86hqgGlu2El5p2s1kirZwyozNXeKoT5PiPX
GYIhulb4/9SkQ5k1OhsFnf/7oPYD5woYuFr74Uh74/FVSuX7f9Uv3TfTZ95nRgGyOgYHoG+IdlEb
u/U67eRD+0n3t2g1V1/l0CRCB+SMWvCGGci3/0CWUzF2jcU6HWpa4heRgy51cKNass4By7Cz8MBY
qreGmFcn33Z+Cw+tfeMVyH8UMAmJueulEml77tO26Ip3w2ZEUT2MaUkYPWBJm7StHpB0BlarxUDE
+hOus7WO4SD86VuN8vIXG1pPPONJDhrqMcUQE8p498kVTtuzOuEDGGCGx5jhA4AAHDwpfexc4cFm
Hita2VUCWDYg5TqpNw/e4HNihZqoOGIsnLFWjjHz7U/Jno0NeZ/AWbwtJMvV5JkCZ24x42sT8dZl
o1eDkzJtkNo3qgwSss34hIz0n7JrWfUlY/T3W7j1hTh3lNDPq6GVW88OMZfFAqjCkF5azIahl4Xv
cj+2cBVVb7cJJedGaITZC98ww8p6l9fDpwl+HuKopjJBxsrvaMMBhywzQ0kL5tlv7r/Hnh9PiV9O
+WH2Ny9NecFQC0toUU1Ur4o/duZzZyA53WEyG3gzgHmwhV0m1HiVMr9Q9DNmsKB3KMrcWkXuOn0e
B5odpJKzEk+cjE41iJOBNvpvsu/cLSDYMdUovjEnhexDw6HHGubGqjjuzWMpUIbHrtDuUF5srq9X
1li9aSIEW7QebBHpHmxivSyaxGFHnPPwgghnRfmRhrNexZLS6OqVu2UXjDBiUiZsjSRLeTpTVhVf
+Gdoo66lZYxWKm+sqCLBfA8X0Ii4LQqZyqOpNPISvXPfDaY+bDowmhM3gkKfzkZtDgYAtr0EvHRm
apUT1to1O6FwKlk41BzlQM82bFOGOsojICyta0yH6UaMkUR5t0gZ2PrvaTg3TDOSmWfdQWwUmhOa
ZoYyCHXifHPBzHQDhIAE8iU5Dw8h8teGJuEPUNjbuCX1cqOrQ7+JvUMc3pCOeYnVIFDMzuMgUbaT
KNeNuE1Zucppm73hVyYFojeQHvDsFGYGpwVUTx0ZsA5OGOAXQxf9Binglwl+rHOf2zvrD0nnJl7E
gjUv7+eONAlNsSQQ9bHUlKioEUzOk1+LmpmsiVaHvMLRkGpYT3wgUUXwO1zN4i7SVh6Jd1fJwL2A
S3l8f3uuLLexaPFAHbIQ3TTk91RgAs1RyaEuHUrpTalVHEpTgcHYw5FxP/Rsp4hIXRqwNNS3SSFA
agPiCXaUL1nR34nRql09wGJpeeFu6IdAusVUNdEmWyZCaOaZ+MU+hK8Zf8taS48ctb1fr1vg6hEG
N75nOW0oH3I7XMrod+FQCUk+FlLHZwe2vFSTznqK9UE9zioKyy7+71xIP36Ckfa6e/tdc0UCPuX7
+8QjZ15RRVyWUZHFG2WRbyER/h2Pb4wmoAyY5W7tIbd5ATzdJdEvvTBox5uFlYl1n3/ag+emqo6y
StIuh3XBm5E1RYNEyr29eKvmA1QJa1SNRj+qaUJ2zSGuJ4Y+evkGyfK6szyAXjFHk9AV8AiBgf4G
p4QGv29H3C0hR0XksYCNiqzIOpZL4/hOknZLJrl3cOPBEuaxXIKThf5FPOZRc5tWwu38wOsdEvWL
NM6h0RQOW+/uJ3Mi7U74EGShQCxdf6nxqUFJ50h+JQ0cs/uH5wQvXSG1tdtDVaRx6mgOrOYbEoLG
B8oifOW1i6pUmlGWGTt+Owa5iHSpRCC6wt1YxSksoqdtH3EDgHrA03J3ZoZkREZbwKNB40oHGPIK
2yyojT3LF1vbwCOcxzAj+RNIOT51Bfoz1U1CdL+XCArDtHReSH5zn3lG7Hy6niE221oY+0zgiqzv
2OlTnbjBj3JATq4uhfMpnN0baDYgbv9Tp/IVwSH1ryfTa1fGggxT0wkg+E59gcQg473uDNOGEU4i
BRoMq8Ou82otJoWNAE7ahf0jLpfEZqnBhR3qZ+EUCw6cV2DedY/j4aZnabHUMo1sIBFWUHnGbURI
4OijCFBH6TWNf69nDrUXBXpWRwem8Zn3PUgd/DXlk/M2AltLBT0VAArbFkQtOrsUffq6Y5VtxidH
ckr4pX/xQdoGkOXY2Y/tnDnRsIT5agFwmMHmwRA2yn6o8au67XLRphKHnmCHI8keLR9DTVwCzT8R
z1DNrTRhca9kLBDe0spmONgxeERaiZG3SpRWH9YIb4wDuvyyVHaKxbeeBWYmNW5LK471bpdbRazW
BEMieG0wFcGQUW0w3ASTxlLYWo9r9lXhhrZ7NVzCMo6MiJzNFDZaZMNLmS5eQggPYfmcUroTa6cL
SXsCcXRYkCGLlmnDs0jUv2fMaGtv8/eKolXZQ5PwgqPiQLh7tAESWk3w5Su6BKYWdhX9ti4bKgag
+D8hWd1UAZ7gb7hPG+/iRM+/RFSBTW3H0LjSiFq2/bkL/xfN64xXqCf4AsIkPMTL+j9EEdaLpvrY
BHBcrgCbjxdQN/8KWQVFZCin7FuZQWWB5dE2rW61+Usv9gwdo35xXstkOp88dOvQReNlYqhJdsPh
ZsOBE53JOOTjApuUTnzIf2+xvPWYiqJnru5Of3zh7cdEHUq8Z7788hI3+8RlCZsj/kWvwx9rhv3u
YDY46lpCdLRUq+XoJwJdUzN2pNgjD87n6smEKKUquHrMFYGy2+qjObiJid8q+LH1YaSlHJ7cDIEc
5O6YSWrUq7r/nm+Hj+Y3ugjp3GjR4DlAKdCsBew2ZsFNirtqVofAUYO9I4F751Ag+5wrd+K4UU4O
ubs3s2EVWdLrNTwdO0VaKrU571LV60mMi9zSl9Db5r/WKQsY+/5DiValQAy7eSdia0Rcznj0G5Qf
WC3KM7H3Q/UtqHkhTv4/2jdJTdq0XnVLyzf0WPlzhYDfDKOTQEmblp5xrH7Wt6gJEVBiCalU9rHR
c25xkhXZC5BsopVCmmKI0BbALWuxvBz8z/7z2uIrV2DaFU+VgLikmIOjrSy+zx2flzNcr5vVnvmK
aEEa0qzFC+XkWFVPKjHUo3KumE4bnZSZd4e26XpC1G8LBMaiA5CaCJrkLHnCj+ZHZgBRhY7YOhAF
+e//UD/V80aoyeWzvtVtnKIYP21l/kURe2KyoVwD9mZqmXNa7Ev0+ApXhPM8OhNezjtKQZN+SDK9
LQdjKLFzPL+3EUR336cSQc6n3W4Z4zBYUnkHVN4XMzTq4JQlnMudLHdkk+VyCDiJPZ9hu2QABYNQ
Ex5CBPtfJk/sE4Afgx13B6vXaPgcit2LP3SELRRUG2f5ETo//hTbwpSVyLiQar/uob+cQZ6A/SKj
hNsPXJEjpa8aMbPxqTdHF8i60TXn2QFs5oV6hnq1uVXxMJ7Cti+6IP/O7bG/ZsDj58+0uI0AmJgK
k+Ri1HVlPLgFtN9C+4ZVFEM5bWjOkuLjUUkOxgjOakO+4rBOSsYIkSluifHqv+jrKV2so+abE7ql
PRjd5eMQmYv/i9Ycq2ITvbxDv+4H81o3Hgt0NdJ2JuU/7Fd0M9WgJjtBmaHi4sdSlEc2DiJ23oJ1
5TI6CZS3Bb4db5rGjIizPO5VyJWHchrXrU8Yn9E1K3AfQGG4fzNpCVFZYY/MEdfvnM7uupKz3U32
OBmeTvs8aIF0hJbYKAVs0V44kuAgGaYBzaoAXrkwDKOQTtWPDb7i88xJc/dWlm2OWHUnQn0firSX
oUOkCXLjwtX+1kAaA553tS2HCGOkcoe/yGIizGy30oDdK6WUUFvKlM/euzm6LeL+AAVxL8XWjBnu
jlw0AsfWowyXrzf/8G0ESdCSpz18S7B93Rygi/6HoLWS0jKgSG/gSFbrar1WfjKcKwtfbA7ZctKk
yhSo5iHxu7bW+padSLYMR70X/V3YcYFp03+asjMpOMw2iluAziFIwMEt/ekDAASZkLODlGo1YfdD
7JDTNoQenr/C7PihA+VdXjsZtOmitnfte/H4daRtAN02hEmAwPnY+xEACyvCz70M7IPPafj5mR8e
XbtByqutC9rTa/vO1h/MCk4DPz5mPtWnxS/y4GpZdRGINetUdaQF7SrJ+g6Dor1yOZmHzLNvpgmp
Uuow1bViX81kgAZvdar/IkPq62WWTv8ilqCoDHQ20fTNfV2I1T895zJillPl4bUBTLaOnQsOIrTb
r9fUpCCqolJxQmr6/F4ESZfmVGvwkR/0AFSqSibPMedbRCRphRclji5f3EqyleR44If7J4nSHMFp
2OWy2ui1HSObiatpUGdheQnCoPIjx2tyr68OkMU9PBhdzcIyVoymUqe5VBHF2/OeQuOOs+X+irZA
e8TVdlCT2zKKksRC2KHi5GnkZOhu91WNLkZGLbYRkw7AW8rDadiPjvkPHUdbXYnSYQ9PHHJ2jMys
eqDqCCgEMO/NMEU1uRqZ7sPQxnqCC6VBXCSpW+PgshU8TZyVTzhk24Vr20+9jgGTxN8RdGgHmsYN
D3b1db4KEVfWMbG9X0fA6GFwMYOfwSrIb02y4bweutOMJHhej6d3poiwUW4uHrELr0K8q8mniHrx
IRiZk6Jwf/UTLBJME0Pki+HBtI3+CXAGdI2jkEbIlhnfsBK0n46Pmbkrem4cv00f+YD+dTVKW0sr
EC2nC8QDCK3pLksEOnMeOn+k9xJtBr6aWBKiBI/fT23xU6TapFbNKdmp9J/x9Q8BiOh5jLgpfneu
c01uInf83pWOksEuBrACJhHVnvEMibxCsysj8MCKwFEzK24Jrj/xuTrwOnTkaWnu2o9mOL1SsnAU
+TVj0eS78TwiQnEIhJv+YEwagZcHeqEkYTJfk9m5wbyQ701qqDRorypHFIwLxUSSmgfXcUGZsCVj
ED2NJjf+9SXsDOh2Sij6+6l507dRlPwHtj8S2o6X3/Ww0PwMJm+pXGmCm+8+489sNVJeu+mVhgmB
xHt3ogX1Xt0xgjQom/6aMD4uUaVCWCrp3EEyAdoXVoumjnYZKN3NakNaJ+j+ASZAcxOuLpmsX4X9
+4fWBioSPdXi5/a20tR7ykH8XWN9Ipl0/bJFu5CUMvKAyFhSTfscr47pX2f7s/rXDcqj+mVP4/xv
lNnGqZy6aBw6Y4f3BteC/pMEsP6bgbXGXjcr/uiD0Xzv3lifn1R/hDiU+F04hVDjnv7yHP9j4L37
gwAK6KHldeJchzts4x8ixHH/h+Q5sX4DcfhMhivItINPWsVRch0g/VPon4lr3nTOgizv+u+Me0L8
izS1pUHz4jgaxGislRECQb0JQ8ZzlUZKbnwXd7fcz+v7V2evC2V+GwZ/VX3JtTf5gOkDOMzdTIKo
vjmQKtJZQuXBxCBgiq8fIjyLZLI3F6nU0FchEiHIM7hiB9ORYUE7dO2vCvVyjfC5Z0II+sdnyNQz
S2kbRTdFqEl38tNRabQp0w3lN0Y3e1syC5HiNtPutl6v8lQEFAlKGHASNgYBsW7BUZEPXMAjdHaQ
cNhTQcMbbYJ7LwkEoPUw7UI8BYykUOVhLeFCCKGW+K/EIbX4WLm+SOWvA8729jKzO01nlT+7upwE
nlERSaS/2yqMxmicyIvFhofC/FSsn7b9Fy4X5jNNsiK6GC27nnARne4p8rEvHx3/hUnEK4YZ21Qi
bZXm7cupVjajIV8X2Lo3g8Xbp0L2sjs7vehof0fhcGztgJ/0SkCj2Xdybg+Mf07iCMtqzEZ3LImm
K4fsYWvZJRfR7h4qhKvOGG8wjK8Wz5aY75NSL3w4ZzxqqSP7FKAnsdCXJ8VU1puAdyE7A84YhV19
i1HOdWghxJ7rc9i90yoAX6W54ddigWQfeFfTsmUYuY+DC+QQeyUnPBsCWJZa1qtnHH4iy95e1ZCn
IKl7jPJj8fYYG4B5AAV2rhs8+zSrws7EilNv1KboThEIQTEwDBciCArAA+mghilMmST0YpzbMvnC
JPN6robyeF6aqBrJRzh3+LcfmxqR7Ex6+0r3wbZ64kCz4QOrGTeRTpzq8piuREdiPut5WOLLhDZD
yPzHoAO9o7tvMF53sQ0X8n6x4jmo76BynO18F4PeCkl6BBZrSzda1tM6/rSSz3QVyY35udzwAw6g
hKERza8Uf6Q7FYhiAfkWiwRLaxgBXvlU4nzbbuRspcz5w18T4kiXbwnrUoPZcbBomYeoq9t6pmRO
7YNFaI17coH1hSfexJye/uWUL4kL2fBVbjkwRKo7yR1LakyJ29GGdhamhTjXO5/cCii9q2ssb04o
HNHsupBJH2MZYmtfNFxtrPEUwxx57awzdh6wZl95xP/orqpCfsssFwHZeZ0CStt8XZOdFB42g4iq
pv1VavlBRNxuQgOIWe3Uk3T5dC6Kan6prpWUX6HwgDU+zGgdc2ZqMw+bVeIrp4LIzLAkLSZm2aq0
yF3nJ3ouXsqb0AaHh7s7ZB/EbhQhpedwOVaMCD5+bWGCulYNHM+VR3WnPom8hkdnVjK83NN5sxnU
UN+5X0Rqx0vNG8F4EWtb33SGKutawUlttxRXJYfN4TK1W/IA4bWuoP48PwumSgUGCZTHTItMd5Yh
TkPBP7OensPnjJQlXVV38Ehs1RDU6DP/n1ZNxz5YjiXkInSqhzUHkNnp3fRwFZ9txcVDKsy9JoC0
aPv0G1YSxJJNEGKh9LixKJYX6eO0eSMVTyfb4sQMX2Ul8VdLelsl8IMUGssyDYHtdqtB5M8ou80J
PxRto7tNzS1NfW1xNkyeN04Xh57SJtKNCLKhVh+mNumozSxZBA7auzid63yK7dPsUpMePymV0sgs
thkz1AoaYv3543vxLZVYjd8f6a5qiFDdZXLDjFnfOTEc8XtH6e9ng9fW5V7RpfqhZZRqQyCr+wXH
uuPUa1PX0NYaA8i960N3DZivR7Kc/PpY8N2qn3ssahzINUJ7tJhQpgYirRYAYM9TjpdFacVslPPn
ySJiSQTjPUmrfZISXSAapJmDcHJe4dHfYAm63THorpMdLZAjDYVKkrxzXZar1w68JDM82OVxvIPP
20QgZaG0Yto67hsHIP7yEthb6LIuS6TFtTLvnqxmGKS359qufBE9+fpCPK97D9tcZBfwvcM47C1K
65R5QvWgsdoLMGXrgBfaX8p4fjnGg+BBp+qEXZJFmqolvyKPOMIlLzbNe6+T7oqaWlJ5lade8mgV
GsMzYmP83C8qKywU8Fojv+z/2fIWLVMrwoLHuMCyq8Rhfiy8SqVPb3uS8xetF3L/vixpzoJYVLZn
Hl3+D9aU3PocHXYKu1E9xKUWOX/QfPa6ViIzleNANWKrHH4Z0rkalYLcLV3zO5SLDSM88DaxoTpC
bpLGBZNGFWDJbFaZM/wYL3+P6IPdDi/T22rPZLt6lyKqoIVfKkaC58lyMzoj+NA2VIlePUx+/XC1
R4QUiOGW6eS3/i6dE7ReBR2T1VBMW2upMu8wbsFT2zSiUUuT4/cDhs7tn/nZsyVHIRJ50o67JmuG
a2mvfh/L+NF2e9LLlWJ6TH7UD33RrXzW37FtuBiXlF7nPIoU0Iy7da8st16lfRtfTSSvnwFnDHz9
tY2Dc2iYqYqSznmKxdgY0yUJLSDpd8OXJep9QhBhHjdCehQxr2UJtBdYIG9ybg7LpeYNUVygLJsJ
Rb9StxROg1pgzvLzwFHNDp0YR1qZaf7Qp/WISHjiAzUbUJCMGhi7nx/HMSWyvRjHDs0nBEnBg4Fx
tqzFGVrvJO4KFeA43o7yH8wGHaX2kpDR/5osk6jMTNKZoxahVnETCJQLX7EYyyCgIJfuevfiWYPW
EjFrUbyrsQjuT7HdACc9dx46OWzKNe54j4x5qGjxn3pcsnlv73XG/S40XUCPv1PEzpvYBabTNjIm
V5j+6Jn/HHWYJwj6OdAUPG4iW7Yf33Sa1MXqepIkPlUGzxmJqE4ntNPlIkOt1bJlyzogIgAUQdZt
9Y72W/kMo5dx7k2+y5OWMKlmLXFMeQRiaIEr8eE9fS3aPijMCZe8B1ZaN78dgJDCbVJ2VvI3/sS/
TkCC9NeLnHeH+YzczoE50JOLhfpDzOyiBSDZQpGbCAUjq4H+RdGdE1y1X5XASA5fatS7MSb5WJHB
7gSjrvCifZP6Hf9jWHFBMatHeMSHKGZ/jg3LMTHACzGUEfZXns2OlgHTew7ZavlvEpo7gAahyorz
siPNyOBAlMcRLD0dbB8kwUod9RnRjJJci1Jqf+B7DoyxYo8cIE9AhHVnmcaSUYbxujAlCtuRimwh
/4MaMPCWT5TBVsAIiyMTk1bkNYJYfeGPlMNqY01G4PyCtbT5xI49lgh+LhWJvfNZZElVKAh0aMCL
LBWX85lAky502LD5nUcpUEnRaGEyJX+l5aNOgVqhu8DXJGs9eA5W5O2DMgLoU0lYFRRDddwBRh2o
NqG2qUxdcXyN+S8wW6D23+LIwXKTjiUwUCy3JclpuOSab9alix9SpFuK3uZANBLw9No7xFGCTWkx
dLELqR8X35Wqb3dyt3S+E/JduXczIIsOld2ZtuQwU6z+m9KX2e0sXxTuiexlJiqpCrCCG+27sVRs
eHF72e/vRmqdQPIzPuyk2PCVasc7eAtlK1c9NOwLxsho9CW1JUopwIHErCuc0RGCkgty/6TbT4dr
F7kTbMX/EqC8jMd7FCwn46dCuuArau/Yi39v6Bwl8KrQlHbU9p12rPOLHSccU+lL5n4+B8LvOPiB
m9Lmz9YOfvSn5NLhrOCBSHLU+nJFHU+31/CRxl9CneDP9A55Oq+kB+gnME3ILU2VP7h0tMPfQUiB
SOQ3wbNBx8wbf+SXLOJiFDlbrIGPS/EPEwURXznRhjA4K/1Bb8Q6R6QzaKjAj/UAwf/5bhOiE2X1
yPnKsJoT2tDoiLym3f/v0VUG1oXKEkSDNpPwCCpkvxL+dQq0ahIaK/levr4pod87b9205hN35V6S
dl6P45lJI6bxYjg85vivV4UGE0/dJpmb+51NbtsgPtODJvmnDSsS9RYHjLFAUAHU8wqQc0Qb5d3q
/FE1UNaIAtLzv+cB8tMLMP8lAgCFNKLWaTyMTMnnPI98AGfU/E/jqVlcr5WCv+ySH7Pl0ymTbuwk
J1vXmn5rtAcYaUUJRtXTGzfY14OW08voTLLBrQKu0Aw6icomolHuLFiyZVUr6wFb4C3dVd7OVCuI
0XRIsC5pJ/KD11u4laN2UGAnndvfoomKxbRzctAfrjiOkFh9LEfsrKMqlskZ1C35gNQq2FCsRXXo
HIMBQ2MvMXyANYdaOh5ZYDDtW+mAR9UQzzj0CUflNxmOUOKq1S1SdXEeCG2EO6XMSmbOs8fZFgIp
nXpW6675X5kSxzcCqs49/TJCXyOZGqzNMxNLKf23bSRvaK2Ea363y2Hr0ouBG7QofEDPfngcuvux
rrRtJl9+HrQDw//DfCRmOfGDVVTQPHrv8Q742yjhKGh06+GCR+iSwSBfXNdmtKLpSMBDCOcht5d3
OvChUkeAfnp+Kre80cvz3tK569EtmAheZItd5f+dDBZOxJckWx/Wha8nVFYRNStlXF8OtArjas7x
q8j4AHHPFSwzb7duqu5fV1gIqvBBnLDB+pXbqpHJV09vpXlujvbAggzaGtKEYGwrIbHrilKh0leq
WzgXM93ZmO5E311o1mmkqCnULh/hXsIMBiUDyOudDI3jJHSKo+y8jrP9UzFQ9kRxz3L21WqX29cm
6z0eu73t6DsZWPw6ACkWN4KhvfF7j4KMkzaJxt3iyfPosurVDf4HehAKKwurgurs7rOpPvkeQiJg
d3OAMpgA3qB3ps2p33VPZftRNSc2aaB+4k0fgZyLxW+0ey0dI1iLwdT9H6BxHsQcSi0y3j7yRKDO
7lpX/NcrjMvyqzxodOOEBLSLciXLtnFooAeInzbKnplLx4dccUNHohPng4IiEQZ3B/hHerzqnttM
U2+qtnV1CgRghXvwYDAHk6sPgcCGJy8XABwmM4aqtVLGe8TQLbtCbrZZ9TFB9wC5clurZaVrMXZN
yMxc9YRw2ZTIBbXKoQLKRdpvlzBg70LB6c+Y7JPKMByIB5A4EOrY25kcfd5AKecHEHBwrxyOOR1d
qr6n0xl9PasIaQTsZUbEkkGlsDXcA5SmxkxQTfwmHN7mv451H/bGTb6X8fu26vTT13cqgskg2+4D
tS9iwryUxtrhphaamZhjFnbBc9a4TSu/bnMrWlFaBKoNVkzqMrLx9aHlfo77n3URLAlNLm+oL+5Y
qr+3b8xw4l77ys11VAw9XFmBqiSoebdsfEA50wvILX6MjsuXaUizuYkh09mlVw0SFaPosLFXZnGT
bfGScjWAlMon5EnYtdjMmZnP9t3sJfi0QIBiDpGcOdgaweA+ZXcMrBoRV+XgC+Os6gHLJHrw+1wU
eCEXqqN5iL9KSi2/DeiIRQiADmuM5Ckie4zIyW5rZMzE1KhVKodE8dCOtuunCeBDqIOHKn7gwWt/
ul5kZkZUIW7iBXjtF+RRAq6Fmv9Rx97t+3zv+dmgMrZAn6TFDeOjAkBThM9yu1kKIHM72LjvCvLr
8uG9Pxd/ONJeq77mUaZRrvFGLocVfd4LpxG3rV8M99cteqDf41ebLt0BhyEF7F+blw081JnUn52f
fiGD2jK4BQE8MZNSqQCOqqZ/PZjyitiCqjSi2vBdf+hE8/w77Hp45QnrcmD90I5tOk+gAmdq4lpH
pXFa3Z1hGW9ej/y8DJfUobioYyzi4IGYT5dWM7QM7pSaVwdEjnQG33YdgZtL766TBzHCcEkncvU8
T0LAUsIoZLee86fS7zcXcH/jWnfpVlHxQpPKBG1dGhDhyqbW2ga6QW//YMlHV5b1OhGMHoFkSxmU
cbz+qZhRx3lxVtBWaOt+Alebx/HhF7v7UsYeE0jXbML26STHp53yMLNBKbt8FLIHnuPFnuhdubNW
GXDDzK0dTtk6PJ9gq6PLe/uSNneQz1Yk/YFe+LuyXeZcwGjhX7WmdJuNVVvFiO7lfUPgKvzsjzGs
ntk2BgXBdivTUXrDZg+y8LBy1M2PjK/FRIKJc2cHVQXJwxTIU73BA79MlAybz0tI3eJNmB61tt0s
jWz2OeIXH4PbObiW2CQOF9XBGaA2VHg60USSGGu0YggVTUV6ErwppFoy5BsHhzGaL9ewbKjxFW6E
oFvh8ITOMZRBEvgMVc1fhaZPQZIPo2iqiJQyIknZgzSZ8OpE8JC6D9Jr+tUuTH7CV0Zl+CLzA8Vd
T8XMlINvUyoLfCwdRESHgM3Y3H8Odg9V1zpL+BqlLFPzShX5igNSPM37a2Rqt784hPs/Fm7VXJRo
OWjppKQ9u/yEnhiAkqj9cq2ZUIHuaPqfoT8tPhn8UPDX0WLvOe0A8f2xR8ZnCdt5Mie17wmLuMns
poDGVHseINesqu6AT3i5yKe9uvO1641h+X45dCHgpqK0m8OUC7GzLQkrh7tJl1vZvo/w5fXWlbFF
3Sroq3fCkh2DN5KZll8+XmpxcKKABPY35DvQkR5dwKv9T7ZxNA4LSv67A7f29qGgthoR5mylAXfO
B0JPcRmPA18ox9oR3UwzaT0raJtn7ZzLaCfJbiZBv2pRRL5vDEta+ik3LLg25PLcLT+Llfr3rGMI
IirlZ0pjYeefqEXhV86mntQcbVlW6IyZq6/zOdhgJJ2NuGs8md+earqYk5+OkObjq53DLMY1dKNs
xSM0/55j1AIOc/SsBAhA1Z/glstHbc1kWoZf225NQZ4SKcnKON7zwf+KxoClwnauI8Ii0SyBCmdK
wHZ+Su25lv/SNE88Q3JlsyCb2kdKprv5F+nbUM6PXYj4b/vLttcWx0h6/IGXAkRR50DXHljJTPph
7P8h+fzC8akd4OUL2XNi4p3rZRvAkLBpyLAInSLruPnTh0FXmtNfinDhif4M5mAiRaFjFKF0OHRq
YdhnMO2zSEaTNtfP6mog31TUcXoHhGYxsQqaCPa3ktusYXV1JgOtuK8SwTkBBtA5eBwhLBcP0d9y
kjmnY1aO9jtdsfNjZcaD35GxWN3wlCOslYC1xMI8SnOy/4ECOi1PGSAUJlNXfwIU97NX8BcspPbf
yQ1ZKrQc8cEqMKgrWxOaXoBocT0Re46lk+c3sNLNnODzegFDIOrJJ4JN9RqTQy+8HJZ02ocL7pET
MAyZkXe8RmMPJJV29WnTbQUgj/fMOBeNt08icCEIJCzPnUWJyNZAEdvgqxDDC3LNO03ryMUNMSn4
Cm3O34mubjlQVPzPIOct5dTpQL+cfDDiVW9+piqa8S9rM1UHbVlhisya22HzzlbtE9vHH2G4m16m
q/YiJbq47/d7oxbitHOHlylvf6LJEEFQA7qZpfH7QLAwEtoYGa7v0sS/Zc+Dwpt1FAzHumSsNkAC
7qdCPF8gOtG/sDdvEhBpT73iEQnqXql3Cu8mxhPgyHcUapPRxK5iqoWCZmBZcCWDHRqe0Uw4Zghb
+RJgPvyK01JkKDC/USEDZL0nwI5XCNNmDf9Wqd1Uco6oQt2VEiImdAQZSrgniLqh68DZZd4bwOY3
+3JCMWDJQsqGKSgi1FLhY4Y9TWNMld3oXPqxtj87VG2K/uxjI7g1WiKCW8F6ah8ei4K9uXpcZzrG
6DVdggIOAL0spD5VKUF/ImNMVWvRJfRd0etOtmyffJAHgUokjH9ZvCgzkNfq4bht/uIRAOGlQmHH
hVQuNF6ToJeU3RSuj/fnobBwDP5WOyqp7+7OZssQMw9lz/PEUTb7vQfTng/nHJ2o04Pgy1/acZKo
bVjV71+WMFBf7p5vG5ChE9ah4PFzJVQRj2tkl16keLag1g4e5ikjesDbqQycS0cDDiam1AY1mznR
uKoEQxXWcpYoZgVTw9Hph6Syxmh+rrPtjdGghUxcBYM0SUSF93gCdsDgnZti+NeWZ0U/iWhcbB8H
ojsy15CYxB3Wroyu8PWghCuAeGLzXBuhrLc+B0vDq1Wbl32AwEMKJZri7j3mH+r7akrYsLK2iAlw
pSU7MirbC+sqCqcqJLxe317sq5rSoT+CjjEKmuCKkSGffssKkk5ueIU+AEZW72LHAoKDVR4EnIoX
8lIELQ2NeUbd5/+yvfopT26e6apn9IvrvBHYSnJ9vAZHzvTFJdUcbDH59bXO1/hm3uf3AaFAHrUZ
xK5/uF3/8umC6HucdW3wAOU4zJMl+DcL5HfR3+lp+YH4PXMDgZGH8KzRM2wka+n393Y6fcDFL9Y6
2NXd4q6H/NOPNSnPuOq9m6igmg5UeQGJqTn37OzfSgFG4KlfNzEvwFSZqiXrZPB5JFq270L0Tzsy
livm7Fzye073O+QS7wH9Hz1UPMlzBojjkuSb4wRaKB2Dom3uTimWvmUNFDJPpy9vT7uRtWCMWi3a
/x3+e645FI4OhZQ1pPimt5ye+HN2ct60neXST/AhI7eoeofTOJX17JDnuQJ78vGXOP1lsl0scpwf
eJsJ3lruLCxMbNMTjS7WhFgVwPlhMgl/hxz3I/DJoJKLn4Z48aymsNDD8Hn0+1yl/yu5bE6nSdd7
3gToDfMZcu7vWQPWhgAqgC0/2DxXn5nloMqb405h92fNf454nOXT/Jc5wSDzg8Ucdn+JnG/7abId
nqEDGzsLJrMxvJd5iU4Rm1QMnzZc/gTM/jzLxsLJUZ8H6bWzkevv1NLmNh4zHtglZRjeRW4fjgj4
U4nujgQ0tmc0HTM/c4/IBApvRiLlS6I7RDpIYgQeJi0ZMpWyGWIViR/gjdE4EbTiz7HmvI9hOylo
kh8ZVS3DWSWFojDFm4BrcdGxQ2eyOV1AkLkaG/txYg056z8MlnFtbhIUPL4/Sli1yyRP8ZTYnOeb
vtZyyTpoIi4SDAZAeqOvxHQ/Fpmsg40ny+wZNsI37ZMzt87b1dHsEv0uTMAxcCijF+Q51jgXWxJo
5OI6bi6vCheYJAfUdDfKutfgfwtHm6PGFfbyh4Pomjxtp572o/8lj6QwMSn8bVs18dzmgWUJBlWA
Ee8gqC8OAyyZw0VRjQ25x1fhpK3NPwjo8nsAT6pNg6ZVOowMR1WDiIiQIdRKX1EMmCVV6UmJdBvU
rc1/pRSQkCLHPoGH4qvvZMsCQzIZLJGmYHS21vwmC64mizUSXHjmo4PU1Zf+Ub9ly1SegTQfrshE
p6jk07NDtmfMrK0OSoCyVG1uAEKrJCUacx+FChlf/VXddEpOrI6yZBrGuVCY/SvETQ24GRPWhIvB
UZelReeaRBYJ8Gz17C0daq2g4SKNBcDnhCHNPQQUSo23Zj8wvlto2KbWXiTGRTTN6XKhlCYmePVg
aOFkIUiN+1HHEOnxSKSw/5yCGY0ffr0fCASgBkPil9n4ms7Nay8IoXkYrT+0ZfN1fxW2nm3QS83c
S7CJqrW27wPIgnMDrVezYz8SBrQthbbo5dNz/VPNhzo4nrReFpSaQ0AluZohvB6gZudyd9bSMyUZ
HzcCD8lNdfd/sQQWW6VOIoWBAuPloURfCiyuH8Ik4LMxPIKFJGkhLElyqWbrSmIgF7Rbs7d/FXU7
wch7Komnw0y+OgzmNYkNykeUUliTif+PTzyK+8tgtxca4HVDKNg6A2aF7HPwg9RkjdqNjpZmNAlX
EYzQqZ71hiW1LbC1YH3xe4N4wFXXbDw/SvnCXoOSvgb51ocg39CrrWFci/mQg8Fdi6Yuwr12vE4r
lSEHe/bT3NkeKNISlZ+VebXuf1IKVTjRsdvf04hN1cbWp4tKRET8OjT8EfkqFbKEqSjVCuobS/yY
FP/127qECWZ/H+YDjQmO/C8GcHHdwYbWE8d4wM6itqZC8QrOt0CANdiAV1NLt5sRth4yfXQXIiwY
HZsaGfbVLqlFMFbwDnZg2LxFDQy0HMjwy4Vdv3kCVZaoavRwoqfHGcpFJTp4nROWpP2T8zhVEVvP
cunhD9U3okvDL9J9arpKerlfVugNMJ64yC27V/sYirafJanJYf9ZPzvW4IZ52PkNf3vcM93e+zvR
JKTu4UXLJ8qOO3oX1MwDkCaH3B8LRZHNBDDIre2K1mQSYgtLOxjWjvSybtUUBh02iiEVSQlttRqc
I8plZrZ9fnleZjrItmq0kEbGsyssxDKBsHAjBQ4Chgb+S5PLV2cbSqUk3KyOGejedEH765abWI7S
TCsvW4ns+7JJxQm96XEWX7CSONSu1/2q/G2NN8IpnorM4RHiTNmTVGC3yhZDAhuuash6w0ZlqhX5
pQ0CRLyebeL/zmcNuSjvyfcD/DLllnCgcEuodl+Da9CuBaJkFYHitRlHp+Idfq2U8zkQ38OIN25O
Vm1eHwKTzM1DONjaaLaA2zcW011155zagfQEKYNbsLMDNvBq6QT9t79FKIOAKgjGMTIvrEuZ6SXr
MYCOhb8Eqn22yNMxQYvBILHjp1zvGhraSDIMXRF2NKCirsZK37W64AHLjh56oasRKbi7iM8ptGnr
NcGI6yPbWOEjXVbLFGOTDjQmqVRGoGb4JyKztA02vloTDTC7iFWlMxN8m6WKsAikXLqJn6KAY43/
CReFmpel+z8pvp3fTaQa9scme4L0H3dwlP3oZqWYQBlkN7FetyiamjVaf1djW0hTlovEx4gIow3B
g9v8DJntAt1kLMlsh/Ng07QjTNyCx7sdGbKJSEGbjwvskzG3oZblMlXOKF+bDNp+VWhNxO0nGwOq
hetK6SQNfGWgdBChMkeQDTH9E+FMSZ03hkc0JufTzq+m2V4s3RJO13STNv3Y2MYllgddf1xwsaOH
i/fKRBiknE/I81do8TUPd46vPriqBqfhn5Z5XgTXH7HgOZSMhFd0dZOse0qX/1P50WiQDC5ScEf2
2jXT417SDirmMiN/jfC3pO69G+cSAcPN1bEYmK4zx1pn3eusQNAZG01DnVJJfKO9GkMrzHaz+kt+
G8TJzKIeLJh0uP369uisu198grNicRUK1f+10J/NGbmpSB/386yTYMiWBdQSSkR1CyQnH5qFDOeI
AwVi2gAHESCZ1azSpqnBAbqVL7iKunm01UZsbasJQujnYiqSrxzfrFbIO0+eMl/ZLEBbpd0Zj5Cc
JlhAsP2P9dcMfB00cec9gH1nyqhIHkzAlu49bpIw+xtL9GE0ovpyaDkXOpsSMs5uaZX2gr40QpTF
WP1fqUmI6AxoTJQ6DB6zytaJNvgEHp2my5bmm0SMi7P0wDM3Hml7SN4TcF0jZ3V0T1UaAZFcoB1l
Y7nJAZYskRwlkJqIHSGdR6e4rMoKlJVIVIX8Scf0IZu0RuSydhKvzjJKwh7nbqUsJyxbrngop6nQ
lD3DLKnxFSiK0SpMTtps4vqicv2tviKfn9loBjYUiV6VvNZW/5Ha1qF9VtrNi1wml2wOUDyaDuz5
ZGqa32KSpybOQI+v92D+aplnKEfWDDqk6yetTaJZHvB3kWM50DZuCKVEnw/vlsysnUwWij60t6XG
HWWbXCXfZtp2EoZFjVRl+4DDFM/xiMdlYIfopzErw5RduZ1q1l4d8yJCCTlZBRCn+5YIh3BjKX7K
9pM55UHXSjSknYyga6baXhku2b4eBCSRTfhkGl6/HWVww0WdssZoyHDss98CGFtBMSLqkQxGgVe8
K2gru3STugyekJ5+G1gbtXHRXpDCaWTwvo8a59Cb81U1GJSiTXqm2CeuYi2wd5MilVA2KSSmFlx0
04cvoeQjTrgz8NKxzgA+nezcrRI9btnOqfU78++kLa+e2k6WRrf1oDhkBhf3ZwItzfJizOqJIBcK
WYyJZ/rdNbKuchP7JkCfVjRrfWXGLLL4GYOH+Ee24jPUYuxNzbSmtEaE/uUPvkrGtFZbIG0uO4m5
QIm5Wwn6hrmndfTU3EFQKy6taEyraN9hkzDfItScQomdbB+FN9bIO5cZvBe4b6wbcvUS9kxY2ry4
jOBUIHqi4pnXsICKkUDZVPg5iaR1N1FOH8xSsNVmHlPeJsG/QuVb2EB0dQtVmWefz/MY/yzGq8KE
HtiFfYLys35y8gxaFPgxOUEKZQV8N6bHaUaEhXfkRd66XDKk+OJqqBcG+avopRjFMQJxyUOrAt3y
uftSjXukMS6FXnPYDKvbBgYgxEqNu+OVk9d3khxi50ZzfOukw5EaJR9OoJBBO9qXB/Ezo1xpVIlS
C7+Heno6YJxeRi90Q2Drn5uyGQKvsdGw7hJ5HOfmNfKXgSAN4GRM+Tijx4v/2CRr1pLR6lLOx+Im
q/tu5qQN4czOrSNbShdPm3tGQt5kwJmh9L21RXy8TSiKDEiqIrC5ECq/zIzyFjMLsB824Xz1+uzM
p9F6OeDCTi6nPm8/LVxoJ0z0Tw29dmjxTmbT2Pr8l6CuzgoGu83aAIcOuzobbFtKT3xJK38dz7co
XnvvjlBchOl69eFb4mT61J6SbvDIMzQVNzkignl5/8eJkwO6agmIWTnWvPAhRmSqNdLi37VJ/5iP
iS/XMkiQeHe/hxMJ/IuNVwv7vg6J9Ti3BF19wV6g4CxCX3CtnYlb3nrY8Go++IFChECMZIJKTdvy
BwOnTsrbDPznY4ciLRy6d0/egz/7RnmH++jjwa+Fi9iBIn5O8eZRtxVZRo2WV7rltZZfwIVEIhT5
SnPOuPaob5aNEN/aUGaJLePkoYcywNuNHJnxiSEnnX6hYMf7zx/4k48FL40bzNefc8YFtKjo+Wj7
SIZXOk2XIRqjnVfCx8qePy58FMu0tfRTbReRnYJfMcjlvX1IMP0/uTWSCbNzb1JA3xvzWDm9iwzl
tssAC/7hsR1VnTZ9sPpW81hx0BYbtiBxEhraxEbBlQ7Bk4tFti9lGbi2mUbsrWy6SUrwsnx94lWk
gyRgz8WkEIOpMWEMn6O3hJ2T3VPtjHNCpRByH1xzgaagDEx4CmRLK0eWdYq+xR6Xi65hGEhYCpzL
9M3lSnLdph+4e66foFtN/fqB2OrMfpLiJHXovuuT8bnS9uwnS4SLeEYavkdar76JGslIftEzW88m
/uCYX0Q+uoD856jQp+Ytzfe1yqYC3mbMhRky+qyiEakLUXcEkWahzgbkFfQoXgAqoJYttHLeWOCY
GdqVFFrq4rBuOUQyQFRPvyerH6sAp4fND0/9/LPYSWy4HU/bmllhLPrVbK8dGeU8XgDTgIMYos+m
uhZtWojL5qN9FA8u0QPwRHnRwtn7Nd4jKY36PgOy2mLzMs8wdDzPMZaouIGmDbV8X8ylbxDya08l
S7PbONJ4lEnZC8DKITiOsvwyRDI9y8DOvNrP8qxkAMvB3hAKtVvkrmbpSD+z2xhg7WEgVMi+EdKK
5YwOzeg73vUP1Xee+jR7Z1KiA7WvIydXG2lM4RqcOM0M3XNfPxm61wNORsb3sJqSKBNwaLgwp03n
4e8MNqv8B00ou5sz7WGMChwmO7inxb9wvj416RtnX5LCie0qmNy6sM9rrICwaOKb0X1IsBNAn83R
orEnc18i2aUU61uRwMH82xprEeUuGqlaW3pwFGZnwPRcztLODMk+U05RvV/Wd4pg6uZWD9HtT4cO
XrAuRZvAO1E49jvC5j3Stl0Tc1fHkC+k7ulfk0kmh08UTSs/ND+QxHy2OvtVCpuDC9C7qVSnwvRR
LeA0iU1FjFgLOk/04TGe15BlFz4Dh8FKkEl4ytX+efyhKAqZJ1lnT2hsRKws0nnda0oVym+SkIYe
msEb0j78IAdIMoPy/4khhtJuZMmamD1aUIiARx2T6m4SNwtAjhVnwOB5OIwstyOzBz5pseQS5MVh
8IeNLTlRiCOFar8els//zYOsQtMu9nOmdyWNFmLYJ2f3woP4bfI+td5csHqcibn4pG5IY40gw4sU
w6ezLZ9CPzMZCApnfKnqgXZH9WmT8A2RHF/fBrTis1fWeS90wB3Pj+957MJ+6ir2A47784CZVDzn
OJuzlwnb59+0GHsljyxSLlunwpo8pUbwHTUOtPD1I/HXCJ/k2Er7zvFU4qXi2XJJUs06D86/Bl1B
jQIfxiiHbszbq7Apg67Z0fEPUrOTLTXCSOInnNcHrPTbhvdvlBDuSLBzYfBYPavKY2SOBleB/G0m
r+UKTbYYFaWG+XGy5DtElzV+RABq9cs9SenM6cKwDnZYYZ8by7h7aFQ/MAoS28vhuH9eUM4rvVtR
VFGroYbzXMtgtFKQLnjD+CX/YYA/qNaZoc2mBcp4zhG2OGGFHdEdVNrbEh3nz3VrMSnlW2CR66Ma
C/vOg3dx3rDqPl/0eUK91DCXQ0T+e7QkTFWBVtyDJ/d+/o0I/Xpz/yX6xlUUEEjBf6PgugOc4Tr3
/U1n7cJ/GfyHcuV8+TsS0N048DTPoFCLz9u4H7jfFlwoDttLshQ/YP2PfI8S5CmHQp14+7kWauV9
IruJq7mtE4LhikORimOeXho7HsI3LQ1xI6H2VWradcqGeG8YDi09z6dJQTqNsqJYG7EpELx6I/oV
K5pVzIm9JWY7Xt/4JshiAjuRcD3JCadBJcUg+9GMWiUddt/qafuwvIwSwLLSNyus41AushWaX5+7
EOhr1/6uW0anLBoTss5M8an9ALhujNsgZomMpltaiqq5ufjoKU6HWcPBIqrOnOrEvfSReZcFfJ/B
pw0Si0oNbpBkpYnXjs0klKX5AVRes/mR3uQ4Xv/NrUCJTWqSrJG6ZgSb6ExSZ3o5hZKR1TWpTiS2
AWTNcCBpFAcfG96Uz4izDwXP3RilRaW0514Ks5kdv+6LBrwzZV2BPm1DnoI9gxacmsaM7bDLNY8a
BWSXv4G4ViBqYJjJfEyV24VkBeQEbK/lL5IeCS308w2FsKJBhUCJnwzJwrCYkYN7uzwOc2AvPpYk
6aLfZbGiVO3MKnJn+9dB1vSSLuRnoJ5KLgBIFjmihOa3671jsh4kDvetd0VH0MrrJjgLQG+nuCPK
mH0kAmaLYRlWl0zUUZVEakdiWhOurhcR5pFpuapDC6kyigQ8q+9PzFXEIwc5L/ml0BOtChROTyNb
oUjzBtGMQhHUtFLcbUR1EB/oZ4viyCQ9FfkOjwNEeA+I1EHoiN5a+9OV+8LWFZitpMfbRXBF1MnI
OiazhqOMRtBishTueq9aUQ3FHTM68tavbw3J+FJbtje8ApEcEYAh1bib2aXcSzWb2HWepkpPKrSj
SwmIm1U18fKPaZvH5qrsTWnIp65dvPMe17ZrhXkiV8+xhyKe3lSKud7fQr/eGao2Xgq/Eatzpkxr
qgZYvO0gorJzY/RuQRr8HY7JPKIYf+io6msBNPRCZydf6trHlLSdJsvJq+8FfGoD/6ZqBDmcok+3
3KxsO0zsE8Hqe91K52ggk/gbH/6oBxDrZyBKGjt1a9sQpTz2HaOXBvH4b9Jsu+AozP4Aj277CS94
hN27oFnBSPzRy767Rs8WgJMFO8UlcJYZJJ+5MnoeoBDtIwLDTas4RH1boav/VbEhwFdMhipnUxtA
9WuEW9jgPhW/xEy2fXmbzbx2i/wOlHSbc3mbebDw/cvo2kIlhB8xnjk5DqRhdXK1eik+RR4ZmdSL
zn7MFlugRFwjS/PaS1s8A/LecKY8y1RxNtA+zcHZGfFBmPNJ0P1d8r8VAgQBKkIghmFUrNfAISs1
Qy9LCAy+OS5zdQo7JKbfxpoN/vNmE4usT62+fpOu0D+XwDyanMRNr3MMIX5VJm/CeGttYu/qVpqS
o+wXa5JMfaQsv9FBA4jOH5PlrybagG7BUUKnxGX0t23G/6H1tg/A9ukUgnuNJgW/15bc6z9S/GKJ
LGQNqr3kt2tGk6/e9v/ic2tvgijDehm93WWY0bCeA/NF8y6eu9R+GN7+ZA4oBLucFkBB6eG63ABY
2hqBlg3WKjQ0WltDgyQdwaTuTQDC6Fn6Zgap/DNftFMxXZntzhJ8z94axxqfBbLUXVyrEdH3Qm4I
n921JLIsZPsF3FiGymQiqxr8OvYDxzgxj+g/xt3YhEXdS/x7R3PeqKIKfy4jeHy2dczHZfI4iyG4
hh6t3IOarrSVs8oM3b4VKN6Ixzw7mgTa9TTIkezRk/VxvxaMzmThyk7fv+xUTTjHRZgjgOtRr1p4
cE5YluTzjwr8ZN7VwW3lzFydUVlxHRfiYwAKpOPkcDaKXyTEDjIrVP4wdmL06hRr805gS7kMgpmf
Kk6zD1RnIlD7QA+mQgAmNN+d9f4cKsuY+EeOTwpS9PVnHRioCzQwEjt9/DbzEM6saKtfwmHKH1FG
HQZHEn8CAfa2gqWsQ7k5NQlTalQ/7Yj3pPXKJj5eUgYUuz18TpXsVb5lT8cHXaUXPncLc/p0f4eW
UHzpdvTFJCDK+MFuDx0KuB++2h8vS0W2kUKCiC1ZmP0AWEjDbSOqc4MFV8I9RetaEPfKBIhL5ptt
UU+7BVGUNA1WdsMADCkh7k/SDb4Ra5Ia56+CqOusHLDM1O7IC86Jer5vS8sAwooP9xGVwKri2cgB
6bTOkOJA89lPwruHNqRfSCaxUOo9GV+zR5ragluPNDm3x8wUjIN03C0mLZChsC7QIkJwAhF5geIF
23tdOGDdeHPszZI7WQQhUpQ3a9JjJeorrHRTeVJvc9rQ/7NXUGU8GzkwkTPZoqyNbZeKWS9uqAfc
Y/Rl8NigNzjAmX5MF0/KUfNsU0CGtlaRrwvo2Pk6gWCIreOaIZN7BQg45+ObX1Ie+p8mw6CvqIrv
ZwJgDBoBSLnCvxIXKJdobHxUn0J5dfRPTID++KgVLYUglHFksGBjtpYOLlGTWc6tihUsMm8ghaBI
Tva/JyB/bnXnYHQYHiIV0sfM1Mn7u8KsPMvX+EjmHxNiHDy57PeyXe7weRQwfsz47YhhQP8pzoBW
MhfD29N88JfbimyxyowmFPbJAZgNpOYIViEqppvxZFLUh2Z0Z8A5nWW4MJGu8yYhqmwiT7wdAKkG
L6ynN+deRNb5XXdyrAj+EVzqhv31ulYgRPD2WGNgxEdaodUuOydG+JPS3DS9vJJNeleu/ojVuQTL
ZqNyRA9E7uM9PD490tO7LrIbnrLqkkeCRBXvdh7Pxqs5LoLnTO+8zaQfkYYCyIADdLFxZp/SgtFk
eZWTnsFwFBsqPisvh26+nx9HxjBFRCPOJcZ5ch6UU4uP7V2MS7PFqyi2r3CZlFhVOJKSdKYfnSjZ
Tk+xYSqejiEh8rju6Ug5BfWS5CQULo7dNIrWH6MYLLm+/HS267Zghs5yFFb5hFlVL4seLpK1EqO0
KcekXqLeFlFLekjCCUjXGtIMjqMBmY0OvBTIn5O0EES3nxQFOAHSInDAz+5uYvnKts75YvASxagb
REDs2F8+aWChshyNwxofo81hJDOVo019RGn6NTmyypt2bSVGkiyhjZp3dcxDHwcjVnllc2uz+W5V
B33kIL4gj682jNYkjRWJ7XIH97XZiDiI+ui/EabmFGxFaEGTTcZGrtI5PvTQFXk3ZsiNOrnrCPnP
CcU1ByL9vpgR6GOwdJRrJTSgj14E4np7yLkxVp70ME4Wc17SLeYOUryUOv91NF5kumWcMHSc8zWZ
nPiObw2ognz0gGVSOZ0rWVhZUM9RRaQ+La/ZqSJA7wYpyX18jNlxdYen2PWz1kLvC066w7dzcDJY
913AbzD4llWbUw4giNUeipGJaQ6eRaw0bgxMImCPu6fLYzRNno/VP38vLHSYs6j7frlTXCjNd0aJ
6KRmMobW2Yd6TuPtqv7K/zzMHRGCFP9Ub5jG/sNSAKMhQCAtWnhLUKNGosXDag5n8xCoeYRw981u
H0tYmoixQvFCl7Ikos7szEMi1ZcdY/sKXAtK/Yh7rSuvKSRTndBRVD3m5iqyFGPUYA4zVNJB0NPT
Nq8x6Zpe9/2IrerDlMuLLnZ1YDRb+kMmhpn3WFKTI7uPiD5Aw9IihE+drO0z9yE6crar+TC6D+R4
TGVvuhVUCrcGFGHR5CRkxEJ4raZHlA3Sp36zb+jsa88vhz/ihMl9C9GKYA3zSsSnFz0dERqpoiVF
fxHorIenVxqmIO4nxaKsv629RxU1lUyDfV3Fk9HE74a01mcQ/poSWLxPHmBF4hnXVOE7tDcyupxt
oIRWo4s0+HUzbPov48qwmyYuUhqVXIosJtNB6RbFKc6ccy6iFI6TQ3ApH1oPE75iNs9qaSEmgYwe
hSgeYuJ3BMkxFXQRvy6gAC8e5AoJKORoB/pN3Lob47nNu7ZqOJloQBW7JN0EPpZuqQBO9fGgFwsm
VexbWUFy2K4O8FWeJ0efDbIsTNsPF7wys4GHzZf1iLfkqNbuRZ+nEoAUVb5z6BqW2ManO2Hm12I0
34L/EUn1NOCMUDYdRPgdt8ptOSdlznb1pF33mThkX9FF7pNEXbNHzF/QFPIXRyRyZoy5MF1SazwF
tIFTAmhbkXvvA/qZGz63zVYbsR7iW7/ntrUlEH5DVt6dA6dnexwlJ6eBrSDKsWP+v7m53o0kr87v
4aOcI0uO+3h9E8pVVty+wRpf+EVrpfGOk1tPvQYU5p/15XJUqUdEJPseO8B7x+25qU1zdbxDnXck
tF454BiDSI3jezeo0qTsPto6KWmRqTkooVjrzNAiKkbrERP+XqhIy7ky/QcZ5yA6n9mxu73zKfRn
3+gkNvKfxiXA0JRhMG16NJg+HQhSeX6AYVnI9LDyTgJh2cipvIbGy71N5VktAsEfaNYPjeRBP6kT
1zvhFNKRKRp6D7Vhlu8oM6/gGFycubuZVex/OZtyB6kXbhb5J490TWz7t/h29EVFd/59k9a1cd8N
gX1VsFirbiu9stR4xZ4OPAbe/+DXy6sNlC18W/Mxb0bBY8nN86ht388AJpp4NHvvDAv9jLeXrKmF
9LhTT/nprm1+Nw4sSgMnK/Cp64TYbp3tu9BxRPlqCfkZAefBUS2dLowWSw5noiG1izvKpz/e14TD
UDfXW/G6RBfDs5wBbzWIHIzVOTHDD3CHWQL3s4UNXBgqCySKzoob7zHVSzw49CxESKSTHGKDpJVV
fCu38juFcJolysht3vb9PxZKGFwFnm2bDDicrfA+K6P9cNcpIN1WFmyBBEGj7OUgnxIM60DrgL2/
HOD+NGaSC+FnFHqNaW+SGAXhHNJ4dhljaV/aQImCzYR3V8FL1pk9G2y6en3pyQ29AA3zznDHZ+nk
n5yXwX7swudneMARt17T1iMUufgI2d25irnyVBrxzNzmVH8xHMMvTAwPwiAFNjPZOYkDI3vhqrF1
6pS5O1V9LVFrfVSqNPY6RtEZCmHr436opyqX0Ibqm/p0d8a8x2TqlOqL059MpXWIgXxdsiYDYDw5
f7L0pqHBWC0lg4+7Dwpk8sOunJLah2GlJpWfLb9xWV2DrmNd21CaG9uQVf8E+XAW437DHk5lkNxs
y+Olf36UoBdWmj2l8xE9BAdUIAeXBy8ys2xPqJRPW5xQWEFE9rZ7PQWAYu3JnCzGeFsGV2hPO1IC
fq7Fgnt3dmFanFm7v0LCMCLziYX1Gra+Kbhn9wIdSQE29adPMpRlYdz5wQV6ktynHd5qfwT+IPl/
5qZLlnjJOVlKQx2zFgun+Ql25Rc/jkXTr3GMkjZ+pnHMBm/JjO+BiKfTwEm5p7ab2I1bxPRlaX5B
SHyjgDgtX565H60J5qPbB/IvJt6xolrbBYgHEHi1jBnLqJi+KGmKykNFR+eIZrnIXqDS7VIlXDPH
LovEIeKthSn8K3W5Jf0RG98k+u/NlmTGQc/8BRMygBNnl5mkfx3rZBUIHF7uG+lSdyEceB8B0osi
QcOiRaPyqDYwtz0IUhyVB8lhyLpzWGXsP8Hs5EYUMr8qFZ8tb0c0cZqgFPX4rvy5p9Hz7KavmVqt
eFC377/QfQpsEwA67G+aH54jpr1hBsDxDHd86+iY3Ade120z3/jU74vhJp5EUYMAPrKn10LVtZvt
7HZgE7n4N2VIujvE+8+hcHcUfbo4uYkNFmzDpDPhVScLkQy4bJ5zXQ0+cXRrgmP3olt0H+LJ2jn4
TT1FGhZrBImQR2p7UWPj1qmAyj8Lo7PrQ7sHWwnhaSXLaTjHoF5YDmmrJvn7cV+N5EelqH0zanQP
r/R1QqZYCuXWxvdyvVR6LaljcVxCbUmPNAJTuU2cV4BtbxCzE/sZXJ9DrOfh7P87B1lHebYa34XW
rij9Qu1fs/O6aL8RLBB58ZFqkoa9ydPomq84SJYBrGnUE91M6KsdTgEQ8x4JLDNjAgi7/2IC7WV3
29gFeW+27HsN5YWrvhLtZasNm9Z4Jf8wB00XhXvtwf5seB+FoEKQHNg8UXYZVJm2oKHTGJ1rPtVa
BwEZuuSY6e/nfRaPcDWXVDyeuWqM+yMgbH1dGCvFGx78Fk5k7gdhVHRwb8UqdYWHgmmMxEyA/o46
WBAt+iRvgeY1reioQGVPjqV8hv9NZIUgJwzs7dWYSOeTj494+gy6jwCg3NjAy2NYC2z1YiEVvE8A
YAT5X0bPSSig5B2JnObet0WPImFXtvueOpmoPsmkRgHH/ynTO/qaZdIIP2VotjbdBNcQ2UoeCE4V
NKNt2nF4rjVLsVNdKzpB+ruPHA0lERgNmzxxaX01GnOXv4ITvVUV2PMd6qj8tIDSAwwe3YhyWaPY
oYUKao42RRanR+JeE0V88YC7tFbXoEkaiSAZdsGMonbLzsqHGAtBkbM1Er9t3phv0uXRUgS1Oglg
/qtvp6RZv3nfUA2S5yQYf15SS+J1WSVeVHaxnhj1l3SEkeTCO9T0btI732kj+/nTOcqmy4Yg2GfK
IwQ5qn1QvI4vvqesqCjxv8slz3iij6cc/VG4SE0gn2hMoy5HacKuHsB+z6REjyDRCfazr75NJxUo
FGl9zlpxGEms4zo+qGPwiHh9rzg6q/BC0Yudloq/heHjaTn7WLjI/EVyMhH/M631CyP7+O3eJamS
u22LikOmHjyeRakixp+DGLpSnWX2E7FTFWb4qTkY3h6RMYIOIyoX9+JHpuX1FMlDySWMWHgOMtxT
CdAwF2qknDZbAPQQirRRw3Wp5bEb3y+Jpxw/HwZiONJ2CBU0ZjXoMeF4O+2n9PX5yH2plwz9RdeH
LjhsgGmnvH6XRkEgXgO7Wq/jEKzdxr1PwnAOEkfXD9Hft7DfRUlZ+qBe2MQ3+KgWfWlH+b4zjf83
blKKg4xK8iYks5lH30s6IZNd4RrsBxa8z6O/vC9hGyfXX4u+Bia8hGSs73XmbYuzoZF8qjRXaDkX
XIwtv/3t+mN3/57d7UW9Vjm0pCELlsp7ntOGZXfAjOT2s3g8sPkbe43Ximns8PeWfvYppBaEBcr/
/f99bK1vblrHWE668MtuK3yRsFPQnJ6WzVLe3SkZiNLgTWw8TfMat8+l6e9L8xft47xdUjiLjghK
BLepq/QekAgTV+k2Q+7P98MzvRXfXDkmAoS6CEI7n22EWxbkO52c2k77fDL5VtxchHNXQzF5Jx6q
VtCLhLm4oAPtr+K+2LI9SkumCg2/z2pIa772MXoQOYk3Dnv/LWUfP42lry94ps06yq8CETEdSXNA
BsILCLI5n1zWQK4TF36XQPhSnuLvCQi6k0x0354ecBjXDCu9rTjaK2JxSLaZYjMekrmxlJB/MxOD
D6cXNshGFzWyg0VdbSca5bSpzMM1cfC//tkK9RXjlW+xu9XM0EDBV5/8i0NHZstHAzgnPZCXjKsl
2NaYZPDJv0nLBKSMr83kxRFT165ePUoXNwK5/Mj46mmAqkLdiRkeGmmBSWZw6f/mHNKlmXzNnrl3
ZIzAYA8pVgupU2myuq6ujqUap27kNSgXKLY4t9Gd5TLa++o8mcm8NhrbgSP8pcqXID9ImrZ1IQPm
lz6pim04gI3+dgEaA9PPHvUGnJNJgfQsguIYIq4STEOkYGcxNNqHjVtYWkTdhKPGfhL9bZO0ohvf
MngT71RUkTIk76ByBzGq3u7Pzspjs7s7h4Dz7acROvKL4QnG9Qys2916DzJkrw3tFDkBuBtJ1xZc
KPKuiYT6wSSqhxsgtJoDZfQymyu5CtDkpYGImp/D3mAbwwTWmW4ZfWfz5tbplrPbNr/M28MoT/2Q
dZK/Rk7RtozoXRP5dn5y1d8OV4cRrPm40j309QEsNXz5Hw0Nfk692CBUwRI+8LLQUk+yWIGhcWao
XbTG69BGRL669nlbQ7jinhtH0xWPnRGJYCzVxukFqrn+IxRPKRVwHHpCrfZE7tfNeyKnu284LqZI
xp9MHZzTJJq4XXkQN1BUxpP1SBg8qE6t16T0b7BpGyxdi7+DsSOqy9m1SHcQm3HFriQWeOleNqNn
ppt0hQ4oNKWfDuGouWgGGfI2f2JegxMWLRTtW1WJC2syjuXedGPW7f/306XRkCYuQSJBoxqe8WZf
GHqa/hlVdzy9WC9Xx8cy9UoujhklIivcHHn9Kzrpdjq6aL9hZlfQIZBP+hf/KCzgbW42JfSHeHxL
EZZMrwHUD7yS2Pq4SE8kCO6iwb/I/Uqre3bE6JWWsN8ne8BxzYtm5/c3ZuWIEoe7HJCsJJR58gfw
z3lLwmL5YGoMtpRf11LxlfSau2OUOUlBufC5DIWpxVXQSrKD3cLqedK13vPu/U+GMRU+9RWoS2uv
EqipDGRaZATe7hxvtWgcbfxvYvibKhDr8NfZEW0dTSvw8YVEpzWk66IHKDqD9Hy5RcDN9jT99chd
jpTuDGgb6ONMgDW5NGEmedII9SznYHzInZ21aVL560h4KA5gKJGh/UQrBDCzxTTSfFWWvpweiqW7
oGA0UP96nJOyQsD13/qhazB5rN7MhpV7iFr885EmJ6FHjDqxsozSQTyxZjuwqLS5gGMD/xE8pzHx
KgnNzWnJXqI39+p66HzwsAbR379PPtbp0MjcFjz70fGF1IHQhgIOwTEJS23B1FVftbnAt08MElDc
aJA9CwFwh2lG/D7xW5d8q/Co2a4AjiHRmi6RBVZs/OZcJX8ibVx0Skg+Wrtfg2YQuSBuzqExZbKv
4uq0Fs/Vk6zTDnMcO33ReX2hbhqoNOY0LwIaDlUO4t8ZudlTkAamo13OI4iZDvBbAli2E6emJrvO
rrsOpoiW3D10qxnK+b0wBgabK3qlk4pF6RWAblbif2lp6Z3aKxoVgTEpBeOb2hSqh+D0sIhZXOx1
cHiYP8HgfIq45QYhSmGSGoXK3O4gr6BzI5+ORjR0Ohue7Mkpl3cltfu21dnrhAr0H8/rqlsCqd00
TB4FlWBkpGY71HFPgUWbJm5u0wWloGXp8jjLVg7SIS6/m5Q8khgUBXSeVHjijWW2D9xqeGgRJCY0
o+5ituJsAiYR2CAjUbRPDNgcREb5tGZM94QTlEn/CINz0meYFqciOlSCiMT2yy64HTPP5Epg9vIh
7+QkFLBMfWbYvYD92sh6JAnr7WwDcuQYXrCEX/c+2Rp0kdPUHm1p2EyX9biffknBOnF9IbLsiBTk
5F0qauyXUCaz+a728jir3ZchdFTYGez8ZPiVDQ4H8rpYy2+8b2CKlOu/rcjMRYJ9vg5eu+7/R/iZ
8AhzRB4ICvI1u05RvGbmeBp/lubTL7BReCdCiko+jysChE73zM4zjkETFBCxQ1w4n0jOkGmY77QW
3XwNhldf19Cm9tC7qvNoEtm9UXNuFyVp3YmS1/zb2JwYmsUDwbpaGhOueebUYgeqibmbLOZON2Ut
etNSjHMqOBg1P/+mkmtZ1kLl/C7RH7xEzvPCdxBKTY+kX3j5yEwKvFyZqMKP8C2R+DKK3zkyPcDO
/UEtzi8ZCkmjMlnel3NDyMr06b9z88CtX9lQ6g463HaNI0YkViMtwBVE5Nt4S/V2sds8CqsdZi5T
RSjr6QYXN22puvMWUQgaJWCofytXTBpfka4AYTYLi0BrAO7ud7gc+lN8dMnaAc3/aal1H2go/U62
IXMxcRFWX3Wa8paUw1rEX8sbtGyyaj+/GkxDU7zoooXI1OgiwllBkZacmY+KwfmanijAYPoWPJiG
5q9J7TCrYuMT0D21mfnLxRjCTNZHAWi780fzIP32x9jyEOWHqD2te/nNUYLBN9ZlN2KlMPLJAWLd
juXggbohK+4LBwUDy4YeixVi1Fw1q/DeAMwb0IIjY7ZBa2KEugjXDV1WthFVDDEz+2/muO+/I95L
OjQIZK9hglNlBusJFdHGdSytbcNkDO+jcNFxydTd5vDEMkTWNmj9kY5PdE4JVjx+ek+08A2GWftx
s6hNt1RAARbImm62aOUSM+e2H/HRT8xEkKyjIcwD8A22oQzIsJLTLC9TrtWzrt9GPyTuYTdCKdoy
SxaJfxDXe7Yh5KeYeA/lqNq15OXAw2kLAjXh+XXt+z4LQ+/+Ls3Puv5rP8t96xNsa/eBJVq8ZKyV
vbMkgWfbCTQrb3AESo/ks525SbPO2GY/jJt6fQDIb48G6nr7PIUKnF6/4DFO9g1jGmfnJ/Kky1kh
9Ul5KmkGw/z4sevJ7qV1rFtTDrmcGBPb2J7pFCj7YL0t0jLmjsQwOXgBMMh2fqH11i1kQHJdk/gi
GWsSgP75L4h+/lKa4O8fmg0hJi2wXBkU5hGlMulDGbEYJuO9/X/wG70elnzlJGMboxf+Ggp24JAJ
2JUF84hu+3hIrfrs4U3r/7js9uwhBg72Rjz0H7mUb32RnlAbZi/zNT7irNgmm2AjTfdFYA1QWNFX
S8FL2lwE1qze7k5+Ruv/AY48eul7vMTFfIYFzZUvlo3CElzFzcqLc74q/ddV1DNh4mL6SsiQIuI8
s1w5UpZgRoJd1DyefnxCVmlOxJZZUsrVLdrKG4AMqyiDl64i2jnQJuSgHaLov+0JdEodfcQm2klQ
7ZV2NyLzFwddjGj2LSDEh/07tFreDIhtXXToU5RMZK6FvwHM9sRisz2g1Q4HWoCHFqSMKpXRk8hh
XRj5AtYWPQUo6XIhpnkuifPZq6oO2MGW9NPyc7w5jVcHBiUuhuKsVvI0miB2W1iOG34lFCR1nHvI
FW85xnojbluXFzpJyKJQEh72Ssn837jvHgNFYVjVkt7zadGDlislvsJLeLsJZKP3XkC62F6BSmQj
oq8NEXzf270B2j42gk7CE7UzW1pNHSVaCWvPDCenkBfRrloaYM6aFriuAivs2DYvFkE3tapUHu77
MFuQGtpIGfGWwzqcJsn4o9I2+HF1QDxhCwqjmLBKd6BJtdDLok4nwE3Ts4vhGryS79GT4a9leN/c
/j2jNLpUde/x8HoIektzq3PWyXjqLwE37iu7hIdgWC3+ae9+mt7U8bC/sUqSdgdd4927asUPxxJT
uVuprIoa09YP7NpySonEIyYkZKfGX4Nf4wqCh7WIk+kMm7f84lpYUr4IOnLxcJwP6j2SZCuikSQu
WCak23X67eQh4xq5qnzqdlkPT5OicrXEN2HTeYgiBs6MkJPpyc3hGrKL8m4j5JtqM9CeVIjqd7Pa
GSuvC4f+JeqMLUgZN5UrP6JT0x/rvy1zoOqlYjCWnlGEODAwyQAk/wJtqMu9kaiCe0XJDHa7ibIb
dwl1cjRmJTVfVlknkLeRGcHHOlWqGrN6Ts1j1wYPTgzFUCU8qfysLdfMbfwEqsAICgjW8NqY2EkV
2vvnnfcfr7hj2AKmg1OMLrAbJ8BG19EjwXxPObIumKUza7z5P2YVR3qIvdwMI6ASLgYDrOJAYgQe
PjvBFYoUDfxoB3abfyPJ6FT27UBaxqSlOeLc9xYuVow2z24R870Mz3sWDHUNgs/5k43UkjncT9U2
cR9wHZQl6l/LAVt+kCzlcbndXfCRNlO536nJPj1psI1U1cv9YI/dOnZEylwhAvYAo9giIt0s0E3T
25MFqdMSNwkse8g9O/D76mP3H/gl6dDXF5uTFR49QnZJZ4Yo4jcqgH676uD3a7c2bJnkGBfzXz5M
bD5hTFQhglP8sZyvaI2DkC8V+UsHffeHBxbMEgIboyMjHxsxLY2Q1O0l0zGLUhOOFI4AGXjiEjoz
RETpOPgyPdE9nxi9S4b7in2nw2+BcdnbJn6e9slAAUAXsZ3YEnt7ZFuJvcJPH7fkILSEKcBhMsYV
Y8RpWDu5PXOkyDP2vQtFeKKWuOMlcBWS2XBVG/m/cykqk0dTnCPp2hSHpP5agR5TCuXFzqip+JaB
ynXvzh5Uwdj6K69Egijf430PvnMz5sWhNuccUR4ntuBI6TDtjjYszc80DEgQamcEo2tBDIGC6qxM
xLxxjRs9RZ8pLG1AFMbwwiE+zVRiNfpJtvawSikFslCRFeT05LpOrd+Ug08n+p00OEIVbO8Rycw9
nFrxeiw/CDCiuZagUzR5Q3UOOZLtFl/cbjNv+4NJsHg7VNU0VHQr5Wf45hgFR8zQc/kGDl0N7hNN
Dktz3SUcf4UB+PCB8kvxLJWW/fbK0HBYseCu8ncpQ2iJAoK0f67oR1h7P4eMay29q860+3ezhSuH
qM6dZxABcCPLRRLOjrmWWejYR5TTYugkmbek1h5qAD211H7C9Z0boeg07En6ukMxyF2njllr3oyK
ACrYWtTy88L6MAzWDPlTBTFMWWEfWR7PE1cqnKy/w2w75bYJFBufmDnP8iBtLO2gvoeOEBWT4sOF
jYrLvYHK82uU3d25c65PnzfXNtuZOaf1k0JiCOsvos3/S9fFBLpIkFngoUAU5oPME5G+RchsD0GU
zNVOLaPszUELu30Qb5DoIUhpqNaXrwoEmBZeeiEntqlVhEzDWZ1UldRL3k1v3e5VI9e7e7vOt4eD
Hqz8h4Cuw2kmqMoXkPj3mlq4zI/ZS+qDQ5a9YGpX6k7Z7h3mQDb6s8B9YfG49kTO93X+YVlIIAYh
i9hwuJx/hs4ltQ1J+gHWb2Z+15L6uUxYj0v6csbli/iC+8lcg4t/Q2L+tyrdcOm+JMVtzwg44u+c
L8RSjVV9urlNd9Co4q6wpC9dfY0O+mubXA6egitKz0fpvqW1DHab/M2EhoMGaHO2pwraltdH8bSG
+484FsB1DqEP2ih6towLbsohPsOo7RZzxafEI1pVaAbRnwwPifn+YqSntYb2iYS3UUhh79XyXuzH
dwnuIaJhGzV3EgyzRNf+Wu6kreBsXxdUASCHIFkLHwXmkgcU3cH9nB7VLHdlyC5C0knMzZV1ymf1
s21vAnqMR1x/JiK+wJFbTI4cS80KV04ZsLqrRdAxJScpu5dwqgfSoFcOh/gJRSBF5LHJd+K19BEI
Xfff1tKYjolUXYvlOlAtrmPS6yUHS9Ef+hES6h+JoqWZbOTNs56pHneulwiSLZFLGH/90N1LrcEZ
MwXDTMltH27R0Bj5busWnBpHovoovhhpRoUDvan37a6XKL5mODVEGA4vJ9Q2VOzprtnYX2ZkJ8Mk
0MTYlUOSj4GjmxtLMHtRABnO9XIGrq/K9TlWa8atfhfxpMmedzbNR48n9N6J6Hj8Ti55gm46vhXw
3D2xHI7+pbgtdOK3fKAU3VEaL4pHmwFs4C+T6Mx4COzt6QsA0R4W/rJpdyO1Ekm8ONUcizptKZbd
mwWAKaShSUCdcGnEon2Lmuo0TWHALHe19FHjn/18Kw/FRfofw0wugEO2U/3XSJjUekWZJ5+T3NSv
Hi6j+RRv8aw00EFK4tp5wNcl0FK04EHR0k22v4BZiOghvbMc6A+WwwhcTDab9HkjyVh+jaDllei7
P6ZoYDnTjaX52+rMnXoush+ib3V/rGDX2l7tgkEp1K2C8jva4dtMR8K00Mz1qj/MRtsd3WPhUAOQ
fGKWQWiJXaIFpiWN7csgw+a0YV+Pe44Ch0/rFVqqkU8eNaA+G5I0zPYICwpd1TID2HqtlQet9z+I
I5S678UAW6k1avR2S7aCX0vS29dm6t5TjVJpt7TDk+/KUQMzJm5MuZDjLUG4xtRP40NUW+LUVQN5
ZJJ18Y3dnt4LXIjCQuVNhEt03zXidBG6NFpii7mdRXYkRgMlxpjxjByrIla0VC3+vGVBfMXQFCuc
rb3u+MEbP2vuC2FHQQMZhibm/YYKUPYT0K//ouB4cc8KM3JXfUGtPM5UAyCYSMeRE17YmBpuFyyb
uhu9bysB8AoKG/AFOMne8F4JQPsJYvRKuOF0yukhzzZiSwOXKsYm01/esG64QuJcJ+dTvgD2ilYw
mMIRNyvvjsmJNRJIS+vVjT/7mrrZFkqAA5ih+v1ydUAQvTk3vmjzzRHmfIgecn+H2MJ9G6vLeduy
G+rKT0LZekehmjRGe/rggyuWybavBQaISTzjPYOTPfBH9h2nd6qZGNvJPI2L1YvGOkf/7+qhmwRZ
o7h5RDbdVTdoc4Edne/yJbxziYkZRCiHj2EyPEp+vSSrobavpm/U5v5fVJko6KT/kOCO2V2bELSt
dqnvlSbqFqnhklDx1uAmFVOqNN0595MfMHMmQYA2zwfgfaGj115GLtFcbU25A+gdVRoIunLa/+vs
hGHoHj/zXArGGhLEJGuWxu+6WTPqGfVHlIedw/X6TWOz+KW/F17MEb+BKS4TehM+81/gYbrbqWcF
tK9LY9ifWnJlDS5IwFVaSOiuPNjiLsZMKl1ySBMQXURsc4+r3VfHc8Nz20QAtQtmzOk//o/44vIK
1iFcRLE5G9lLtsmUG/gZl1jzrl4TMt0Wz2iUPA0Y0PTA66RDPMe6ExvNG5q2TXGUqpktw0bQ4ngR
MhzFTxxgsKEqQ7Kh4qx0E+xmXXTzhwVO6yrKS7s1/lZjC3R3nD640U+XWKkPem3e410U0nySFyrq
A21Qhl+dDJCO2A2mqgmfr5q/f1xJusTRxcQgSE1Lm561hMFtBic1NQAv1fMR8ixoFcvI8GqUDeA2
MFbT23IPp3wOdX3X375j1q1isBNMzaYg4uC0lSueDAfKjvWw58fL/zFmhfxISAaaKFhx6ad5RThL
7QKiAl0b+Xs8ftaY9sXMTd51w2eNTCaT1MNtNNIWXtt0j4+uhUSz9DuUlH7CymcJH0wJr1PUXMUi
uPB9HBoFCIVu4+iJd8tpd6CPDrDxHpLAlPk/E0DieOgHc0NAV7RQ753Ks2k7iClA/CgyWdfT/dSb
GK7Au9MPzLDpDHyn7+JuSoIC5enBNuNkUpmnAIIUoad0/oWhOBwZLyyIQOJd53CzKaTkTxn8QIJl
UJyXoWjpb33cTSaZ2eUdNHrlOEz4Cgqd/bUHmbu8GsnPcxTYkxUNgepxgdvOOR1n39GGTTq+xsvZ
th4EbI623PflJ1/xMYK9j24kvAiwKaPGsf71t1xOqhMX7N80vjKVftHkJ+32khRQ74DIH55TVGzV
OiXXZ+nWnIfT8waFD31vx1VFS5+e7zoBX+C2MbP/lQN+W4UaZ/FJgt7i20Iyx89iUO8yeyhtTPU5
wr0KXY09YMTE/fyfSBXxYJZcf6TH9Qch/Rm3QNcxl7EtchcDCkhSKZsKnmMdm+EgNVwHiINcfAj2
xBS9x0A04IN0yKBxy+8nL4wyREDDpIRk2G/7dlZjGohTmoL7GC+0H/OrFbunc/O9g9G7PRoJe6aj
37EqbXgxsu1+6KOYWSfO0r5KX7Umi1vOL/C/TvcAHK+H6GhGZXk5PivlwOXKvj/iBBjaGx7EGK/Z
pgPTznJFNsZJc84bSpHkr8GBaN5tu4w0KBJmgIVTLufiwBDxM3xeqteuggmOntrY9l5qIMxBypRd
ls+GJP77l8DWBVK46lB3dBUL0cxuecGAUUpFn4mGODLHMETH1lr8oNyOaZ9rrthdeUI2avff4pVK
5ooIuwun5ga07RDXD20djqGBJwLyV1bKel8r5v82ffYfo61Vo1S28QbrVEV+342tgHl7FNOzw8fk
L9nwUT6kYtSR8Isq9ivIQO9zHMDi/s+5lYctx3ZnaZv6Xn/Uas374sHnl4wsVKHLlzQzKgIZcYWH
f8bz3NHD91P2d80Lh2GSGY9WUo2doQWI+8+h0jwz4kWHh3RzRGANoah3ki6nFk00UjULSf3UKylJ
YzPezhnarlskOy0ZIzR06BTmG8SOl9FUOQmQTKAZunBxG4fTLsMYe0S4FO5/JuSWk5ZpYRuLcJo3
F+fehspG4Z/zFYRRYdFvNnhgcqxTCo7VG8AVTI5LcdnShv0CMMoOlgiKYxc02XApA9/LM6hV6OAD
5oI9MmsJ162FZiLWCj/i1X3/D9KAX5Kh+1T0UKJxzGSwSFsCUeFeZRqq8tRJAAPu6T+2PbX0FHQy
DRBW2qc1jBUoYjXquT+yJ4tvV06gPeO259ZX3fYkUj5o6L29qRkPQxSXbeOQYtFKGQf1mANgmepW
XRBKI6EvS+v3fpbk+NDi4DZHs5mOUmJp6Mhmm11IKuSXMtULSW5uPL4F+68pG9GeffXatQQpKWnD
ewfFAE4HRBh8C4oa/lLQND68bBeuZwHtyJ0pf8EclxTYa9LxxgcpywXIuC3d4o0y7I96Q4ftOZCj
P/Wf3T7E8GgfXz+XtVLkrzaqybvtDcx23VxRE2YnpfIVy3R4pqQ8KccH8IqDLP8/apZJh6uysoiz
9qaWI5EvvMsCdeTEOPxrFVGeIAm8ZvIYLDI0j6VhFYF3rsQLx/FEZKBQ/+OpGkX/5i+uVP+oMNqt
D7Vp2iMofuuGrLJDv4xPgvl6N8F5RwZ++4UD7JYbslkKsMzGcMDNmXAhbAQs8z2qWrPn35lxCZVU
HlDXP7oEThuW/5pA/At1G1EFPIk1GLHkGKCwzJ8YHAtcSO51l/TqgxpHwVLiYIqBXT4nT8sbteGY
tF2ZT3nLnWy1dS/BeKzHnooj6xb4ehs3O9CvelKL5eZVo27FPALsrCSX9N9cGP3AaO5AfWWTXc12
S2eUj8AYW/Ke1GcOelZxBV9CtBUGwwXkGHX0bKmFr2Zrf01olgp4TmmFChhHGSOdCDTtUecuhCVf
1BM29wOSc3MQE6W+dUd5QT0CL9PYY7tz9E9pDbVvq8asQvBB6YvJvWpFB9PO2UbuTbjhuRq63xFI
uafMOk5iAQXlwZNicZzhylwt/hleNVBxXpb+tviVwOUlP8bKObGXYiRRvT8Nd8cVsZ27C+xxrH1Z
CO/v8MEoCplPQF/FJVfKQhEE1YqnVfKL1Usbab3Ls+cZz+h/gv8VyB66CPW9BuSJUK5OwZ6YFrts
cc4P/q82C9pJL72IrkpLpTqa//HjMoHDk/9RUuOzKr3DxSGQ8WGMrQJTvxOeds/4lr+WIkywgHfi
phoC4OPZjw/xsOrofUCUCQHcCkW+U0YnJx55IDLVOJma7Go5PvwVdFfyLuPbberAzOHib+Nc72y7
wNP+u3uo5+0HcYjw9S9PhG9FeHPuHEQQUmg7OsldO94e9xQT0rsABphZ3oHEmvuMEC5IBYJTW1Lv
b5zhsG9Akm4/tc7kbuvRdJqrNzlv4si88oQP74Tup7ZYkBwiZGZ1VOhljozrwRvyW7mV4y+IhZ5c
0ylHNCgUiJWe14It7B1UEV8R7eqg8erNmXTEU9EhZ0OfjfbZR28jHofhoL2rPfiy+xiBlBb2ceOA
pO2UrUjDMyVcVwAzT7EbSMtpVzTEDJ9BYSBdRxSwzz13zRPMti0RyoBt05lx2nn+cMSP8J5nzteX
teLKNehPWfH8gYBFZigUlvvIUMLedeJVMtHom9ZSXIRU4XgFn6W2jLJSB3A2aZNvhgy2n0sGdhkK
uQAqgqIt5Gn/sDSRGPLMQUd09FaEj/c2RQ0dWjW0Ibh2U9FQi8QTQ7pmwuNxvtg+5cC5XUgzzV4t
hNUIOJO/x0SDNA7guta9QZAK4fvnH90WBzg2l044iNRrTmmrN+HtAFyzaoGDTMWM6pd01kI+uTuY
WBxqGpYt3MI++Lth5BQelQBOLlQRuZvdLD97w4tUYdnOVoiEDxxa9sZh+VwCEqL8lQEYG7/ldTrv
5El12/f5+L6jo492TGYLcc6/bf5qP77S89Y58cZSIq7oL9MFQCFW3fIO4zTUK91DfPWuhJC/bEMz
5CLCn1V02/qtahcBUTTNSVB7vZmrX1BGFRH/Kp8qomXD7/j1hwtlevEQMy/s9EWVAGXEHfGXKQAf
K32r8akKopgn7Y3WjiyziGmRpcYSZmaE/+UdrbdWTRtrMNHasNkNUkqfR7P/unwln5nVCAirdsvx
CZfXqo9YQoJ3yfKUIX70lTkThWuqUKfIw2jtOcXNGQKfF8sQfk8oFGOxjGwzn+CuMDtLUHz5VFlh
dxQhaZCJqkcrNrPbkLEiMMQ0Ga+1ckWHM6M3tLBSVx06N5aFOkT/iqcIazo5ROb/z/2XQvWYzldi
mpf3OSktohLRUG5wEpNLH3oOmclcVyRCMo9FsXcMm6HkzecvXFSJFTBtv4UqddcsDGouoGfT0xcp
xPvBj4X3QhZ6qv3m00Rzv4aVqGDgL7uhxE2e4gwjmWGLgLujaeUlIo3jCDY5YEuzIEIUJkiztlLG
oPB5taGsqvPrgE9PhBjrxz4nXAziXb3EoY5nbkrYWkXoOfuccla3uWcDHRAE4ActhT2nsnFcw2o6
mVXYr0MFcKDRM+9c/elfUvAil4BTQFRmCPDiKwiT2KtL+sSHNjX8FGRPz/I+3H+EiulqVlVutK6v
ytGmjtIYUZR++A68QnvGJEf9ZHw0Sui+Y52uxY0+XNOe/Op0P9xb4UTnpOCB4jgP5i+k4PjwRv+j
eaANmTy2pmZOydfoNrtdVv4WL1rijDnxVKiTFmPu3CTsL+JPwfWlP721BVD9r7cEPjTdVdLj47EK
899f+Clh4MDuB3HhMRUFjyJFNb6tDscsG3xCpW3pR5c6/o+/51j0bh1litJHp3Km+Pcz27hod7ZE
WYqGKYYav9+5Sh/z4q2DgVzZmvn7OOVmlOSSUy47oX39pcgs+ep8cpwZDXeVcoK8pi7mfL99s9zq
+zfpLtKFkQPh5JJD0OCFCZdWBlf7MSNYVegvk++wlSMfjJH4Q27wqAo94UHKIp6loEsIzMYab3hw
X6A8D61jQe3DpdVgval4fLc9dZsXVDqkmhmDrk2psYwTZ849RI+GnLiw1FMpTJz1k3vP82EMsarp
sA3iist9Y9HIH94zmWKJi4Ff06vUwt8rMlOpK7dQ8FP+DyXSYzWwr+gvCLxVWzvU0zy+f0Zrwjcw
mr0fIeQkVRg0SttVTjILqikWH9SfUZhXuUI6nfIB+N7fH9UyyVPG4uCeEry0f7X8Gfb1cwunkZgv
fPnVL0pBUGh7nl23jgK2fr/ktd1FlNwDwQFwmzov42hro1caEIh5ETaVsqIjrj/oJ2s1oecvDcXM
hCN09cv9g8LImz/AB8LJe8oza2XbGkucNNJwoNVcnIyNpHhtNx5OfqPJKg3n4LoCblE/T/UFeZwU
LEXS1qzAI5pqtu3I8nQvSGPmYUACKXcb4kiQx+wqPbAX2E6cD3LX+3K7ozjwSaEl9YBlUQPsFD5q
+QVOnYbf2i9sfSiEQGD8s2waUIXJsY9FRFEXNtt+qQabGIlxB1sC23jOuMCOqlltrnIwLH+MtlH+
iUE1W1Hs4xW/I8cL9YGSdRzgog0DOqs4+XKLREDIcarVoKLDwhdNjPalB+EAz1hu5Qe5KQJHouoT
Ud7xaZL7L/RCJjPVt8pHzyvjL8y5/9kOgMqeUH4b4DJg7q6CENLlIED4JaTE/J5UmAx9nOqvU3BI
S8LNkqtpufKUqJXpoE85Qutl3xknJ/nHbusfa9oX6FthDEeirsVHQ2E1/hhkUBJztctkDw3UGiao
36p64iOUbq8fIrltHDOVj6OKykOkB3Pb6gUXTUuadzn3ODiiNDfQYuVhaaplFOrPICr+lGfIF31q
/ySBouS/icDvz896vW6WjqzRkpvlRdwQPRwefEUJIiJpJy6Bl/qeDYYwmccxa5mPqDq1Wds3uhYz
gorQj2rdqDDbqEbhicuWm5xvABzzx8icvKp9N+cw9IrQ0zkCEMf+ApqcOvam2U0cAds76Oyh/tWE
d7w1tQ4aWIvRVPH6XtO2ekIA/dRouAIzFzwtg5O1XOJ6XOoVHLXiSyax4JGP/1xy6/+upUUxum92
wy1SxqntdiXnDn3qVjmtMY+2SO0zg2KRMvkGYFGevVQEuk5S94W5EFUW0Na+YsAJa5mBkATftl/7
XRgked12HrWzZtSHZqBrkCqRlF2Uif7zglo5ZYb7o95pMv+sVldOXUDpmtJ1leKrN9+j7FquZeyp
3R3Sw1z6j2u8VHRSMFH0FfcYEJ+tGVrBumxmdCe1H/YHvxzmmHTKD0PcAP9ZriiDvgQjzN1G7SY6
5iecua/GbF1uBS1MVgwd3UgBUgpGaUeLIrDputSKup/ArcVArLiOQf0Z4IiQy+WgLAfIxUr0MS5v
/VyaUXoXTd2hM+Dp4yLlBqPis7zh4RWOstEIMJE/eTaqlHHALcZ5MKda4YSG/xrzJxUKhRfcnOoA
beIR4GYIkA3Pu8zi5K8c7+igpD0dwmqyLQW/zThwj7ByT/9u3kAwlYhxSFyGYnW0mOeHO0VsyGPU
EtDAS5XdSqLxOhJxAN02Kzdzsrnd5OKPqoJq/X/1bQd8o8VL4YP9b6V3THsp2LuMm+Yk7BxkheuQ
PmQGnD6A9fdjR0mGVSGKfWjPJ77aBcRXKSPnePvxK/rtfYKSheyes7+DFF171sQAEXQdh+w4b4zA
kPWFU/r+ZV3IWv3IdFQ2K7AhV+XxoEuJO8VKMGEla3knh0mpVK1BdjzD+uIoRC5934ug+o75L1iI
X89czbPMiDz0fFyb2eEdXkzHT0COqE09a+CYZnFu/0+u47qjH2aPyeDZ98l3bekmLJG73x+JLC5Q
9Z64cvXRz01CD6QOvUYvZ8mqrCa3dWxEUprK0O7e6HdMNz170KnFSqNQFk1GyXujsIM4+nRwyvNY
MC+WJm6ylz6Xhzjz/LHHWRDBIQaT8jdtYhxV4gTgcCfXJp5D3i4O9qzxaWreJjDYWVCP9zaGrIic
tkXVBp5HJuTeJDZdmACFtj/7ai3y6OV+DylgruCpb5jKTDvagQETlqPY11Ss7rlW8rlMsOO0dcBU
7JlUdAeHrdCf5HRm+j3Qvk9dqb0eR2bQbHeUd76e8lQpINBti3UEpnBGjkzIQT2RiOQkj7+qUWUY
EXFr7DI3y+3eise1nOEgTkny/6DNptQD8m5RPFO8mH7l+wRpYeOgzDE/B6/GL0BZdOJTtFr1q4wJ
Yy12jp84oRvkYGlpohg/PUlkD+8v0Fm/I0M0pTKBHZiZvV8pjx7CJ09e/R79IVSLQhK3qpdyrMuI
z9k7kSnu8jV0KifVsaVvAgWoEIyjGTzJBKSLxF7IFAmRG7s8kbldbUgilJNA8JCk0F5dMCseEauF
VhHXzk9KFpPzyjLnKiE3gcfYSOUdUabCpuxuCierB8jMHBS2Fxv2fAcAo5VBUV2HV2jUhAiMWkEk
mNRoiY+ma8WhPq2Iz1xRKlFxKqu9B2Am4ZPvVg4f0nl/AidedAShH3E728CINfzWWI6xC7arhn3J
yQ/LSojyMIJM5M/Fplou2fTIUGZvwgcL2GjT+XJhFbPfgHehWaGqEViJSBGv97VxZhzD6XMHz0md
tndYcB289E8dODbMhUbpYMJ8zip26dof+7TV2f7fnBK5g47LCKCYnBOSU5yVUIcUsEJ9/i5+6zx7
Xtqyt5VggaLxJM0W101SQJsqtKLseXm/BQh5zZNyiLX/+WjNRw2bh1dLAe5+ZOqIBoJgEqpR4aeh
MtMXHnw3tS27GDwtdtlNRk+kWx/VQM37EVLXg9H/pUU7Iv05fiedv3GXzJgsF2yxM0c0BltUXm8J
OTXL+bRWNKgq2aKzSrs0xq3i4wuntv1UoORHtd6Mvit31frBPRhUmto1xoQT4Lw/is6+1aI9GfTY
dZ1MbqkNxhYPifWCSrzVogLsR7T2gEFbfkwrG0OIU9C+S1GoNASDH3KsIOZQGAFlxc8XHrZgUsR9
HBikMdBUDGNhlcOqEnrmugAbxsQH0hWXaK4o3jAoAkrTLg4dFjcmjdHD2qnLyswFV3dJo+BNdPaS
Dz/u8dV7ay5h21y9n0TBLS43CoDGMbApXO/oi6zsLX8Je7/6mEDOr40bUHWIADw7e0WuU/zWGuEK
SSLAXbjx8LYBfpoK2KfHVAVC796mxdD2pAkV5McnG/u8ZnZl4YNUACNes9MJ8379GZRDLF7yAGw+
LY8hMNGQjpdp93TqAJAdHfoccdRA32T/GXWIu5m3BTsKjv67idwKFaCHmZxxmLP3IubI6fDgsy+F
GizajOwUyfEKIeCnPIzEVO9VzYQBxgJ47YAW3XIypKNiuA1K1sBhjIXtVdKiswGRIzQDxtVdGeqr
TidSQT3whMkJ9oplRh7q7oIjwPyqniHB5nsyBEzm4VJPlAfkeISMmoPCsU/unOXegdHeJqWl22pV
yHw1GgF08cCyMzno4/GdeVLv8qzV2zaVyJ1t8qOGTVEz+Yj/MNLR4oWL8g1pFdLwMXh2Pqvdj/9M
tG9sB3IrEX9f35HrXPZeKTMqldGXKzwbm/kdZ+Z8494BXzeOVQ1mcC6u2Tz4O5kcdQ1XerhLmVPY
lDwcXPsrXcel7wcmTJ4f1obdmsuPwRNlzSv5Ol7R6l364B4HeOtjWPIOQF34ADkh0JlbTMrWyXBt
KwQAXqXAfCWspiuFRaRrufcTaefQRKsoU4fK8/tnFb0IIFdxxMqGSgzjnwyfKdaUz3MBl6DUT7Qo
KGohIkoOy1BBrieDBC9K6jW8EaR9tV0Vp2zUAYe5erDgwNCxyTs0AG/zYqRxWZDTQDIy94xtE+zl
ksyIBcfaePoguEA1RKC0843tfZo/BkBKCtzne4AV/HuFL55q/Yf9uolFA4FggIMIpZuMJXj7ePTO
Adl+uvRJzM0MivkL373LsWLOwk0cyfMpIaVPo9nPWH8LWhYhoByIaVo8U7QDQ2u4ZuE3OKafjS4h
Clf4wykHvY0i1UD5zCrszWFNn5srb+1GQIhyGOcz7/L/UulvX7B29380DRkVHA052ILGICOriDUZ
t/nuWJs/ZxCDIMwru6a04RYnZu1pZCU3YcAf2hRA9zKWyrRn7RioUaXknsEFnpEDeFWikLwrCGY3
JA+xpZ/BO8bjyQ1oQDaXXjHXOkJgld54hlOnNyf8HyqFr/sHm7K8S8uXIdSR8049eK99FqbB7pKb
Q7XCDe0x6aRgUUbSQ552RlcuhytsKL5Y2tb2NvhscN2yxKcArcnj2SieOBQn3Cj3ZVwFV89NNBfJ
BnU80KwBm/7G8lEWg9ZtkEeN4HxynMoDZVTjI2WfEokw2XiCMasE2gU8V1W28rRzzhts8Gz683jy
NuTT9ElgIiRfM+ZQXFGKuZyEVmtcd4vMcdhvuq1Xrl/L3l8hPFWKdgKUlQuI8CyGeKGz/zczysoi
MVZmbyC3GropQOSTVX3dOSllg8mYQQmrRUwb2UOler6Rv3mCwtLC5bbEnMuMhFWt8XUL0LxyTK0H
fh1NQlBMJJ4H6KzEOpIYo2RYV+1JIQRWdtrYEOe/hS8pHTtmUFYKm/nWHvRBEFgx7WPrPXIUZVYO
MPP46kzWAEy6qe55qlh5q3JYZLdAMwOs6ERFvtkAsBBgDI5iQgPkA8hmK3OFDglyVWojZZJskKj9
mloOmYPGShWefkykkXVDVM5zMRZwMWnqQXHiz4TpUTthm2kkC5qOH8N54EA4dTcVmSyPbMb4XSDu
9j8QwKPHxFrsSY7P+lwWLrOroj0X0Vx7Y/ZbLMikBtvZlYGf1SVJYtA65sX5tq25EVn+Y+8WnS1F
DNAhbIEoVBNsciMf3ZAKrsoHb1dlYc3LqC8fnYEYpYyQGuH7M0AZdrLxNb44bh91nUolhFZG3kPn
SNdvO6NmCz5H/fPiXPSViG0pQcLX1SNI5hchTHuB3XGUHpmvYFZVPxl8Ca9gwEFjZYIYrCNSWhx4
YfvMzF+2tXCFJgRxqiS3I3yNO67/FOS43RxPOgYSDC9vVRXIhxFip8hhKvbqbRNagx3QakwtLhXc
NhU4hD4orZpODvp64mVU/qmc6rKP8DhE7Nybb11jvr1p58nTbgKmn7+sfJVvAJ5bnKr6S5SWOs0F
eO9YONI9GiV8uHG3AQ0J5QXC1Wftlj6868awwLn09oH+x9e80ofA8SJ+ghU945GAMhYufttgKBmx
iX6EdpFTE4yslC7Y/JZ6j9HEQcGbPuTB4wVZWqrFInSYNMKQDtknY3q+gJYbIEjx10AqS6tTudO9
79VHpAsOyKg3HuJCWuKwaLQx81nnqRcwnyAoe5QOol+B2+ZFCK14N1YD+H5vJfn0h4ajznIt7nvC
PStSfnmvxtjBnIQmhPEpuhXK5qWwpEkChS0PswyLqZw2Wm3nVRIGqy8KLrnFV7H1WbRD2T/wUYGv
W1Ft3+TRWUA1p7wYowX1lOIMsRHxsxnffDLG76RhwtD7JuFO5FurPH9KZ5TLi5Ui3So/cQyWq+Of
2ROOEFyrG7N0MBnAEgscNulclpCmJJ7JQxz9ltrQ3kiXaqERrbu5y9lOY46APGjcQt8958KyLxoJ
4rYQQcGJAaVLeFOdgWprKw7fBFCR4hrbq9XLK18xennu6mc30O+VgXmmx+9hCwTipd5DWilfLu/R
OLj4h5pi6WJF4oQmcOgTUlQLnW+PYZ01pfJlKdh0SXXrBgSX7YsSF09K5GJsyLFnXjwT9huO6De1
UDmiXkrgMIPqPkYIuoEXw2gB2s0TpWENmKY4aQwRBmewhFgjDqDiYxRV0bDa9OgLHr8hG1wdse3v
6UTWcsorC9Q6s2ZhSwBMztY/vWG6a/LVuF1hBwjgWnAA8CCmiL2F+SYn7wp+C+VTqHEmij+Pd9vQ
wwyFJTVo9B1YDjYvMWuyXbvbUprxgXWYONO2Km1I8pd2jDChcDOPjnGTTRA5sIQ6v82gcs8JXKH5
RvnTwmPf4o+jxwwy6+AUhF6VOaLdM1ZdZqZN3sZ7Fwm4R6zAmyCg1e8ABD27nsUxblQ9Q5h61pI8
vFwbqWQ6toyrBRiZXKzXAYrFRt91RGWrMnK8wg0px4AydcxAIndLtnVbbIZ76Rym5mjM4Dnh3hGb
wD/7XmqWHbILrX2BC1tiYbbnTm2iPZq858WMr13uKMlgB5sIY+FNrMx1bfHxHws600eV9v1TXaeR
vetUvWS3n/y58G3+LJjTQR1pmViRBJX7qtkrleaKIqSKHOCSNIMMjuMTQnVXGUymSnwkheDLc1Sf
bnaHsuPOSxdyu4XC7i0wCMt2ynu9IPudrHqkWuWNcwdkqXRC34Rslkxcs0YPX5bU2ixpG1N9dzyC
rP1ExPcjzmoNyDFjEgDjZPWD/9Ljh2A2MDb43yWGAuJ4PWG/n8kW7+ETsSgTNkO4naM/2I53dXMk
rsfhdG+IrgUBuoLUv5S/OtGZCovRym7IR2y8SKBKqOGayvslzSUbz/h3+NsgX3OSxl/j55mpJIgB
DacAe23L36NtmdtKZFIWCa/pn7+Cp7445kX/wrp0ApR6SqRFGITJn9gL1k/jEFP5itvxZDuM3S5E
+aQ4jdFHBr8/CmkCDdbgVK56LAci9tuwwmNdlfllv4e9yYtHVrg+vZtshrq+y34A0DEsM0B4fh+/
43oiZppVYsx3DvXx3z707zydpdcSkVMItydz1WUdzP1W5iFJnW+sr2ZWpW8vgBEAY7LOyAZ807hj
JBtyFymkxRFes/Ud5HGiTlR3Kp8P3IpIEsff8awOeThMBEBcPGjg5CEpTVpwsCXE8LoQkURt/WNh
WTl6YO4pMgXdUWJfNEkvCVPbWdizlaSQHeRFvEr6hclJVbAY2py0fIZrZXSpgXKIn9gJlaFCI9MY
zHjCGeDJfI7SjEmZRYnkhxSeG9St4AwTqzbhD+JpLnzTa58+8iXp2r1P6fxbl9jKC35eO1yphJiU
kr5/J1Tw+Xhi5MQWV2pfzvrw/UHw05O8APNcaznaaI6i1ANhDPZTuM1DrPvTkLiQXsvx7pHRF2T5
OS3sfzV5hKYM0eawjEyCznF8Uaji5etQtJcwjyoYtgcFqzHe/8OR62JsJ5cNXtRKqQ0feg6L3bZP
DQOUvxaBoMzMq4Avm4feuf4YtdKvnhkRnJuDVUovB3MV6h0IvVQDx4OnXTu/HaRRnjoNJdEoChbX
QCCIQRU89eRkR4Zl4M1iltoB1tWHGL8a1NsNkHMfI/3/SID9vR13eT20OcTkYdlMdVa5WZqpq0z9
MKktf76W+KbaPrOXZroON/vktQAe44/cWDduKW0W5Q8+Dpfl3RKH0zX7yoOyJ1KwCaiIR4U+QNlb
YNBHBgjwYm4IGnasWqxahddey0TSnNs0TZav0RQAT29A1Jk5bPZUgQWlW/3DsMODEpbO0lIMq28o
dUDh8Pc/C7VpdUx/BJHZ0Uwm9Y1G+Mb9Cnr2w72s6Nk75+glsAt40iShs2LA5Noqbd0AyH11e62p
2x15I+V7t6r7W5VuDlPMQp29l1R2uNnEvHU5eIqwxBO+pn2Wg3sSRrysFVd+atDmCTZgGA2rG+XP
y0uu9pTSE55lioQ3kWDhAPFGOAVlxBtHKrfWRxZcFSduPz9NWDt5W/ZS6VH4B/oTOdVDk+ONYlSf
l5smRIDvZ9/8qhHvv7r3D0V+6mloS0w0p8ZX3JLJuF9SdskjtQMXDnMLk6+PkF5deYOiXuFWmHwN
qJRX6mDv/qhKeq1v+xxVQ4DNNr0dYwNWZpQ+LfgKsr31TrO7CK0PVQiDDoA+UCu4gedfq0pO+WuS
COatRLQKrJOr5NbmaYjh5TxYpTLr4fdv5an13O66ZNC/pBv6UuTlT6ZOtfZqD3PwEu0gV6d56yHj
b3opibifcMaNCkiD6rF0RUcDoKSWhcbj+l8CJEZXTBeXkHqFmP0cJxl4Wr2lGf/MA65wPLWXZA4j
EV16hEJd/GO43rsBvfZbm4euPALkcEzf1PW5aCbQ8IiNrYF2+OCuNP/DZQIxJck9uM2eZ6TkOZTZ
ZE4w553BDadMoffwK65A9tbHiybbEocGwyfhNkYaKjgfgEP9Z8+vP4FIEvRafjRkQDV5oYbIOZUZ
SqUkOLem8mdVYI2qBvUQ3BpCmRebnPG4wZvTPo7hNAZf3zWOYHeTys9RsvUQQguSxO82gICleQyj
3lUD1+BQnPr0wOpDDa4qzrlHn1chYRmPge12WujRRNGjR1lQzis5qX0hwQnGTphKi66fqFoyZW8x
tJkVxUKFxWPM1yMRgP5bLVS/43+0/QPVzcyQLgYvaZ3VGnC03yrAaeXWU/VoHrEG6Z8pY1A3Kh64
Y/yirJgsADACRmjzNNWUKq0/gda2RWRLVTzkZIHVRLWG2ey4OVi38Q2hoUA+PNHJlkTUZXyBT6Dx
5PVen0m2M5Jt7apif3Px7fo5oN7ASrnv+AvTG7Gp3Qq74O0R/Yi38Tpw/Ymo+/GHrYTTn6h5j5Qx
jONM+3IOChgB3rMM1h83pADPAsvvorNYTHUp+cMntDquq4mhF6LQE66SaAe8BBY+X4juCWeYgZvW
oAkN+qzEu6JgL3QIG2lcFc4g47VNBOfEXJ108DyoBlrlzmd5aGTsX2CkiT9W+EIUTHPtfyY9oByi
NUSmFU2WQHXqcmpUyRx4dqEcS//bYRwfz/TS/lJ5RyR8OJZgaRaK5uceN7swGSf094wdg6B5+vi2
m/59I2S1Xpu1ugEHqhdEK1VTYpvlUHPkfF0TaRiIxMQI2p/3gjRVextD2ae7sAR9YLsZZ5FRb0Pu
c/vQMdNtGmWzwzciKIatoutEupeuEa6HredqrWczkn0aywdy9Xz+Mzwh3+dg0gA2zi0VLd+zUJ63
zi+CTh7RhS94bjY5XxfY8fXczOcrOKZdAD3bA8v8pdStm0OZh1O6RfjhbnmAa53X9z+QIQBawN3S
j7RDmokqd1rKG0xid0VkaNhgCoZyfnh0SJDFLzRN0DE5qyBFaXsBOh0zkE29IObPr+f2hH9JNVzA
tBpDA1nY34xn/LUHrpqN1CZb4uIqx/SfoWpQuR3pglyL1k6Yxa0mzwe+R3HN/Rj4z95IGZNDP/W/
/UIp/XJENXKy5XiN4MCVfSOBgYpcSLhpkL6NozlO6G1rtVx71kzJ9/8HZIMCivra6/zYAuhAllr5
VDn/RPvg+hDJDxJZ9LJAaD+ukkevK+0HT6EJ/CK/l0wd+Ac902KKuxTp4HIIga9tCedG3b4YtKeC
fBKXanbUyG11DidWM8mro98tF5wUbeFH2LMVzRLxMEDwezKef26KmFGkqWsUZ4eIQwRKAdXl8y11
vXA6o3j8ipZQrxRe+Eg5+4fYRnhUrV+1ZDqltbSS4UVxrRcDL+5bC+n2AXkWrgF2GJsVfxXrkVGN
lWUIaxpimwsL8FSp3L6KqtsuBpI1Kc0B+UPMFkyoHw3uqMgR7tCuDSsk134g5xApFhnE+3HQL5zZ
T8S3QCaHhR84nQqqM/6FNeHVtZoBkbxiyE1vsnHMlCXEanhYpjuKIiD7ggBXORTmjVu3UxshY9PF
wj8cw6NRs845gX26cl8UVNKdHxJO2DIzCCO6kX1TNjWckEQyKjUewcxCLtxw6Z1KrYN22ZHCPSwE
p5MbHqT0uTKfE8VpyODJLiChpej3dpCa38tW5pzPr1JOMBaKOHmY05OqRKynQiRxHz12MYVhFzQ4
NSkh1CO3a2go3VYmqpPhbOig8stoq5Ob9mzbQQ2eYR24CrZ8fFKso+fepb5Ld7hUROT4KNDRjUQx
jjeuuVEEryLpa+DWLbP1CK0FUkGq7qrOR3tQpcAV9YhxaG9cS/rEtUAZ57Xqs2CEi/vlDp8u7d52
qjNTSoImgqHySgjYf+i8RLVlwgJ0p5hgc5qlnAn50oSxaQvsqIaY/IPJnrJg66ArNmotvUmDu+zS
9adJepC+dGgNo4PkFRbZVOWR6t3rpCoC7S2xRh6abhc70i/gGGS2wcoM0QvnT5rVzNw3+XJjVysH
qY/7xw8WjzHaE8mGYqOI/D7tnWjS4T67de6FY2ykyR1Knve8GkrG40TnbTCi7xIc0UeOWnuO2JPv
FdWYxKdy1CxvYsmGCBPxLLeiwkNcMyx1LpfLnnc4iuu4htWlLTj9gI5XWAXB9F28v67odHyuuA/X
AisUuOuTZnRC3aCkSOcRoA1SQ0p99bsUI3kJclsvvFJ4w1yx3TEdpZnF/cvFt3rkuC78Fy+74Rnv
ubk5Yc75ZMN7k6qTxnoPQ5Lm/QPd3KujQSjk3/u5ODSvIl3wsfpfL34Mccy68MvVdZggOC0kTMLC
Zdhsk6LEsmYp868lsEuQjymc40sN+iWE4PkWwj9OqHgY+rjfrR+6P8Qtm813g3VR0/r/oCsH9rwf
tOyUmoqBL6rPUN1rVTgd2YMB3foVJgwNJUlnhRal9n3WSxmdLGGen+zQfx9YpCbCh9pB00rnBaFj
GbODXyHVQ/7lNB5YoapUe+g/ESVbn+C/S+ZwIhVz8j8xkrk3xdXFZ4TwygsRQ63lA+RtSv1vWtwk
qO/z6/PgTzn33Hr90RZ6GIKihBfOvSM7LzdnUMgfJb5+BSnqkMuLeebQWIWXWmMslxiulj/ghIp/
UpSBRmOFmdUZ+zzhbWVZMcYTlorDfIIjpB0aMwn/qo4mBb5SQnvHEidVYkkkt2yMh+2072soXm5e
CwDNB0ECi/sVTQzw4wVupdFiHGNJ+OxtZO2lBFRSIy/XcP1fUmzrS6TRkuJpaDo3B29nHdeOfvHi
BLjBUahOiRoNDKZNLVrM9Ocz04njDflM0PHqrQe2FQgCOjXYPAJv12fOj32wqH5H2Th41T/TrZOO
GHYFZkY5ZRmli0dqDdPP21Mmk5dyxKPCxOyWCaQggP8H4AQDD+pry/SOHZ5kwKqnZCw+LU52oZBr
HKnE5hBxMYCBuD9ORcskcesAwW5ROZZb3zexZKNRl7Q5AH46ONHz5vr4HgSG6wfAtcDzZ2kmHlA5
/tIptuvJe8KUVTeV+vgffT7YNZKFqZ8hapEH0m78o2bBlO/vCHLzhsju9blCDAnxcJxF0NojZNtt
QCBm5kVgmm9rMAoBRngvgtRP4smeAnQqlUsRksc1Gzo4A3Tda+nsygIHyEzF53+ZHVeAPoRs00F4
XIqXG9vTKSVMr5s8C9NpnYo4ak8Lo8YpKZFKCMXUnqDMunY5RuMMwFREKy4KLCKFSLAvNMkNCBKd
stCRO8xJ/I1e2sOUChTkcJf8M1g/ll9guXE/ubrhLHy29O90kZ1zNab60BWpJSRTeEINRPitFL52
NVyrujAnYRQr2WCBLBggM2rC0Q8N83DNAciBtuUy971C3MX+HYaQpINgJF2P9MIvHhLJgy/XMVhb
eDk7S9iBtsyxs1+qs/aVwhGM/BTKcZ7MOSEMS5b++Jhiu5t2X/QqgRUlYrVzGsxcAGK6vcv85RNo
9zRSMJiwWpjRKOeud+bch3S4XfnTmGZzxT10QFgGvIfohwFywHj4Pv+TqbBTz4r+CnU4sUKT0CXl
5Z4BJZlr1KeANsxEOH9t8EmhJxRMh9x4UGOpS0f3B0gCmQKra6O3aLHKDvRUvZQ2KoIFsD0KM0jp
lW4FBvM76noylamuw7ECIsvaPBZaJdjfaCFA6A9Ff+6tsWywZQGMTWI8+TzH36nqcWwapO7V5t4m
TmLbW8bjCK5ai6zo68gcPh3bWXQRt3/fP3J69XrAbRA+oc3Qxp41tSZABmfgMyY+54+6Mawt++4V
/If7+H8+2mBOlT584wn1sjowUyMo14jox5XslMAfln0klnzGk4mb3bNMznF/170oh0ooIeJCFpk9
s4Z6fgH7ALn3+mzof8aaX0cp0NyIYCie+mPrpp6xJbKnQWcJ/A3nD0r/FjuR0kTlVctRmKYEn+m+
L0i8FswyuPINWU/ZU6Acr+wE4gpGQWv9IyJsDu704KChSma6gMBnZnBsweQnJvlnyH+saQc3ehTK
/DyPvRGFbBvRXqlg6xxD2/BdVmHLExBpwA2WTIQT1RcHaZMUoGANTGp3SUVQwX68wWzcrRGA/PMX
RoWiJmWfrvQSzyM/wIcoALFe/9J3A4tHWmTy183FVLETW6i+JP1DF8VQAx52u35azRxZ8iR4jnZE
es58iVfudVxc/7o0re4B/U8tWOkq0DpZc7fOnF3bxfyCR0f4hp3O2PpjcvtLlpzSyjltURGCiyZZ
H5wHFOClosUrKF9E01d7SZEYL0HuPybyIYW8RDfFF4jBfvjKT3kFO9r3OPL3xKEkkjsc/nBQnA1x
dYJXKUmDb+djnEaoUNy0nn4XDUD96oAPkoBWGzOeK4XxKlvgG9SQIQV6mQwtPWl9XUlx1YAPEzr5
bj6JTlgo3J4Tl516bFsqIdVaY7Zv3CUbtpq4KWWdOKr7vQDrkcpIxs/EycDH9f84niKJMrUNPEs3
PJw0c843Fk8BKKAABdg83/29IogPkFqGHAqcAxfHp7U6p4rQ/1dKsctfyoPMsASttXSAB5K2/YeO
ddr92rlcLB242rHmbjl7cM+I+TfEsYA04YXMUNBOZyp0UDZBRLquV0t7Kpk1Nvgx82kE9Dm51faP
TW8Mtu67w2TvQuxfJijITn5FKd0sS58sf+eATjaIwODXRMMNsVwyd2NkRrYcSOWy7Vr+L1HMtneJ
k+KV7TsT2SSLWv3I2sVbeiOptn1GWkyH7D7slKoSXZ9B77syPqsp5Hnq9vzhKPhwFaCdP+tMZP1N
0OR8RLccIkmPwIVGf9I0J7pqdukHjrlAt0C/quhk4HU9dysX29c4QuedwsbQ8AR2PW32g3IrnGSM
A5Fb84SVceZ2I7kE5F3QKpuYFYib4jNbN517LsdD25vgIV1C4+dex3hxOBp23TwPsAj5VHI2aX3K
LcAyS4E5ZcguHM8vOH6mCGle/A391XppJ/ZA6zqjEJ9KLUvOkYQyoPAGfuLCvjIZYYLwJCJKeLnf
VcNQwKgYwBXXDkieddyILPFpGWNO+SGoNHrnpNruPVPBGjugLb9bnIJ/cFBzq4+wZ5CrpD9lR5fW
Dxyvxz4RlsDug6Z27lCNlBsKfso7GZL15Ctp0pz/7L1VFYVUgvhElbmrylCpDEsZE3o5qXsT6p2l
xeXhL72acu6cwj7Ym5q0r55612vOODpGEqVRz7sDcRMO/gE00a4cRcVZakTnLpdumO2QxkHP4SKD
xTW6haTe+KXjEu6QbHkjeyVU2nMsVHmojHb+XzeiggA91BO0LuNB8ZsRGmh3QlgdCl7PczvvGpQW
mlSnJw5ICZbJyK89UHB98WMXkLsapAIDSDivYwsz5TCFSwF7A3LkNbQvcSec0fEy1qUeGcNhEXCb
wg1gQmPdXhHZI4yqTSmbgm4uM6lKejPz95rpHKkbN9U8S+yDDvgCG9MkHInvWwevtFxMilrHrdPh
ItAfAnnYYYqrSIFB0cHqfzkEWW5Knuv5jz5ByMjOBEgNqAC/rP9XI2OYLVog+JxOXgvH3Ckk1DKR
ZN40KBCDuKGD8+ztkVtR4+ioGxrAuw5nG4yolSBAwa5Jm99ZJLWr+TjTtzq4dy/TmPnaepm0F+iF
i2NuwiM0aBHf1QNo0tpTYEUTPyECiPbjUYzAaDXkKrmSf90xVUCG0TLnVG1WUm3bUyfXJmS4MXLv
4K8418WyIOxdRxvr+RsxM2rnqLmIqgP7VaDVssGzEtOpEl8q/bQ1ZLfQHs3Q9y3wopxv4OwocyfY
OA5EuIPQx6SEID/8erkVidwy39Bid9qT8pL8c5vNlJ2BD/XVmJWWu/ksqobtU2qxsUvFVvRbMqyP
sDGLXKVdii4u6S/61HajTm/FhxnEKgXej7XJeHjMGCKcJVAyuIi+UzK8+jPsp1xC9aCDZUJCbkHi
cSlPAB9sotxRxGYDPtjBbHbEXWQ3VvVnmbXmVvUlGcLluufnH4yaXqvH+J0Cmu92ICk4XRcbbhwm
75TAAR582wSRbmWdgVYGqPLJKWwFxYUQkYmz8Qrh+f/9pGrBuky7JFuzU9+3uXu8dG59TZLpy9O8
+V3H/nEeDXfrkqcV7TuyEu6QlitAXtayQj0U+bx1zReKbAEKBae1no88t+ZcG2lbIsMxma0tsMqE
MXoPxTejdLPdTGG8zE7lIAX4RLb9xo1NyTnZlX3QmCdxG+wYTlu+UZN1ZUbR1rv2j0sDgwEwHN8o
a4zxXSJnXMmcSfqYVmQASJ6/v7U1j2C7dsQtupRIVB3CL/iZ/CtmWvKytmibMLjgFoc/PjsagFCz
UT9+2RxqURK+y2lJMV+zOfhm6m+DAIVq4en2HP8EXRW9t+Qtwh6A1d80SdSw7lGCH115oQ016smI
r53mdy0/lZ4z+xYPhyekAZxTNJVWPvwzXOK/XZdWs3YzCd/IoE06lSytO1+8QjgwFYFVJZxsXkLG
PWi8m6/qRWskuzU7FSYsdDiKFxSqVROEKN5ER1Vthw9Y1+HiDXW95ibJBIhS3jXHmpc6jeX/bQ+N
hFH+GOEndHkNt36pFGwyREcqerFvvbvfKuX4kqoLcflS2gw89XnSd0mylfREAFXRgqb0xMa+n2Fx
LchypyV4jx3C9xBcpe+XVYoP8r4DiYQ3RB1oTXw9gphte9MIlt+71gWpTxn5jG6Yxd+zl4QYmgnO
qBwGzACvJwPXhk3zaKlJvnZ+iut+YMutwLcgE29G1Od7Mu9W4RfnAcBF8SFfbe+u4RVSZXc75ECn
Rxy0Zw6zKtPhzU6Vfg6o/T+ErUPvO9+SiVReGL69PmkhPn3I40IpmP8WsfO81NWRWHAI5CML6szV
rS/JLUBk+3aWtZ5XIc/rk21JKFyjQZCqcz0SY8MgbFRqEJKToHbxESZcVV6seVB9pPFxBjAlupAn
aJuUAAwn9oGuI4UyOTbQGA7+j00GLqEhJgb+x4kXXwGtXO6dZGH4wpJaz85NbBxsdSAE5UNSGRIQ
E0OlIfOpmPnt3tciRKRbKY/sYiCHZ3wkMzuaKpBH3o53mWugbe3Qnz8Bn52E3WvqLqclZfLEwShC
PPJ0n7UWmarK4VuSXBeGdsG8RqRBDVyJJyGsQQWyMZtvnPsqw+WL2nKbfipydzo+UY/iSk6ZKBcv
7cMtiekgfK44FrmwS8bZkpHcw67WrznjWjPVwrT7dndkDAF/b807oB8If+GWPP5TLrQYYrEeIJmL
sriCluM0gM9xNc0qXT7DSyB6a4GJ7WSXUFB8UIdfXrfm7xPy8/kxyYORh8D9RdtC0s8Rji05edoI
l4nxR0ZijzrUt2ioeb2KBoJVbn587JEhr2IxcFCOd7QrJ6iekM3NDhhde2ccXCgTuIKp/qL7yKic
iTwCpFRje7L5jkWnx/NUDeREl8EpoyunHzR2OZUlH7/VKGsGSPZPIL1yASWKLS1paH4aSkwshwS1
OTdIIQe8wz8B1SbAVqfQY6q3w1eA7tlVfzEpVY9ypLNijGOYaI09/VZkzhzB31u1soTL/eZeMhHq
uCETU7lXIQu+A1jSxtWApGuW8JAaUCwkd6kkQUkcWuVmOjqWoCZSXgJEhGtTpcpmc9Eiwg3NR5No
6Q/FoorSsqjuFCvvrXvA/hqkwAEX33TdcB9YHL5EAwXMvsaTd1tqNx8CCh2FjY6U9+YYeUViQHNL
pEPucGKKkLGLV9Ni1OdYWezcwxE5ytnDJkkfZceaRzBAPreapAGb/eAdsGaRsZZtsjtRaEHvM3z+
n2b/lkzDUgTQA730nOnyHo4PUezQRTLK1/6aDYNnUyG4XhriU0Zp5K2GyqSFV8TdTn4+aob3Femu
p2xtQfYM7U2Cboycj3zb66R0aXthW0MknNNA9KXfZ/vZI2lJ8ajiS3vwPw7YCyb90flSvS4l7jRy
Mo5Xqo2bEwi2WvfD+UYwv47ItO7KzckTHKX/3uj2m8PBmuIa1ndwEVqO5NQVrYnZPpco7fwguV6R
nx6E/kTb1mvzxy8tkVe5PVZ/gZ0DqTVN1p5EsvASQJ4bxML2OT/RvoAkzTLpelnFpnokkMwc7Z+3
rKznDUk+e/ukHu09U6zUe5FotAnsHKrOWR19WH+fZ4MLOD0OuLdFR7GKDTfgimNy796c6pInHPvp
/2sM5rkhyp0BM6g3XGjL5e1puNR/q1rfcYlAcZgKl5mRkeY9HwwTsWZdBH2cL6xa29JK/BJbuup3
nOqY1lIED8IXFW2B33qWmI7WAE4gvMcrZIGYEopDZ1mX0JKB2wSe/4GuobQfeTXrQfKWeoMZfVXi
k+iSk5l7Ztw585HX6ij6sbEuMYCBMBwoa1+vfHp9WQLx1q5pIqgtgHU0mZ0xlaKRCUB3u8q3HuSx
p5EU1RWPl/YZrIJzskCIv0PpBrHvx+KBTis3kIeDeGDmNYXtWVQfm/IacWFjU5zavJ2V35JalaTG
EyuGQpkvsiiqDIcHMP4YcSllESLC1iE7+G1uFbW5ja/G/CUhhkM0IaUmmKFzyEAu33Nv+N/X9OYQ
iKwgX8fbP7NXlDTgK2xo16O7BaIv38M7CkCxiT6YdcXCGvFyPbPQgxWZWQMm3MUhjMecTncCeLdN
cDlpBxwbM99LysSAdZbdQEBivTW9YGgGXGevP0PMRXrUdGLidA9cb9nCWM1/pJNjQYxUnkVT6t/d
L+ysz61P4Cc2lUIDe18tDyDCLVJneszcp+Qfad7lpEO/W9LcBlBytO4BGoJEGiqYV35UJQBMt22J
4OzBxcYLIiKcAWfpnPmISAaRdkl1jhBjHKQm0hscPxJ9e97xuGUpuKLONKGheSTcppnvqObDilqH
4Jz4tpDiQ53PIMKsJH6lLfmLvPuXmwaoUXvL+lKqgtjRU1ZV6ZAgwVnvl83dR6gS6aI8/gjR/hhe
pXPg+ZT/egFvnhXHRv4ynbTEyrSCg1FRVHGuzpSdC5qlp9PaipfdqEBqSjk6WLmuXmOdukrHhpSV
wz+TZ5nsB4D+JQ9NradP4JS8zi4AnJ36EfEATxx/2GVjE9VlWvG2iOYJsuaX88mg68DaFFv3YBoN
vvZB6VSRSBJVR00kvCpocjb9vZ7otAKsqnbCNoGVU4S7PEsgLs5KCCKoUP10jMvbn0PIDaTECS+8
Pn6PQnLPcMQHN14oSFjzB+OkOgcMHuR4yAkQvBtD9dGyx3XGWkei9VOemDqaNWIv6QZLZndBJy/N
mWAVJvuyQbrJqA6aCjZIVYKqXlb3nyRPLXvIsOU82YFqr7edApwL5/GzNST3oVc+4kEBJM2eWq0P
b6T6g0Wc1u6SnTHXHzp3p18YDQKXM8I/4zePCwSkbm+ChSS2GeL28iuieXa0xgyYkVGWzUSbxHwV
jl8WwK3qdhTW5L/NKs2enkAvnEa4sFrTTgxKFq8r/zslVClR8htivbeO+24vJfx+ZzubgqXXszvt
ZfVs8YE8G7aRNp67Hxx3gGN7Dr9vaQy2kHEm2W6gF4Oktucrsh0648lGxfwTYyWOftMHDgH4XVRL
55wGiICWyH+MlmCBPEWnQ/rpmSKIpQbdu7WF0NH8HjoJu95r715AMcvG6qxSuslJDpwBa2iR0iCl
f4dTPOY5i6vV11iriSRh83kgPhFr9XUyEZcPIanmOVUIIefU+uPxfMPrIQg+I+8+e+SXpieNej34
76hLosgFJ81QFvTFMyRn3kTjd1mahYIAjbkEHc0wF6KTc5Yk0bIaE85Pbht+W25nEksRVbFvCTrz
oSbs2899cWAmQvFl0vneay1wIqeARM8bOPofahD5pIB9FYM568qggzg29OegaEJcyy12wzkxeS9f
A5M118yFqYg8tkhskR81AlxlGWxA0olsQA0iP+2OncNYmqyx6KOVBT6YVJSO1YhdsmZviq4y8F9v
BcyelhpKcSB8jmxg8dVmwuUfMWmo1hUb01JJ3ug6Dp14gpTHfGI4rf2dd681QG7SfaC0aYB15TLa
sTBNSc7F/C5YWjZODU4Om7OfVOu6HJ6s0yJ6ml13amd4xc545D5eKL6HmRXCfJIRfKgZgJI8s/M8
RKI9BrsdQecM+WCiAn8jmUTpyh4BfEvVgAaZzDlbldyYeLb5FJNZTLOQkzpMf9fj5dQDg03EmfV+
gHfNmloHaamRYUM9L9pSduWRUhifJwA7FCq76RCZ7vQIceZVIqqTl2v7fMUhZ8jUsd4CUgf5epN9
NaAfXsCqLyLOmz99cvAFcqOcS8a2lae2tmTUzlopcrhxW80eVIxCBKehU4n/g6Re895c2wGpEL+N
GlexptQxJ32TPr/i9qaSupOzpzNOyfqVqWKaGVOQxT50WjFksqF09nWxdk9a1+fBOiAYFC61VKub
Jykts2qr9qP1o1dGDVuCMyheO0RNZLcBvsoAE0IyVsSBjjp5/84EpjsFLO9jPMYR5pVEd+j3auoS
3gIzej7cvERvzZ0KpCEDHzpbDpcLoc2vAlnwOe7gH+PrLHw8/1wP6hE5XYqfR5Cf4gj1E/lCNhJO
O1411F5A1BXR4q8hG/S4eTpj6p9+r2H+Pq6ci7ZhbSRmLBjhXib+zHUT1Yf6VaVxhanrzkSVcs9X
L1uiLg8tMZo5MbGW27bU92tSUR7m69k2DHBpC/6aofP5ol/MDlNtH8G+ycbSWdMqgAv1K6e0WzgB
hchMmwsZ1zwBog/8uKia+P+WD4Uyr/j0wxe6ZdJRBaUefaYSVan1yEMfki8Te2eNfe8A/Lpj6tjE
lREdg76wT+LPwBuhNcpxSZtSOihFIagFr3DJfb7Cs9NsyMLYla6uwZdXf/6bJKRwiy8PQEW8/CmF
XY+rXntxXt4OLgug1x9ky07J+BbgHlKH3kfba1MvJx6AggZObyKvP8ygFy9Iwkd9P70hFXguxLjZ
xWjvBBOSejFmy/dtAFn3u+M8+5XMWygfeMXvMT1/4+EQoV5z2OVRKsvOk5mShtcPTfjb71JoW8wT
yNpz4CF4DU6HZ/0wyNhcjVAInIC3nG4NWrhy+rZTransPvgeyjM9AlbswMWYgP6ySDIZ/6JUnH7i
5ypJ3G/zrPdgcNxu6c5VxTN7lmrRuu+2x6HYM1eEJrIUd8t/tkQk2RPBAAh7opRcpDwOl+Q2oBF3
CiLJTVJMtowX/6mG8nDF3ofYfISvXzRYikJHPuhn5D3fyfKiJLSH/tfwH+25kaq2UqctgdXnWbkY
PpfJ034VY4J3lfLMCcuFjZW3aluWIjcWoPnH1mEaw9So9thi8zFKlQGFJai+k20+53279zkYgABN
/p4LBg3/o+latY7DVLWsAFGBYmTHU5kuMlmRf37CVN7Ntn1etHWMKRFQ7xRLxCunvarqGDN7LFev
ckXNM3Zm8xJ7n+0W+K7EEiTWWr+VM/2pTsqoTpCqjkBerODjaE0istwsMWgCAL8CLdRVWpZUneC3
MvtysVbDS0pyiH0NJJyk47PPlIqiLWzb9fOOCzkJVzr35wxRY5raBe5FGtQozrr72kKEafKvIanH
RYHpeETmCGRpLMlOTLkvMb924SZF2kaLo3tz79dYfZoA5+xI49tbzl/qulaCH2yspWkNCEiVkI8Z
MXeYgBQt8QZq/1EkjN+FjWc+VTE0liNAJIS9dMOXBzti1ZfN8xB8VE3jq3oIIttKTwJxsG7nAXa7
4ZzO8oi3FslZ0HpzIC38V8fU3bcwSaW0NiMdKmMNqLRVN7yU/FZKZqYVpYb3PLEFahDkKvdHg4zV
BtCLStyiOnNu4kMw/7Lb3iflHK/w86AdJtYDG+ZPKqpTCjM9HBn7IHt45qkbj7GBIczjiHYU7exe
nbDG3EQ0Ely9obL7Dezw0lvvifGUT9zjdg6IOxLimCYUgczBISNdMbCoOxAl4PGxFdw+H3VMbVY7
lVliRaKgjL5kHgcJaXjIoFgGZIvQfIVsNNXeZLAiOqoG2LkoJAUNWNPNGZR66QJUthlW6BWnFhUP
CNiE+EWRkDoYQaqUd+3SCWnmDOAhLO8hpfz0lr5ggim0g2tkX0cgKET5RMbr7Znkwk+10G1OoofY
Gy21fIO5lJejhX+mdEkQ5D68ausmVS/x8vxE0dEPCK8n+IdI/wLrRTqi1TRMKSC8dBis/SNMfGJT
YI8VzZIREjBO5m+4fTSIbAFOMrXNdUjf9NdvMJjpkoVJELuHoTC+IfNpzZ6Kl7UtMSytAEF9wLCl
pbuNDzHGPlEQoDVZJSRVrTn0MojLRvSnoVdA5IEiL4iQderHbMMGU1ezPB7T4qFmLYUssnd6yumk
h6TFYUhvgLlrc7Ls2Y9LJ1MhsMX7wfS1/Aeeu1p+vmPnbzQn3JCzaciXFN3RGVqG+6HMlUfePOFB
VZxdAjmMM52TXwnvTFldIssIj660SeKZoqx/rNNzYXEIzc+ploQHkxcWY5BEM9k8ako17Bfw/No0
b+MuhHtXDoCp1Ew54HKnK5LO8q2q3KfcOe1Kx/zmBROp2x88BC8S83pR+zsvcHEOLoaqNBFaK8KI
D/ZEokidU/ytQOQa7uMffvvhDBxVMN+KM7a4Iw0fOfTd8hvxFxQ2j5vS7OsWGCfK2WiN1sfvOL6K
8tMOfCMECxUS5Kc3svn7fkytjiHVfZfbQgzKxsrcFlFHGecewP9VYBQnW6ngWhwRCAUpY65GSp2x
Jhu8mZCHrKURyFLsZLtVXJ/H5bafQkES+fplzseLGf4Np+bUgRdWe8Fkj5OJPL1vJwPzJcLtBXyh
y+/J00VoYkqEoZbCmougBUvhBpNA9aTaVJM1t6rl54HglObWK8ayDDMr01kEYoOEf/AUuyFW2Sah
y+Inz8qqqH/ftktK1Wb31RRQTmm1Tsb8TjjU9PHOrFjcVSFZSsmD8+cpOhyhtDcbAd0kSOD0/1LV
+Iyg/R7fDVhice9uy9HcFa3E/cOTsNEXcApu3GPoQZ8srt6B4vpBVWM76mMqDn/s7WbQYU2cdl6S
LDxADikg+8pMF9i2TdViih7JfTP74+Ax9iS5DQ2UlOp3d0tZcYjZLWRUoIEFNVDd5gzhfCXQ8ezz
+7WrarzuSH4sBy4FcBgfNpTWo2pxEFkRaRFSPCu1kkcmxG45cYbPILz0YjJsyiRVyWGf9TLTVO3y
4PHhoOTfxRLq9kP/xFwyHrNopxmE/laQIZpo/aFbyj/txss02BtuyWAAZPUPNil2yTXs7CRUnals
OGX6beY3vSj9fj3+pWDSUQ9ruu9bNr4rM3kjsVKHF8uAC+Q3elbJnsACwhV4ALiGqFRdWrBVrvlI
ITsBDFTSiLTA9C7j0MCqk9tEcdm1VqK2RWVzl2Aws6zNoIr0qz1nwpj1R/sBqOIiwwDpJCcrJv+H
9nfHNF3l2UOswJ2Z4/cRqL174Ok2sI7K4JaSyLVSpShb+M9cLB4Sp7EdYIwWSKv2dfh9So55Iq7n
JoJ3D5MApvwZqbCdYb4m355xZW7g2tgIWVEnTz/yG0+JGxcAMTOS6su1AkfUCf+yYsfqWJgTAw7i
sgrF4AUS3bT/cJGNaTZRuiUfUX1KBAYBaW2iXNBiCAM/wECAHmKxrkbBCsu/GqQScGy0YvIh5Hhd
5AXQfNsePJSON0HqqSRsLdw0mSLTPBH6K4cuWPAcIAzFQK5bQungpuAiMrD9LnaZPrKOlaHk9qsc
tkqtSjoTHOl7avRZYYlGANhtExLxpvlYnzffClPUBRdsQebP3B0PKXegUY1Th7HbG7XAOt7oazDJ
OZVkz9r9hSzVHNtBLMnXae25gYgoEd7fEJiWsBAj4OL7qFqy2nfNpQcXihyNkQ79EL0WwjDdhvJo
usEPeEKC26tOGCQy6nnH2wfRHw4RS5D+GOg/9YohNps+QZK5+yHb+rO72iR/9Myfgk54lCdFHxAB
ijl/VlUsW7UKrucE6ZaVW1Tlvc5nwCmjsKbo0PNq3rXWg7opZTitubSut3R66ZpEf6g6TRj/Qk6b
nbC3e+vDiupPx9c4BXSLS4MBKZ9BH7HpInGUiE3EUfAD3RiFnTi8fX4UFqHryqBl0VU63bGyZ6wF
N6UBF1HI41T5EPbtaFM0+eoRJG9EDKwCsMWlZwRlOQ+IT582jAJbgOuEeJRBIYnyWOaOKjLDn7oI
svg7gRAwTMIX59XG+E0UuqcOEi1zl8uJ5e4IHcsf0CHtrcsLxo66cH7AWh5jLiq2CRGY3KFErQqo
QF7WzGlKIsBKmPIkWrDxMbYTmDF0XcgQ+FnHFn3GR47n0Fn0ou8EamlZeQ+fmHXN+qUNazbHjyYp
lqOngAOBzzvUm0WT2qQIeySQbBVuS9Ggo1RvlWucZjMpvNv0dptHiWRhdsSc079ZrpYAU1abxhD4
S889eoGMsT08fGRbSvmOuI8NiaB40EUdfWfYegOZjsMWvhV97rwwS0EmE36p+zuqdVrGAq6x9tWW
BdbNJH+wRQULgsj5SO9Pyif152X944fOGqFhqnQEee18Zh5q8iJSPfSEcrcMe4RQB4dKlc8LYpcT
q6vFXpqcrJBTJeYxNeUTeGN8wZ7Yc+ddERA31AFv6EJEorlmnSAY9J4kDVzJZ0ObNQr4FqAOexss
7FLosav6F9Ch8rEw7dVwz8W0FW9VuRu3Roa6OO3J73QTc4sKi5HklBoFgpScJsuzr5EFX6B9Y9rN
L6UeObxKZPbbs+BWPGsS/+1KW97jmuEsB0Z8Yw5K6+4qmOj3ioLd5wawxed2z5LZChFuvr48Z+jb
6OiDRH08zk+H+YUU+w0YonXOReZyF1funknOUUGCq/UEBPiQQZcXeMbnZH71yMshxN5vId7PL6Z4
F/F8K9zpV5x/3vXxhgVJtEYxEyuqKhMAuzpBBN0IlTB/UzwLbevcDzTzSxiOsIdmdkpMpZ/0Mw+G
eTVakELAVeCXqmF6vakiZx6Yb24aDSmPqqBzUmZGuki8jFcqIDIiI1JzrnUgFIorno0muyKC3u6y
eehS+1LL2QwsYlXulvKp+BwFtcrMjrOAPvHzi7gEJHeMM4BQcvFkVJreMRgODtDSWIgH3h+3EjjN
zgd11lO7pw1ZV6S922pAoFsKJdXEFWQlCYrOiKgHcSfPi3l82TdvMhjDzIHYXHY9Hkm/cm+E2Ldl
sjwzrFlo1PrRgNkUKCjyjMjrqfBeppQACqKpXXe0IwbxRUhH0QUtCoRGwj9AbeOHM0naJXNoB5Ux
J/H37o+ze+fMvmsX4IgqTRDbPOHTZE4HD3UBfUh56DmrM5v2Oa2k4Etm+KI2vi1H6pLJGoxsOd7Y
0kyJwXbHzYa/WssfezGkMO9R001ity9QSHQY5LITH+v5aVS4LNonXIE//Vc+Got5GiJ0EFGjSZbA
NMUwr+Wv5xiIYLrkHkp5tjIgXd2aEhCbU2rieFU2VIyMytZltje7e9nEkTwW1szWtwi1kqWWiQXD
DyOh+gpDCvyHHeg+QfpjA9N7iYBs3/Z+AUYGNEoza7hoU/ycxoYKX30o25AfseHbGkDRYFcllU+R
OQ9nTCU6lDwZa31weH1L3I+k2GQ3hotlmOzrfT/6BK6g32J+yuJnYfZ9fWgd8Sc1o3LJibIcbbcT
9tyDRheJPq3G6VVftioF7CEhzK6Wv9KenBxTdVFlQWXjpxQ8N/Aqe92odXvpgb7vA69fpi0YnA9m
p7Wjzyv1WJ8JP2gmL5MCkCB3klReLgMeX3b9zvaEFvBhwr8ygqnFYv4c2//woLlwKLqofpXWdtCn
F7WjwUdyOtG/64CqkhdO2mQJlNSXKk57e15RmibRA/tz6iatooEDcyr8zG1k0jMi601Q2R4dszf8
EoqfJjaYflML/UcK/FRZAM9+cVQgStrsmvirUupBCmq+OptKid9PBnlX3SpvmwR5gqazaESks2MX
tIeuLk+7mMBgoACZI/bbY4GgrbLH90SiZOg2Lfn6kPfZ6gGHJPeMv6oeG+uZ+KuBm/x/J9um2pbN
Js5VsWrzdh3f8WRMH7a2P9uWY3zoQoGQbKYUlVPO4wVJtRvLI7wlHQBT6unb7PtvpdUB7cOymxN2
929oZOgllhOx9ZOMLjaAiTgqiUZ/lvlXu2XOGtJIV82WWUC+UqEl2359CuExYKle2edMhi5YszpU
eyrz3zY2aKDF70fclcrFQqriUaAMBkCdImDaHhMA8tqIYQTlw6ms/YKfck9g7h0nZU8ZScnkGkFL
dwawt54wX+wUC1wWoPijHyCvB5CcVo8SgxWwHHh9jnc9gTlQRi5XqaCi40jS/Ve1LBE7tTnGVGFQ
qSHGSeC7oLMvKea6A9gry6Ohs5iRRvYvdlwrcjnhzS0UvzsT3wdQ+J82koqH/ZsuWUQAoTzbucHm
KHfnq+i1zCO8JnUIZxstEnD9msQbv/6jImHvufzT4x4GG2PjneLQpzGC3mdTzCR/w4+7+VhyiIiG
5piYfIlLVG+aVg/4/gAHGeWwEw5x60BlTW2jDjHNub7iISP/SCIC/xsE6ZKwXH2unYN4LDQKux7v
pYo3+8eUMaTtOWvQxe5E4MbTwBmwVfIKILMRwvsN/z0nKPmocTpQ/B1MohQRFu9P5QCej1dMLNAq
Es6fPIElSHy74fIKAIl1TtUBQBy5yDrIphUXjFEVTEPlnK4xtKius3W1ydb6brSmHMmgmhrtVpd4
KkI0Fo2V1Wv454D9ekwA83OOjjLgJM1aLnn7JmOFkDaneypzw6rGNRXvX5nXqswlKxVXqXzzYz8L
P9GyZy51WSVlgmR3ESCnH/ndMrlDDaA/Sag5eETSHUzVUvqb7/TLgnz6LsN4BUaSOPrKiiwzLFIR
Nv3RZcsQ+fjyFsAo+i5CSbKExD5tpMpOxth318lsIn5RhkphojEdvf8HBSmuIYGbw9sKr7e1Z0rI
UrqrIy+aFeQCOvFEV0GlCbneG1XcNvlARIAayWhJ+ZqDEnbhduRRAjLBLa+IIeatN2L1//6KqYjE
t8Di+B4WKLWDytrDOYXvJg9tYiQRvZHvz0TDvibPG7qdhGQE3cSPKfIYZZp+/HBLp1SZ/7RdllY4
GaCqCki/tptoPDENNtWNJXK5uLFHogKr0bix5rsW28NHaZ6JJd8+CZgFxGs/nxUYg3HlNdk2rLQk
Zi+cLNXjHKfJlY5sBZdOhHuxKUSUG6WbILqbbpdeI5nTVUnBhVf83a7dMYWkhbsOo/pRfzkcZTr7
gWMVuWocEtZytQJYLmH3C0rFaIBJMzKmVM7ZGrDeBRqllmmqDWJDRn9uH151EzSP5YrqO5zwhsEp
10C+j2ihzfDzI/Kjnzm2CExlVY2aJ7yrWQUt5ZXqLSG6+zXZfZOrnmCS+N1gs+b6na0O2YiTiRaw
P2s8TB5r3LaVOmQGBq/sd3MrSJwz6ugXxd61mRFPsnQFRICs2R/22cT6lb1o5YTAaY1VdMJ/unMf
49e1hbKHZ//Has6i8PxQjqqtodWGvSFTiEoEngdrUmYigMSVNkm/6wINVBeL7Pg6DXzmplzhyQDK
53Zeoj/8+m73rDT9tNLH93A5fJPhBseYkFFb3O4KDV+DLiCK1HNfiYCkaHztAbIJxbdbEknnP0Lp
e74SDNjSjJ6sgO7f4/DsAr7LJg1ktlswjPjFhGUy8hxWn6A0Jszcl1RKjIejUdg5Jn2I57CNPUJL
2IMCDuzYJeyMCTSLHT146gydsw7lOdlekHoxEjMrjlIncG1ukEvmSjxIVqG2Q+6jFPjuMgRYdkMo
W/6hobBfgCOaej5bWksR2kLBXxWSCPNWo4r8AKWebXFWCvqwCX4IqvlezSvBsZmYMeJaJgimvTU+
rc0MbvvjnIL5GejvUyAcbcaSBRwe8SYTuS9uYbaLdsLrJEG4BHve83G2mZ0rwQtTvITq/1oWT5Ly
Zy9MTOcEzDdUSoqeBoscvFB9cQujXdSShO5yOWsIv5GCOBtRbxtOgZ8UUPYnBr0aRfoN7L3D+a03
VQVVToAfMxiPskhoNXoQ8BgAIFbF0bYV7JeH6odh6qH7P8VTMt0F5ArX4lJETtCA5UQDYs40S+/9
0mx8kLfYL5ymL+/DUmOG4ysYvt0//aHtjt5fBf72lQQERCu2h9cabe9rYjQwo57UYegWSLmJSSQp
CqXG4fX28UojOT6Vq1Y5NPTM3oixd/pLvAkWMdu8qMIeqAI3qlibG0Z6oJpPmIpxC6zu8ZYNeSzt
rkLvcj4tOGNBNiV4OExMAm74RUFXEtWaQJUmjjYlfnZwAvCQ8A80mbEuHldsMBJONhUnsNr8WtOv
f8I9lmRY9Fso56xkKg5tqoX/yKelJ+InWP5yZFnqCZJANS7gFcKctLv1+tNEsKuJJHb4hJoBccWP
n6QLks5yf6ZbmSiKRCXhmcvqdz9g8lHOnL5PO4uEs93H4YzvvG1ZzgVUrNVdR2n4hSAIpxgwz/X0
RaX4r57ZYqsfWN+j11ABVFNX/dnVYpqJI72ANcPB9qfsrvn4JyDpLuoxkbuwAybHC8qV5zoaN34i
9P9uhCy4lZn5gwWbaCrWlybB1N/d80+HKzCcWR4XJ35w0B6PRK6Oug/Hcy7vht1tZdUNUSXwZWLq
Ml+hfzSydmGuuz4w/u76LA2TOB2sskLG9ZsvYKnYU9lQOMGzpiB1TGoSTvgb0LRimkjnqoOy3sTe
qZbVo6yI+eP5IlHnifMmj7vx4gpMuBL8NvCHTpxZgcPWP01EY7YNEOz5/Pzd7+Nu6BhuYJ1G+c3t
NTtK5kY5CxX8pJ+y2mqlrRs5YXzRNlLNN5NWohbV0C+pajIAyhkYfvKaNsQcWUBoQIi2u4zqFXDi
mrER3a/2P+Z4musmCqsy56rcydzoJUBOxwhPDE8cawm83vdyWe+fWigGd745eHcn2Oc/KgUlFwqe
mAED8Zs9cUFz9Wm2XwLU+KpLNpyqp//3izYnDPgveeRjg9ehj1gIvWktC75B6qZZhz1l1Wxz4m72
0tt2NmaRHkc5whjs1ynzAddgRBBEPc11JUS8pl/6SSiNezze36s/cd1aIS00mqyMBnO3l8c2Ty9f
Cu9ktO6xITFubACWDtMWiCPX/smBj4KgmlLHcrDQNZiCJP0Ah2RBcGqMY1IE5HpG/12SNND+f00+
ZzBflV0HPp7GvUTUF7mFiz5Y/UDmI7z5hRZbP7KRthf+Sf+5GRgC9zN94JDPNpSppWoHCCFg09/r
34iRIo5z/cPNBwomZlVyYfICXR6JtEMtcz0IIBSHxmC2FXJCw0rSFUpxpr6oy+cEhOyK6/SVXej7
akkthaHslDIxRbG/mCnLkcvpBBpUBZnBGWgWVxrJso8vudgc4fuBHpUQblisB3TR3ekE09D10M27
aY2IV5FYDF71wXqsBaSlirDr0cr0ivPf8WyHrjYCEwy2wBFpJ/GGBBp5XCNXqcSK49gQtE/d+AXU
RTMHYx+Orel8yF/KYSE0ghnkUOGEs8BGjQjWn14EzRJv6CQ7VTreIOVLMTUdHn+qIxyc67oH+K9q
52kjuvmTFfyM61fWuHFi6KKqtjIPkTQXk/KlC+uefYM6gamHoVq/pI2j+Str9aF5Wbhg2OsVoDCZ
qdaRS28ghNbr75dYVvuvT74HiawmCgscbuybpfTTyJp2R50g+bsIgbUyqt7ZHkAWz/DeDTfP9jG/
wEI8Wta1oTk7BZdKIFQ7u+/KMwnxf3MDsolZbYSgfRdCIq4SjOpBtwo3JgOThgoiputrvZWM93HS
avWDmIutYZUGgpd24rJB3ZzE4nc595wO63ynmx39GSfUhfLQMyRSBX1VmTpIlXxzV8dONhWoC3ZX
6YfKgys3Rbp7+m2MT8QqM6ivhxjBik7T0NlyuudHEvpAGCdZRgo1QPaJN1su3R2L2fQOKK2QdPw9
w1S1IlQpoUOQUHfE9fk9kAva2QlaZl3Q/94GQ7Wjaz2gOMP2LiWW86LFyHDD6AOk/3tWxCPI64So
xJDNvk45L9jFPsEeW5ffXoOsZQ9jBR3cMsicRGKeFBjgYAP2VK8sKpLDNgnC1FYsnBbAJDN1A/K2
L5tBcPjz2dl8mvUivaAFxg2CJerIRZya6rnlaCcK0QPe5HPrY6NqB1LKT9Ddrf8zUGtzCmfPI3d9
1M0zbKkW0XspRb/RK4QLVJHkTo70r6uK86u+9UeVO+2ogwS4vN2qnxfZkb3QXaoZPOrnCrSlsy+6
KbwnyHCJMqQQGOQpZ7XLDnPHkekBASUGBK6ISbZKLQ12PiNrQ7YFiLp/+Fof+aqUBXgEZfiO6cL+
bUkoKtx8p004E4JIGjXrThnbQhohmaH8ZNWDoscuk+CvKpiaFhm6OMZfqq6tog5B24on5IO3m5kZ
B0IQNezy5YuzNGfrmle97SnNTWrbqx/6q3qSJKmSd6K6gLaNikqlMuCJdDe/Vulp4G/6ygHTrJvU
jYqsDqJLP5LnW5EE1dRSmGwrsjORFiVhmAKncMpVRs4tJaswUE/KEohyRLJwXzM5gWoIzeKVA3Oj
soCOwJ3e+KLkyfQqQO+jlqmtqCs6UZ+mcdo3fZEV3ENXNYzVNcxR+ZXIBjCf4uGQo+J7GptQNniB
oS5Y/MIBLB1my63hkTpZn5+AtmnS2dhrGg4sKX+j9+776rZDzeHXuwu9+ub0Ws1NeI92eXjsyiWO
sEUxrUd8OB3fNa+87kfoN2hs1ddLm96gjYWIadgDUF+8/bSH8b3sY7mKaB2A+Zzghqv+wokqBZ4p
52+5D4sYKqFrClrR8MTawwnytrclN5ESh+CxU0lTdk3PEVMWtyYjf29kGzNAN2ZRp8v41ELdF4TW
vOKsEpL6oOVfvHkZiQJm/lbTCu0Wwrua5NWH6qNvsOLJ2a5BxtsFVoKMze0ddCk5r7QlVzI68lWQ
IW+jaaPuUHBqraQ6/c8TCiu37Cgz9B+ZUMjFQPB1Q8l9WZffFenrB7V5lvaJA9efbLRXo/BrhCFS
dq2xtCJ8+BxZYpn1fQXC5NQsXcrn/tZLG2ZGOB1mii6efzwCvc+IgDq13x6AdHE0KgSNggHpo9yN
H3tLwYcFbR1WjaXn5T3NVjPJGFr6y5+n/78/5QRUZn2o4jjxnw/4DJfYAX3hTw1EP+5zmY0tTBFc
7cC+ajGgSu1acFvbapEU1jjmY3htcqkAG7/s9Ep7+S714U+oCQIqrcjtoO48FoWP5cBEWdX9OIjw
+PJ+owV+AhqBJMiEBynyiHwgk/QpRc6petSfeL2fXbiIQmfyM6HmkQtSqFXlvIWQKO7xvnogsNvO
sKVxvt0lC3XaptdponrpFWA73QJhuEUD7JRsvWLI0x/ukSt4cQPoohJiVaIoJnm5WJYienlfVziX
/83rdY+bcOLGUUpftE5Kv0n/foFJ3iHaBZGIWEZPdXzfAkxhoruVm1Ebr3lH41QNOf5Xte6cvVrb
CBsUI6QnzOC/iDKT5qQEiuZUlI6KbqXnltPLB14whdEjLDX48J0tanpW3KRhioQuj+V1WFzrSNtW
fg8VTrtmCMBRUjhlQTz2+rYWGRtT4s7b/DS1hEj08ddVRRlFmNd+vk5vjbeNQFBpeI7uJxbeunhk
Rm+NaR2cvPe5sMKdMqdPeKVVK4PVrmCyZKQ/9LiX06RyqFGBwuONT+hCyGMPF+V7AlFE8w1TdtFP
oID9L3WOYxBMWw8sLNz5nYCevrYPLRUDabPed2WhYXg0zi+IVX7MKiNOhD4H/wbL1DRlUgacES5d
5ikubkKgLcekc/px5EJJE9FYaV+00TkbRaYWXgWX0bBCRrWx7S7+yaW+ZRzpc731LdCsfsABJJ/5
sfZ/LsacmdOacsHKI2XCyLP8WaZc6ZqqpGDAVTAebnFGHKBFjgKhIN2Je0IJGSA6nLpa7oRLOKF/
nJw2JcxiVTReJMLznt/Y/SXmfMz20FGxi4psKmucCcCvtpX8QfC+pJB4QO9lgOPhdRpzfyTo4wTd
zTj8Sl9gX5oxMJx5OSkQgP7xDEOzZiHbI5nqTAMTBTQILPTW0mgg1sAloxN4aTigwVlmKZsHtDpL
FJMOGg7sIOwtx/RWO8n3m+S0LNDAjwUwMq0+P3nkylvqoJQeKJIyWEHf6yjJ5DjpIiHXEgpEoH8x
ry05k7lTJJ7RYC3ULZ1iusRFiD1wGMfKNYb7i8wSBzjFPGA96+jW3t8OHz+mc+3MIJEp230NTVO5
bw3zQczNee3nhhMtSC5izxy8b9urAFSWntrBtMpzndXawMZyJb89XHF2cWTLE15mCDZZ5gPxWLAj
mYrlA33RiNuplQJduK3xWykawPBuJL8wWt+r/KluPQ+KwFfbDzLh5VLxlOZPchTqFU27wM/MSkTP
jX7viTfKFjMV89pOVAe/SaZQFOEdEHuvrIKWkLU4sUqb35nxi76JuLDS4nr/TFi7alOKg9vXDUe8
nt4Yx5k9s6Zhk9OA3wjvJTozKT5QrPDYJPjx9GYdVdCIU78nIoBV1bj6FWPsvEWD7EzoyFHwBP1h
Hj0431pGnNTooX978S2/+3BQN7J4yE7boWgM2mV6GHvJtZHfbD/KzUxbX4L3hZgrzG9PkmNIiVuf
rh0n4p3GkVap9vevyFsHeT854bammCrrjJV4tXDyIL78qOXYkxSml8EtTqn3YVMEFaU93JaHLGk8
Zm5DUjYjTL+qObwff9nhgrZOS7bSHe992VbiWTg3PBQwu5dOhFsXUfFyLVN5/iYVN88mz1Ytps2r
ztlNhC8HWSFgPMWoUdn1simq3AikwmRcNRrO2iBGYV3AN7s+sjm/Vs920nBY197bmR5xELEfRQqa
Xahn2PlW667cu7HLNNEBy/5US3Xmo3f9PahD+zFJF8Royb/1IZtTvPdVMCQE1e1K5P67kPEnrn4I
SR22kNWciVcjyprRyd91ptiV2itov7m51yzBhHayosXm+QFmoWFqriVnXhhevSZga95Rt+aY/Oxs
j1I0VuYGniPFFoOKQZSrDpO2mWIp68MtnRNVng9ryU7U31mAzqxHkg3R4a1jsChyE6LkkFqFySOI
7F3542QkNQLXQ0IyNUxQA0ZOmHQ7klS7hBDjs/HYxVzUkrssyrTMnT2sPRscwm+HQz6nsOKXoHMD
/hK2xeaF/2Q95Oynwc8qQMl+aD7Nu23xrAx+KR0HT2tqiITuuAneN9t53meDb5sq2Iuzh7r9WQpw
2+ghYwn8033aaYHS3cl73mMXPUbokxxsEE1pRlx0lsZ1b/E2iHWa4oXC0J1lyF8Kos0tMgJMczwW
kRbqamNr9wbYkHl70l+/gsaVla/J26EruGcgJuN+NgFyIDoED8XsES20ZenoGYfeeQh+67ST8o/i
NiKD94AK14A+YA+H89THldgqY3+27yoM5jyFjmAyxWgOFlPkGzlaQa4y1jkoCmred3U+XE131rb8
c/ihrkzWwOI7RPfVCHa028k8hjo/vmQshMc6C/li7XLkChlIKE11+uS0K6r6tU823gNgSwZE2csn
0+E8g86U+abgmBXqQhVRJYKguuqWRG9ZAFCbxdH4B0fqLeBWnChUFM69JPUG5t9M3IYHyjf+ISEl
Zt7h1RISd+X4vmxpFDO3/SiQmcXbnYh/KlF8NDi5uinuNZOswJsJ6HvWRaluH0RY1Z+r8ZhYP0sd
kk6WtKKmlR3xA7uxFZRM70P2BCV9sQh9zHUEqdhUOKPclYBPZbWIp3kjv002IiRz80ZPTq4bZtfp
Qmbbz2guSDo3TQu2SIKKpr4cm5bia4EseyluElV2GJZzMMTrzrQkHohEpTQeBuFAX2IBIYH66t15
aEmBKFi3WxD4xIImbNBII82OjQY/cY3MUirEC78hs4FXjFHAnTT2M2nZ+IfyVTdxntzJ6mDDNmLT
QFtFk6IYMdTLxy7A0wbFP5nzU17UwWA6Ct6k4cZ5okJ1dWoPFKAi1LqHHlPS2N4kY3Hp5aO4HDcL
mcUjV3nmlSwCMdZb2sEi/MTqSeAi44TmKzPBq2I1MyOALhxkZi82SKU6IqEbS519qQUbdA01PViZ
WyowRw3CSVJl914UKe3vM6+uzVkaqpfEzcd/gyuVaCgXpsnyyLtyAMg/6nJHsf1zjW2ETN95F/Nf
f9ogQnXNzvVdCdoE4l4wtc/l3p796yuJxdnZiE9k0GsH+PNYTnt0Mhp9CvNEDW55TIw/h/QwBElV
TsD8IUr4MwZFvECuro6uas0Cz+7mY3RfX7i2YHr1tF6SLsuxxnnUlRxY3rrAHhK2exclkNGTtalS
jZhz1fg4UxWFKKqShFN7bpWeUWxwzOcLX5m+OoIfYj21F5YNMOMwYaENyW/Su93R3gRcIXLqclin
Pkx/K+dNlhIhWcsZlaZXrVdrxRb6rSq2uEmvCQw7PcKa4jJuCWzf9jCYnMb6DbFn3AlvnpBQks6d
gvN8e4sDHtC6/dobfwecYSh72ewfWcMST6Zn3y2/iTCZZssP0ktHXUaQQzaoC/wv0xl0ncRcaeAS
0Xm3cAMyJ72u9IvAYb/BkXfSI+dVVDUYpkOkpangYqRJLGF2L5+Gf+fRck7dw5HnIH0ouCeEZBmt
swnUQoA3DnhqZWiXTxMn4rX5Qkw62Jee7jtAtIa8WOmlbpUJ1E7lm85bN85XIjITASNCF480cEXL
X4l6HumrB7S9DeCj6ZIFa+HMxje4L4ks0vOuZqBUFqgZxYX4HvFcpMv4m2kkRu3CYCehuOxxgzw2
hc/pePU2MklasVLIPAleesTv+F6lsNOwr9i0eGaaoG3DLU6nVhw1v4Q4+ioe+6FqoS2c9goDEUjL
kBj2Qx5wL1jpQr+83rbw9WR+hV7gAIXmLi8NzK7/uwdoO588uCwisiybfud6Ix7wKuPuBjaNH/5N
llQPHPI1oCEUwZaMy/Qo5s701b0b1Q4Qktzb8TD2C4vqlYe61vqqWae6UivSK7+sV/x62I1L/q9G
94Yb3bLSw0tK11IAtt8VYcm5VDHas24xQNxXJ21Mzs151cUHcney2nsy/dgv2HTUtvQNNY/DhWJw
nxycmw3hVcRvGM8ImX4peM+DD4UAOqq90qQn+/P10CUrYczqY3Cl4JkT00FhsKKeFIxqIq6+O/CJ
tkAybAfuUQxscUMEIyYlNkXvP8g7gUZQm90GGtM0BwOUZT3IzfUMoDZ1XQdXykVTimHPo2ZNuzvp
JoIlLTcxjyHfySenHS7HFgelM//LwWtzSYaEceFP9WavQUZiOpLij6UlwvdP0PWA0xU5idH4oBKw
MdlXUoxsYt7JcwoTfJupmscIMEhQtWbMeAIoA/Pqwb/g85oW24DMT2+4jw8G0nRC19+L1uhsBUDO
bLgWMt7YOBm7B73IgeSfOQW5ZVwKxgA6lqzwZm7r4umIJN7sRPli+uNMNWwxwooggWf2bftL0eQZ
fG5y3SkOmb11kKWO1GKo72yfRI/0oa+jNwiRPPbaJjZb3x7FchZZPLISP1W1L8BVE5KMxj1Tldk7
05ScPdICWr+hZk1La0Wqu6tOVJD3Csa2fXLACCElFpzSXs7r4dAentFlYpPCDdeIuyPkrNaDIpUl
L5P/F187ri4Cw+Y+grtICaJwYyZmnJbTbv8gP0g5KYRbGC1l4HcPkc7I8oViOl5GHkTWhuzRWbgX
9U2B9ctYxteiNQQS5c6EG7UPZW2kJROqvCjkUHPUXaft3Q3VW39NMzpQ3o7VWpJRyaGIlQqoyP6W
Oq1GHf73GyRj6QG8RVHxowH8IJ+wymbsUKBvJYhJr0Erigc8rhGx2xTt5tm3Yuw0iqBvpb8cg/ZT
/PkieRY7ImF37TGsgMisH4ebm/U66kQzjc0mrHITe+LlFSHRi26vYLAW6/IDU9lG+BhVp6FFAytB
vPUp7fElxd30QEE4LNFqI8SVoyMkHXt0o44w7yyG3340OK/xx+kb3fDAh+L8m1Tbs6erBk/05FWw
8ZkOvUqPZKETbdU7NyEd3Tcx/mnTBl98WBUZFNaMdn2p4hjr6SOXlPwXbZfIsgkk1Ia1K6A4xKpt
5cfzN++ACkEe+hzt/WKUYElcMHnaf/Pgtkd4NHau5JthCHMoma9VjoTEq7SayHLZWsKbGZ44MTr/
ZSlJh6JSUYSqkQDxu9pgLtCp/uJPk5eb+sH0dcK80HKPMNW5t4VzD+2PojAls2uo5pmaL0bnbd+v
nqjuC5wIgFvNE/TZxkQ5FmA2jx9i1xkmpI8XEjqcvRJPx0ValdjFceIWsonHyTsvPvxKVNrk/V9D
plzyYT9hW0+SdVk4EMysK/7OVrrs6YMdUBGxF6FIQKqXD7mWJV5Yn+GNVRxCmR7MryG+NTZ6K0e9
Gh5n6KybhB5htbn+kL/8rRKfUWJZOzuPucdo/ywTC6JHQ4y2yw5djz0awx6QNYvH0iJeDtuzI9My
oUV5tBU1vgZtwR7xUziuIvvAGW43+mWreHAGd1gp0G2g6089DTB4RkiEYYR88p42/XGKP7LBe/bs
5ueYE3pV+ds/D89WoREHZMx7FaxS25IbTV1pPMApCLWTou1Jbae4z6pd8bHsqCiTC5f69fvQ1+Ic
G6/2w1cvwj0XKCkVOTVL+RfbKQpME3YI4okWmXB+BUMkweaxEb+pKWxIDMPE/VGOA4Y43g71l0ka
7rJXwYVUL0XUH+jqVKAaGLJY+Vs3TWAjQkr6KnSY/3ocRSk0SjqQO1OoijNfRVEAh0t0874H7e15
3tVxjcX8YbID2bgfUPPD98b4jNQEX+KjtqG1svgBfFnLWx947DiFpI1OT2bCbyIrXLTpmHuAkycd
E+45vMiMapGrOwxEdvJKM43Cyp/Bj+mOz8TjgttJwBiQWGriMfHyk7Ou5XfHPETG8GKuUzXAwgFx
VJCVZ7NWkLFQ1/CPGq9lGq7oBiv4VQ1eNphLq2S1YN/PryGv3D/NfvYMNmUWOMpZz9DTmz+qK2+f
LcCCh9JgEDkG0B9ExRtU/0bZcrf2W9RvzP8/2my1QTVQH7RQmY/1YiqXHWpBh5T5r6pvm9PyLIBi
aCCZHrCVtnfjKKrad/Gxu3E4BFYUOhb+FzRn23czWG+pE8mbEpTYu0Tp55/xtEBQnfiQKjQbVskA
FxIi1awonEV2xbXj88PQ2vopyscbzlxoDIoLfieBQspv7vyw7I4FtoOszHOHVZwi0ILuFsYkKF2T
K4o5Yo7H/pdOybFmgKtGeDV9u69LHCwG00XDWS1ZJOTUKAyu6CsqdSEA87eJmCvWCABNl4xb1MCT
iSUeTaUAR7WH4kBY4kMgXOGjB8T8BAHTDhNfxDkZPRghOANfLnzeXKnOrYFhRnYlAGKUEoS1ry7h
2XrORK+KqbLBWjwdm7DM7Kc0WcHDMbZJkCUB4zgyKbvEHYnBAxc9no0/8rGCvCTt9yD7BfQuxeQh
bnB5qoyHQs7hYcpZhOn/llYGdnzkuy8Th1JoMYi95fyRU8kO7t4Yj9QNG8RBzqXwszY1t/f9/KbP
7Ke18y5ndI29FvBjxvPaoyK3Tl2WS3IE1ekPI0AiKPoWU3vQdu5l56gMYzZg6kVdx02KQDyQBS5/
wWLDoyX6xWbRVM2meTlRW/uWjiuHmAe6SdelQXdnA6zOkZHuyzw2kmxs6r671gNCIsxdJJWPpq9U
1v76+HLyEJ6fSm2kjuUAfSmr8vbl5EGuSFePAqvKEIUefJMqRBptD+8iQwtZpm41ngWsTlMQ76R1
NxLOKjV6/jHCyozUk21smMmYA/bNF7Yx1f3I9ec5ZFzsb94AaUoScPB3+nH8WBnHWscnU+p0duur
RHXiR2+9On7Go2Y9zZFEFNVhwL9TtoDliovTxOGtVJKEdgS9HRz+CFD0Z5DYII1CdtcHjX/qv7w9
RJwNJD/y49q/sIGgr+07vR05of1O3dQNOHUfC2y8eWK3HserP3erBXNd9ik+zGOdk9X2N51mceiD
w/HD1CvMN399Rh7toMRwW/HpiLqv2MqKJ06M2gaDp6O1hJt5Y1KV3+/PNLWswbE/yTiWEtebpOSn
6lPV2oLt1L+ygnL0A+QFdhlYf32JjNCVAILL+NE1MWq/VXBZqxcNzHQ5pcIUL9jsNEINFxkMKADn
LHWXvFTIjB/zVoLqhaivwE90gB9ISoFd1emi8Wy5eN2+mDyo6KDAnwgmtbK4xq93rouNywilDSOS
UXfjjSh5jJPVf6iD2VXfvPdjccoyNa2g0IddfwprImi/o48bvBh4yzdo0i5rCq0X9WQHUs9DrnD8
iYHgqWvWLxMyU+maoCdYT+Dp/iF3BhZUfPjeXO1/i9oedTmPosFxnX4wcYC9XmeHEwC6STqJ065S
TXAbN1tf0c+WzxSK09R8IDHkah8gVGc2DUFLU4VLYWGR+xLSmDejOoYlmz74fkj3NyHQVJWed3ui
54YBBxr56rfr9P3/YZedBrd4tO5DuoKHwtU3++zqkMgZQ2c6YTNrEOhVejaOZS+727DUFpyjK8NI
rfPd5V/uzhIIG/L8qU+rnjfVZGNhEENuhUENzZjvoI8zX11Nmw4iOJVT57COW3s2IdK7QQqQQpTI
XR0Jv3A43U95tV9/idaT+3PjkUE4AJUnBpkaKJfFhJivoq2CbePby7wESliYvI93g3gFqraIFGdP
I/iiCC/Gv8xMFRJX44gFsTO2e8uGqEiYIwgxNbvKy8YcMwQ2ZNFc6oQVQtJd8z2oWo3wWQRmorY2
3QeoR951mXzT7hI/IFipAiOTqvuM+26X+RLBQ4MOF1sm1RuZqhF3yN71gNY1NFaPFykvCTAkSSsV
M2iv3oiy7ErIwFpM1LQdF0peHLohjr1PDhlqLC/zIDlN0LfoJ58Ig8GJskRM9AuVUJL1jT06i2ln
vskXkXlOP5Al9JD1Ys87bW/YIYq6dLduc4kK//aAPSQmVxGWA0eFbGWE2u1tmPoA0ynXfDAe+lQ5
+cldu8HFg84FP/TW1in0JVCK4EndmFRWjKF84wfXKK2vHILvpoN9F+2EuCxTkG/KWmFsZ51Kt8L3
bqPW8SaduENaqsKQvrqb0GW7pj0JMLzSgGCHbWIMhS61HM9LpIbIA3B0qe7jHDFka/FeasyQDP8Q
fGX6toaF6cEK/rfWoANARIEmfDo42Rqn3PZAOYSJpa9g9FcL9XF/w04CrsRIUkiP88BV4gMHPlKr
HwK6iCyRq50IIZPDQ7ErW2RjzudDAX3HDWHuNxUD9lBjCabWyxQCFWk2cpJklqF//JJeUA1WYYYI
WZkCzMDQR/NHoqkZ+dhjGDnRn+YTd0B5z4ep/e1e5e6EpHh4cRHqyLDjPSrorkakBwMyoHgLW0n9
JIXXCV7pjYPkv6t/2QyxtrLRGfl0o4cJfUeFrZkCVL+S8gmv1jIFOhXB5wbwgkzPbhbWI6kGFdCf
k1INmAdcvmGFL1A3sy10Qi/08Ezn5TtbeiToQyC9LTSXLI9MJwbdey0aVB6YhJfYcS1WHTBH2UzD
IQQTwlKygM29nfqAXpPwM6VRB2aM84tXa49L2KS72Z2cje3HFGMvf6yp/o//uI4v34YwWtvHiUro
/eMQCjuSHPfjqwdG3vRoVPCx+omIWfFMdvt4uUMgvArTnMtG64aM+E8opKuhNnrL4UvT9F6O3JAr
FNc/ywKJw6zK0QfsjWuE74ZEPXe9FDzpLYl26BgrfZXS/rNHSnEESEmR9WvwnFgBwBZB33KFz3Ks
O+2fOZylRQ8pWnhvaTWozddt6nPVlpnRcCWZWWQwVMmvvNdtXtpGblzG90c61VT2l+ECPvP90dwA
OIP82kYJ2b2Uhw1qbZbVhaeTENyPEy1SuYbTOAcFhTId7PGiy/UmpmrAYrcexFJ17XhkeQvi4pBK
I/CYjolzD+jrcUiDQa8JlfcEO52mIQEmTZRPTj3t9qgmeQmSYHDWLu8yCK35c0fsg6MABeAiNz/o
5U0LQK+gziYmshbKFo2dyhoeauFYCczAZhjCxnlpbmqTicd2Sb0pwf48YI1ztKtMXAVMg0HBWAG8
WMxGmsj4KETiD7SQMOIAN1gE+6Rwk5Mhfzmxp4sdiek1MIH0d8AsKg+9q6EKz+lr8Gk6OYSl5CvM
wconSJYN73Roy+MD9dO3mCZh5hDvVrMXoB9YjEmv7VI0HGGN0UAEljGXDgQ0jLw3YSmjkKsxMziU
4HSKRwegBrh3DeLiRsu6k2PIQo11xTOW7MFDtUFafZ0Qvqs/58ofHia4ZxJdkQoDLAZA5fsXDaKa
0G8//KSf6aeUdnUE5dZBpv7GY3UXVxhrhEskRJv23Ez7NDwyIasq2U6bQb3L+lsgDDdV1hgou1Yo
UmtrZ2374NSkGGDeloPYYztw7pU4dKQ2Rw+/if0HfHSPseRX9omFJ8Zo73rTnmYflWnhNSd3TcZB
4rt3ZFrfkgqBTRX5oYeKMBI6vNHCHq4aumwDOxkbdN77U+I0JQjHPqioh2VSicBjtORIS/K3EWlQ
RGEHkG4sYB8Q8ruVDqSjbDznY0Wn4tWy6dIOcHFY/3wV8hPVVDa8W7SzOgr2uLL923XYkP4V1WOa
FBPj0VLPWBaXLRlTrcN3RAxMXG5abwq7DtE3/RMXJPxOugVqBrjV48EUvMvtEIWtGG/FCEdFd3/r
hltHAllpuKZo7Hfr0w2uPX5Gw49BKULbwKqp+o/W/XBcakf/XTbt2mA2kAs+KnygV0Cg9jDHSWjd
CKUUKaJz6+BI6qU/Je22vFg4i0lSp3K99DJ2vsifR776L9Q/sHjQuKhFDKJviaKi7nHezNftec+/
pGiVjqDtZC+aBq+2/4phoKbe2zS7OZ68Vsv9325Mel9BqOBjXdqwk43vog2baONaM48AxE3uPQXA
sjS5EheswjTz5MC6HqYr7ljCJfnq+a5rtM7bBqanA4D8ThcrWkHw4ax9DT+EIxSHGHp9wuPVf/wD
f6T3fEPLP+Y4K7Go7uXq1S5H7P24Z99RHV2LEUVYm6B0R3/701MBGM82qd+55cR8ZHa+anbvb1Hb
ev7tUIMO5SDbCdtSkEWkIC7+6BFzqGKE16sAkQwhAEBcv/IEuJVbl63DBT7JvHjlixBgVzh+ez9K
xXbxYTvorQCh5EiHNq08bl/d0CzYo3mvdQqtZRDtCjz/J4T3YJs3qO6NIOaHZZBZTKklRxFhhAZi
KBttRIFP4zoi5UjukYQ2XGGJI1nv0/e+OIbhGLde2m2ekUjRWTop78OM1iKduclh+Nu99CSc/Mdg
7n57yMyonLlGrblsmrClkfnVo3aM3R2Qqb/mAR4qg+WGp7188V5oAnHFtY7b7Ca45cQSY7qj7PNs
luHasOSYDkZLh+llysasfLog/861blljZFacPQUnHup7nZfbEc3Lblfj8yLusdzaciRBPV+q7igj
QJGoh02ePKyZveJQ6Ok7vvT/CpD/bpsxpEUlF9y+SiqiCWBMVTlUfLAg2CgAv8uACWwb9Se6iF67
BUbjT4oYtGaSS7yM4FMhbkGnwQJv1PJZYQ/GVra9Bnn23ahRjkig8m62zQGz4Xv5XxJnXjrmyiuQ
LrOmsyPFJJ/e+J/ESff1TMTUbMwwcuxfzL5SCRTvMtGFEHXIYhg0RUU2/ZH9I4RfNInCe77dF1Bq
Lww+QNxR//TOM8Tn7gGCgROg4H0Zx+mL2tF+NnMoLHzQYeXrr7D8kgACR+gFTLaVSaCZ4GqRZRaL
I9CDksIA377p0cQtgSW2vgVnZZzKT3YHR6qrY4+A70SeBBTt1D2BGk3mdzKIa/5Ogb7Cr59vvpmY
P9lSihRofJzxm2Amsmt3r3aZBUESzxsNublfObaCfNhcQh/+hA0zx0Cs8/ZJQ4Tl0aE48iIPvaiu
fHgsip/S81bkYGufa9vE5Q1oKGyZXp7xrEZQ8EiAepH+QDKax2toG5JYhIEYJvs6rBqVTvUNOgyz
MrC5uqQOp0dthe4tuujptN6HSVw5+B0quBXvroP8YH+qv5Wr0fJwYDGkSdaFMCcv4+uepR+Rspz8
Ve5GVUzONW2h0mA8GO2PArjJIfcJAqt/dLYhe1A+xk/9r9g89Hpg/yqoZmwCpdXOnRTL8+dNt/6f
+u5JHwL0nOqm/7ZXvXCHpNYq5bKMVV4YrJpWGYh4K5sVX2TrkY28AnF3lG0IjVxnGK8Hb3vL62zT
pSUBeQzvxiuysMJFYI+73DhyyaHexFPYs7qhDfLjVjapBC/AbIPq5mjWs0S7WtSbLJ0F4nonZMUq
r23EeP5vrgnAmHMtLtfuCFtuY7bREcVwyKolQnaXU5FTLSDe+iSPbmCfcxTtywIAzJr15c/oVfYc
WZd4+gq84LOgzPoPO8g+6/Sj9SrKV5rQBVuR9M1MA+lvjtW68FVV2Rtypog3r6zM0yXO0A21f9OH
eEQvI7AUvv7yji33UpU/5zqwviaz/Fhfdya749m3QT68I4e1JcYQWhv6H/XWwfGxf5vtJduQNSxL
YBKK9JSwwjLGQGR8B35Pq1kN6v96TE1HuimbPzvaYc97sbzlqEOVGdR7qDiOhfbBJvOt7oiq4zU0
JaE32IRsFTbKKQcKzZfMLWGtOdg8QQ6jKhW7XUOrbvbAfL/BjB366jxSJ3kaeDU/Q/8KNDdjvK1q
Stqhs8tsmJHYAzSlmJQkrMw+VERpqh7NzC/y5Pg4sJSP4+mVLPQjDVgWMzpAeJ4sO64E9dr1vQ3U
tJ1row0dFWjS+WmRFony1qtlz9QmwCX67knsl6HcScoC9OmBs+nglN7u6Any41kAzV5j5kPRh8i1
gGC7gwirDRAzLXl6jMLmcN8hhO6pLqm90O1l44QoTSJfeGzfipfS1VyWqeUC6eFQKlAm5MFtZZsi
lbi7NMnI4tWNEiRbGn/SEWsidsOzivp5wowizZbeouAvFwcOPg1zw2D+Vu10e4FWoisJZinExfIr
39prQGUaj1PESSZmrhnKfNZdqdX0QQCoxjB6PgXxSH7fSwJHeUJwXAvbcVemOsr2n2Ik9kNadklx
zSPRWFSUdhehq3IwGJdZ3x4TrnFF0Sifbb5zOEleDd/NgDXFVuP31vNxhUu9BaTVeocvdDMD70da
RxXNDr4kiI5RFsrCGMENKCJsygimQ55HrKw8NntdSMP1fotXViynSGlZgsVr4KGtYW9gU3ZEvZw1
HBTkb3RLJeMRNE7UQE+Eo5JNi3cMoos1eZ7Cgz1a6Curgqg/xbDyOtmnFJ0auRDrskT12LKpO2aC
qceq8B4KTK1byV3xO47L1KPKI1Db26jaTp07BIulE94U1KUs6cduf96g8SHKP8WUi3fBn5RMs9CN
sa6M0GIuR+T51gE11nGCPG5GtU0XMpDVqa2bliYw+vYi8TVjMC35IgzSeQNhwV5nyR1AnlsCRbJC
t3Gne5BXuDIOrHNRiiSuM0LsQiZdWNfkCcD/HNavjVpqmiFz2kh+PQ4dQfX4aw9SSGlw19MYOIkV
xmNNZBBpxwRg8HYazASUG7nw3Moco8pJIz77oD4N4JfkfcvBjLz7rRdxyMFUt1wlMoQT9sdolyDU
gfBmpLWYbsle5NgSDvbB0I8Fi7nt8PrCOAM/6ftbKD3RHtfSF6lx41vjdGU+tRy5NKEeE65NXxiG
LGnnOna5QbGw0uCr+wm+DrDlXqoe574vrU9HoPNk5S6/UFa/iFvBy6J4i1Zup1RLzg7TRN9JxnaI
RlsU1AAbfg8OP8ggLaqaYn48LQOIyak4LRJtNnrvoZ52zp4Pklpb0wWeFpTZghDoyHLWg3f3DUOd
FCYkRVHSJXomKYzDRjVyNIvpGPbbNafpbyccRfUgCD73VYAolSNcrZDc0fml0SfvmeSXEomXbJYf
7yh+DOzOO0x9m1K75xDCC9vaaoAytBhqYUyFJCfP2gy7dCWXEXhJWpHDpffJ8lBiE6yxZoF4Wv70
3UZNXN9eY0m7B8ilYmmdHsBU4bu5fAuuBJBlAgAocF3gINX+rsdmOjNo6kb1iSVQsaraU8RrQYh7
4lC6vlM+v7hS1gqTkUoDtnsyPLMYGjcfnftUWCMsc50c9h9mgm1WLp7vcd75Jrl3JQqrhOWfoW5X
oCObylsAwhXhnqugTUJlJggIUextRhVvvFsnHTFCATWveBago6Bw4XcpbIn5xPBk5bMXJpbXGbRM
mgq3Dg0t39I9KQuwEmbRi5IQHqlhL7pDWQBpiyEFANu59Sd0hB1HfDOFSJj9g+wFUO1K9DAnz/dl
r31urs5n0pfczQTgjhDeWfwB3JGY3f4uyLumULl1xg7xr/HaMgXhEWaAXVe5VE9ARj1Ycp/+J9Is
WawxTMsrK/kET6KXU/HF/7YcZr83/pmiaDbjLK/f5rLw98xGNY46SfaBTXQQX4W2siC24+koir0O
hK/rtLiaDkQ06H5bABaN7dYTxbxchAjD1098g17t9oVy6GpR7DAAZhFXHVJDCijCEcc4yKDICU3q
QWlYHlTYjDH7DpsKlERxeWlVxq8NkayyPzUXZnMbUEEd3yyrDIivcxLtcZVxTMwcYJwUC1IxAC/x
+6ix/SmqJy8LkXJVG9fNX6s5ZiznYt3JsnebPr5Zcs7kVX3B/Uy5/g0ltQ8PBUW/rW3LBD5hvbKa
NId8F5ITmYQBieLw4lzXI7gijU2UYv1+7/JbdgrZNhGygFdi123+FSS2XEt4VG1vBTxN71MAyGLg
YnsksqIAHGMhLNJ+8GReRbrsq0atvLW056hNjHkt+EYlkDWUe/Z+jFY+mm9bLwO1XnpDS++nkRLS
mOvrAuB6g49VNZHaAMOKZ/MMxiHnhQzL6bTTIVokKuChQ1C8cTkCM9k/6MUHmL5pwBIOH53pyCEv
Shb/yaikxJoHEjv0qxYHVGa/tqnOKpebsMbwkEor96FRihejVTgdjxmFLFI3bZI2L96c1nfgCra+
YJRt8nW9kin1WlH+ArGe2a19yoSTv8EgEa0MJH7m5MB4R1qMXRJW5FT19mRy1kAnYReZWm1qWfgz
RhFMTZznb7zZN6Q1ajDyn+KuDQiOQpVe92tDCrHKvQTIsTfBeutnBlMJqGae5O+CwXxg8QSXPJrr
z2kf+VbaXEk5SCC59FwytHY4F8OwULCYmHWUgN81TxgZf5kaAcMswNiGAw30e25mM1BW+OPC1G/r
iMPHUWm1+9ljlWuQruOMWW88ClfzpkJ3u0KwiLCarWJoUuww/EeDU30ZyiQ19xSzQOIInf9jgtU8
l77XPEqXsdv/9l81ADNZY80t1irWTKxDrNs6wtxfrJhMDUNmcv60MbnwdWmE7aKEyRSl0mGhABW3
6wQ20NYDFFGAA4HIiYThRpUvgf8ZgLUWpJDmCcxm1IxHHMafuhWnQeYsNKlYCxgeVN7dVuYuBSjh
3B28Y2Sxc9nlv00I8zmmNFkA2MHH6+jj0c8EXs1sNJ2Mtn2jVJAFn9WKEYtSD8sU3xAHaOMgUt9o
fBhUF87qQpTE8ESQm9l9jDUxCEX3LLSFDhIuYzRPGN+M7F0xTv7LoJ9PIZc6+0F4ZSoe+k1J0Mau
sanch7NKxZGX62T3LDGBIG5fCo/sGrHkcEAl3/6gFMBWpnNQGiJhDz76CVKk5DGTXG4DPr+UxJR4
uAGk4BUnv3qDuZWerdEGPhaXdQ2FPeg3zWaZxJwS8GEDowWJU0cQNxl06SIBWG7PogHHKJNeSSkP
1pw/IRD74v7XKnxv3D6WqqIu6a/v3iiuEwMZb4/w2H6+xPdeevYPO6bbqiJC4Ksyct7P2aAM4ZWa
Jh+v4bM6dXTnPo/xCT+m9tIupL19oKdBTOpgQQOrNfjFbBCaaKKutn2f3Bhv2qg/RX/M+SS+sx+e
IhokiByEMe1XkKYqRIC545pyzZ8sAGPGqcCqJ2oT5sjWSamDRDMjJHaZlWd2j46Pfls0r8iXu4EX
lajlMuDKmJ8g+Ga9ZZOn0LtCnD4luvJahYzRSO9R+0561ARGVT0hmWZe4oBNWLuSfelSrvY+Ue3+
x2d+O2mVyr2ZfRla7F+svIftCm/FPqLUP2ja4cJ/6nt36+j+/8ryxyiFPBc8wQCkz1E67NYxD13C
mJjK7UJxmvjw+iLqimuJZpRL10QGh9OTopTN/UJeBcYBPY4c1BYPjbGg3oEl6Rq1/7hZcnT8GIGH
VZTcOh3jk3LdA/tvXhxI1W3072PXX321iWADY0RxeMU75Q2iAWsVr3kbbR4JKySpHSXdjUxd7b1R
V75J2x+7XSluLotxqVvmminrHPNw84UML5p+MZM/B53fNJaYcK8Hly0lmo0LPqpV9sihtBltEZMa
iPh9HcfrV8rlflPPTKi1XcgPmi175m3OqZ6l4LLuOnRO7gKKyFhvWDkCkY8XY41/aS05qdNNeAkJ
WFTMaH+xDMmmWCYWYtCbs7LGDYHatMCT/h4UPxDFER/D+XRBiy12h9ZaHpaMyt+bg65Mc4fhykYI
620cCEOxQrddskRJ10xzdAhoM4RVBrmLhR/GV1nDYS7upYFCycT3tDepmO6zh3LOn9xjvzurKcE7
9caBc4wq5iGWYvXpG1iNbuThm3OCFOLXMsbZk2zzAzwk3pnAYHIiIjGfs0zpmBlm02Js8w4zL33F
gL2JqaiRAnkPfYhJ6ixSdGiequvJ6g7OYtPdd71iFiN6IE+f/zBi7jHdYYBy31c1mTUmCkRc0Mqy
4+1shzBL96qxb7HAqeYdbJLRENenQrQQ1jKtMQDdKQX0W6PUFXDsD51cQ4WLWmI5/Fa158Xx2Vs/
P13XTWvNGX9D0vs65QDmAxeQYovYAMYhlcvY6BhqgJlM6cPtQpPBJhp2KBdgpQg7RjHPVVZhEp4j
/rTRamnkbvr322mkT6UIlAAbTd4qPb9aMPMSGJe24gSNyNyfl5TyN3eiOwlsSeOIC8ECoWK+wo3s
vSsPuYVmU9kM5uW0x2Urorgv+5gDzovFWf2/kk5vhs4mxl039saagUUDbKbFFVwZVfkva/fZcQrm
ouHqVYbtXjAz81oxmpyUjno/JqeO13E68C01N+kCNBZDRIoHsT2Hd9sEbz1IuD0PQIngiFU3/PaK
t1+8cevEmED48pkSGAMMkhP9dl3fRnmpF0FXR78qQtgRauuhg0D9C8e3RrkROBy5s3Oze6wkw3tq
dpIucoXRYnQdiOJ3B6PMPKDbhqh4BmukqiLzH3H+YfMliOcdWB8gvyEz0gMOzp2wlXOwoq6oXeBG
Nz1MeIFwP2jvnBoPFqC+4p1CTDZQjN+97+8XmZ/W+scxkYnd9+tbg8Am3c6cNo+Y0FmwsNnfNtXQ
Ib4ufaFXZazz0uEOlFZgfgPGRuizaDNNXvfpBfrQ3kWP69RhGBobguqc9xtI1eBU3V69uW/7x9DX
3tz/vDuc43mVRk8lhYJkbMF9Kw2+IVKLjdUtx8MMGPT4tRmFRDBLYSYxzZUQ1azmhKRGjiaobY5q
qkRSvZRKzYV9YEZg0FC1jpwYmQl8ttbMOMwnw3GwebS18Feb72YDoh/4OYnygpkt9o95dBVzHSSl
RcOplzKSIyGmD2TVK4rurSpBmK9OzBIAVMOoJaX2Mpvc/GL/CecZudT1vQh9DzSg6dssFMmL50dc
dIX5PwkAbaXPxrHWu4BFM486hCC+cM0rgTpkgr8F1h3MG2WKzNB4szxThtASmcFAIW0S3AZ0K+Ll
o45huFhpIpPJfRdSmgMNZfl929HtoJ3OfDuqPvbi265nkPuPpLiSiTUY4Xm/XmOgSQy/SliSB2kL
7v8oJYVnHE3VoUXvhNJMSUTtGUw/zmDmlnw/9b4wIi4Bp2M3+DIG1RNg1dzbcUMxYEexeYvR8iOj
wbdA2vc0h3W2iFV6tGpm+gIOpSxFJG/8D4dj4UPmYpE/lrxs704nAfvVWmU4W7IrnyE0JLm/dN4s
2LvMGb6KUsEK+/5rhtCq3Wmv4XCXl+apTTtWfIVp4q8xdW7R2M/gQSqSJlLpx2o7is0Rm8N5dQDI
RQmO8kC6OCu/+HsM2/ixHnLeYdkKUUknxol4KudjGyz2ST7yjxrw+B9mgk+v5qoy61ry7YNzhUHE
h/Pv5G1xHnnIzVaxCkHaVNEAN5RAwQP8NB6V3VrskTIQE3We6EdBFbS0GC7MS4swy98b+v9krwpj
vzMl0fa/zXe4QrZhTMTdhG6vrkt+smHSpbh6L4sMPya7LKmbB4/9SI5eB8OBG8LYfmz73FEddWKh
1CuWeoQoBa3fWLNO2rur0aBdOih/7Z54wmjl2OMeHzyearZiQYIezYcG6CrzptRzGIGJPdzdbI/A
VC4u6nlkXQfP3ZqD5UWoQWYWnzp+4l2jcyFHsrZGSsUqTx/B1M2TWEjZAghMge4mPEg3bOfssHe8
OkcSjSu5lxHoSX1A4Nu0LTlidG90jXVuFS5NeAPCA2aG3NSc7GaGxK+eM3AJU6vGbM2EeYKzXT/h
HxTwHMWlxdtXjA/wzDc8zZwAkI3j76KqEkpYL981YQplwiQb92uJF9LaTLP4ePlyqqwvscUVRVM8
NgwxiVOUxjp6Q7KxtIkodfu3vz1mXS+vh/yXnFrD50+1LPbgW8lWlCd+FT814/jlLSbl63iacPPF
1KBUVb38v014zR2KAT6PClJv4IugXA3i/XGcSkpS0KLy5Gt+3i7hc34w474EYNKaZEluwWNqolPX
tu7/Uk/b7ccqeUYQsbBh1pUkO1SCrdL+8biPj57M61xgbwbzFcs0iknz1NMQWPpxGJtFrHcfEoti
jfb4tm07GE2WWX/PGxQZlYPkwW/q5+5XFLsdCA6bHaCGn20UeVwoMYaU6P8a1AoCKDOB4sCckie0
wr48slAU6yU//DPj37gHnU8xDzKg4/55nfRqr9nIUF3sFCp4GiAaJARyTl2mh2Esg11seNAY4g7y
1xtA83q7Lg9HaWOjh4++8cClyOIfKJS6DSeW/WhzcLgNEDXSmJp9CoJt7wn2Z6Kmkd1g8iqxINUT
OAJjHNCyRFh7d66C9vJTpqJQ5Is1eYdqGb2ANdVuFgmv0aEJRrq4bhKhT4LFCHmfUfRD7lZWNTev
Zq9BEeAb5gIGQYRRNC9Xfx/f2+7YsY88UGTDIFQB2NIbiMr7jtPn3hMW194o6paK8ZzBruUMFL8N
3xYSLM1SAyeZaRLzbbECQL9PtICVPPQy1gpkqxFcQNKEKCcMbcSY3Ff0RNL4111jGOrd+tkC8QOv
5kDC4gMMrPI1+EN8sFEThqNysp0OdCJpzIV+OYzy01+VgeU5OBCS3s0UevdezGFOYEXpTbgfmXaQ
y+07jTFLkkmqu4YbVGD/AY+UOPaeNFip5DEY7dl4mgiMKGZbptFV8IXjnHlKGRAvyjR4JUh66614
BsJi1Qs1HXAs3sBlal5Afn1PPXCdEE7+1jQIZVLz8OKhGvHmri6bsXmlS8YoHSFaULiGwIgTXTPa
E0A6+XaVQxxsRbr6jF7/76sTWSc83zunKecoHgZfO2SsRPB9Q8ZsxciEDYbpe5N/OFb3kL3/or/T
QGXhK+FJx0LsGUHEBoTj4TD8ExwmNiwA+7JLbfoRyhrhcWnHRpdS2m0F+1k7rvKm/JXRHhON850t
l9/vtRyn4qnWeC7f7q8KxJw0u+uuYArpY1Ui7XT6LlxhpoiDDcuX2PxGQXRvD/jVChCC3ohBBis3
9thdl+4c63xYSfGkG335K1aCSr9W4UsCac3zSHqTTIyH12cW8Wht/AHdWDKjchgqzZu7YZU3pAw2
Iyxw269rt9mtljrVzlft0NYiTH7ZY7vXZIhZMZrGx3tD7xE6U7+0BfcoXytJygcGp3NmhlbO3Sep
NouBa1yKUd6NTqyNJBb6wVB1ExKxeDJGfnBxGSO2x9jXUTQt9kj644o/7Xcr+9LmS9Rb5qFPuHkV
BPoA3OQXgjoY+J27i9q1FMq5OvNDCHHEbltO5L3RTI22LY4K6ispkVsy22gvcMU1LgrTuic/aHdE
wg9FEuSTXWZsm3JHd7pVkUBCxgMBoWV05VjyEzt/sLYiHMtNFHcfQY4AKGJoT/rA3JcDKVdp9o4T
X56fXRpCul56+rmEamfLJ6uRCoOfB8Hu+RJozneOlRNQEjGySfLT2foKzgk8KcYhFQ+XQj7ITndt
74y+gyfCWT60Y9aS7D32rQ37JRQ7V//XkQPt5+b2dTHVlXWuV4Un2kqBTXurEGrqt9O8YR4pkCLO
oiDRv9nlwckKLWkoRU7rg9UqTJFbKG/icm793pxVchkehN1dwn+UfhOG+BRsoZPPLzQzxClfr1JB
tpcCSOzWh4kdLoTTIEsWf3DgrAQDZw4lnefjc+CflFZz+/kkMLDJalL63N/cIHTLZ97fNq40qtHl
Sc7nO1nDoxe+HFU6RQPp3Hnam7ueaTZc9GmLZgv/9aHfU8eFstwVDO4HRVQFVynfoFb7vlOuaN40
jVPGFyt9MGjcuNyruU4w5deB6LcSHhKJdzVaWG7TZmCZQhEB/oGuxlHEaL80hsKcHzhkylN+FTJd
mTreMuGx7SbDWAscJ/LSlbiYFKUu2hXr0EjlaKJMtRB5LAjuSZtwlHq6OgP3gvwVgQeqK2kJVOiU
WSylKL9EBfIwVnAe0kLulOIb6DAiPUQTyjgMbilD4/oPl8+X3epetIFyECj40FKiDGUuAxY/7UcU
eUqMyf/iHO6bpXtuhOSkvxzhpBfv9p9S/L1p8AcQNUB7eIr0ccdYj39g/9mnFL5yohSBt6A9qw58
Yncdi1xuMltT6PtWpr6aa4RXMYJAYdc4APaBH/cjn+uYbDZ2r4NRETnEWP1NpK82b4YQwnADN3Nt
FEPMVpKmtU7hskNwU8ZsSWzMM6TXSWP/kfTGnHWAJmCmEP47kFsr4iviQ8bp/o2CBPvNlDZSf4Le
PK5KZ7s0jPC7PYnWtPymUItPHcGKk7Dyod6982sivyuLfafEpM/WAtorbsYFauabGqGbMr4SOC8v
oPVhZvwx/PG5qOmWjV0PwQX2q/pL3owX1XGlBHHGwLtlAY1PpLJEg7jb9BTMgocJHPMGh+3FST2F
ZVI8gcnLR3f2uUfbQbhTqDzvHJrpwA7uidp8siacCRXh2mDX2yUZNopwFbFfSapeeIeHRbOtr/Au
waObMWGvXDj5J3M25LLsVkeJFwOn/OBCl+hLThnwJ5TIRDHJEi9nO8D4bGU1lUPTfxNS7NZTpEcD
13zGQGeDL05tzYmTEQbArFMlevMjM914KxN4b6tR4swcgaJ8+Jauv00Xc4yLaSG778HovABMKkcg
9l5FM4tPlf0oXs/nqd4h+27W0Wi5R74wqP3G9zod7yXuiY3lkWReUiF7pElX2SKffpo8x/SErf6c
fHMy8/1TUGtxuS4MzA69uQEUJ8tXu+WVIQAOMlweIwjITPxFoc4fKiupCgLoKdQNa2ixDMU195dU
vn9blPI3DwkLD2e8BbgwJRlrKAoESiDup22Gv3hP7Akz58pz99kNKMwuOpxWgNABTJWYcJ8DtZdV
9uwNd/Dfmge+v7pk2UNVqKYmcBQQzJF/UIP6F2VRcX+G1H2Uf6CnZU04zRcZ9tX4fEEPUNUusz/3
VrtXUpYWQdjGbId47KwH454xoqAvv9ZWE/b0d0yvYr4R8DuD+MUjRaAhgQNaqRjun9mOkxdjuVXS
lBTq5OEXr5Nta69pc+2XBGxMlfTGI3a+LNgoTvd28UymEQ5uKSBcSJN0f2ibMAq/rzyEEgeH4AI+
PVssJ+pA9wrV9hXVpbc15b+fNr8DBzorffQCreFjTCmHFT/HDd+M6RxXdzIl5lpDls6/UmMmu7pI
9mwuSDytZptwMx9sxZnF4DxQInuDnen8KbUenaNE0aUOBGyP9hMB6QRPge6yMYnKoxZUX4B5S/1d
vkOMjFvOFhitdpZCePBfGMyAfyVZYa6fOlVQjdDKjZfllWVAXNxsSr4YtsUQ7ziZB43OlIeVuB+V
0SoiNcyM6mXcqkyf40nMksyVXJP4pTDXcTj83fhzNSH9DXqWOmYEcMllpKhJ2fwOBVAyQZjTPtZV
IVgEUyMr6mfqlhMyMpzeYTUEXXcNmuHYg0tg2AwZI7zVUtgChNdbZxxlMAc49CEaDJsW93nA8/d5
A2hveV4E+6xZZUygW7R1d2FtCUPeDD4CCheXu0xdyMr9DrE5eGedEw5Q/h3cMb1yOstX5fL9kBr7
mi3OUXSulkDxA3mYZ5v5CzSOqJk0sSN0KdjTMtJBHJ8xDcvCqYPZF+mSQjVbhj1YnoGzvcnQmaE0
HHrjtsdxgrTDgcHayK9BUNxIEKX4lwG5BaJ2qxokbVmH1+R744+/60EctyGHD58hj0Bi7qrqomVN
zrAU3+EkkKGQGrE2ZnOECiLkygf9VeCYW2OgljvZDgFFeq4rYfn1PDddmHIrXijd3DlYRVE9K6Tv
jBh7Run3vmenckk0LiWu+pd7+Kx4K0W4K7dxE2wpSbTyTa6pyseBy7DOfHNNRx36QFcQIByVr3aP
3DcQRPVzUbJIKi4DN88nUGmXoYgtBR0ZkRVZ9rzCH/T78ZKo+KLI2dYjHcyirkWRCHZkDWBwJOiW
qCNAedPPb92chV1UwQ2r8j2++ZVjXDBBEAQRl9lAFdxn8llU44749E15NuJeM6OAm4q7w48m9e0g
hTsZ2wYjGtH+5fj8cP4VfyY1i621AXpcJYiuUDxzjQnLpW3Xa/A4KdSk+wVgYk48ItN4XJBY96jf
1awvtAs6kK7CwCqaJCqmt4qW+H9xpcu8p7YcS88nWyHeUgZP49FKeKLYnBwmpp8eBATC4NeJ+fPe
On4t/SAVe9hLZN8MPQVFf7jDkmc7FxnZY2Qgfw7cAmnu1PQfaXM3YJtDX4lLhIB/Q6GOkykSmbhG
730ohlCCVJhOX3Akh3+J0H6Y3539IdTEBkpHomst3syt+kZR0ax7NVSiAvRkAbInVKhaJ+3IA6mD
+nJHAGWtNoAGCVbyypY0Ofj9M63kR/o3zT8dSGfQPR0N03YT4i0J42LMlxk+/yxgvXo6lIH5IDvO
Qh97rXzih7bwdj9EGeL+1qWmLYNzQUnw8KGA+R6labdI6HGpee3B7A19kDNSw8RBhh13N+c3OUZv
dogw1w3jVSGQqdQpBM5J1ZBjRr9SLVVQOm8H7dl2HdrDSQD/CyKwYae0wERiRLj0+uGdqrx1mAe5
pWv1M203fVVkZh/VW+KuuXwIWTdxqs16B+3cDBE/a9Fissk/vat4XWr5BIVjZWCQYjUQhYU1PKdH
93r19COFaPhU/hUMM9T/1Ryk1qU62yQwSwIVUZT+uvYLGTTatLNXxBjzKFc0JExCkttzZWASqHw+
Bszj4O4zAs10t3ESwAoCFOb36AoI4MSnkBtFH07fio7Zn6hPS2QE1CEivNADbUlpEtwW1GS3O6Yd
+Gr1wfoba9Y6+Bi+gsvtysJbgCHcQqL8vrokPC7NiJM70sdX0hrmMTNk07rVkqfT9IEm+RI9r7Z7
omUuPPgatBhWwS7Row2w4MBc5ljiM9LOh8jIElrrOCFh544FWnhg/PKs+JRBqhAQx3r/vi2TA2Mx
gWVJOBrxeoyHqSXQf022MxIhkDH2S8EQsJ/t7waZ+KnNSo/EBJgqwxIy5EuI2ouhUzk+swoCUwzC
efB/gjn6/qt8aTqmXxmQuM49/ynzym0x4nLyVp6RQNruK3Fs8w9ZFuUP/8W8zKfXq6Kj+X9cQmkm
tX22MJ3/lCkPMaZaq7twy0Y6LaH/QKrHMsdX1Eo5EX2s3GZASR/SZd85ZjZ5War+JnAe3BVo9Iwc
QZIIUuOodlOVmyihlLWKkkPukVJOyrm1+m4+01izYPJhA6RpihUHLUjvknQU6jCJT1P9q319tB5i
azUP/JcK9Sfjm17kqSeq9gg+mQWC9mOvNDlZ1eru8IoxTwPFSfEdJpQjP3HnlBaI0OQh3CFRITwP
rEUw8/uNsmZT7H4p/FNW9F/t5kJBqL30MuulbH7FS7wpjVjPS6qMZiMSlp1W91vekCr/1niI+hoA
X/KjiD+dctzrKTl4qrJn4DsFSGxw7EsnX5zVAUMnm+xWlAJ32DexkHZQgpLz7FrHDx3nkOBiF1vK
N9yNteHpGDCsHfen6DT3r8utYCm2nnppyiXaqbQ3GxvEHfMGszAg7JGDNQYoXJFELqWJXharr3it
R7nfWQWVkqtEtT77oin+y2HE1ymTurf36XWyIrvoKt/fMj6Z8nRgBkdGw5P3DtwMXGlE8VDkLRfR
89WhemyvONT7+vhVdhWy9Td+Wufg6pwzKi8PGkgRlzG159NzYaNacieLZ7/289q1ek2B9QQB2gMQ
p14FlRMU8OjQAMVxSrmbD15NaykfbNE9daI0DYoXwC3jDh673aMqoKZsyFv1jzfHPJFLe/9ztVai
2+yn0xOmJ6Y5UvPskKemVBhMq2MRGg4Ts7ZqBegqt4do8fuoFw5mmUduEbfeUxA93UKcJvb6R7sU
DqqSNGHjVkfVVyfFi0zEh7YMODA2zIfoh0WYOPfVNHVuaqX4kvFZNLWRBDzJ+KaMtOpUNPypHH45
j9f1nUb2prPj2U6jgpT4YhyZJaQRssGzNly/S2KKcXgX5F/sC+KlnI90xVv6r8oVdHrNaGBfLfqc
qe97v6h+8KiOSdJCPxGovxnAZ5AzLHtEQbCBG1X+eF0MOLNGLSmFV/nG4adagvPnGyjBCOUOc5eW
R7KCrMgPYbXspnQGW9n19SiiP9vnnIRhIenqwSWKeNQrNovIUUc2Iwa/XGphAmxrSKIkU65X89Fp
dIFCXOawUEbaV7bALB/QC/QlE6DtgYvVgQKVFGdZCZKeaHpQqNIC0vbJE3Cc7g8InLv/3fyqi8x6
wSRvgaRh5MqGlKDu/1vhsHN0X6lSU53PsK4xDGgLiF6IwpCIDuJ0IvnBSXEY38X5bKn9And3rmyD
YBjLcWFl20NQ6RtTntlhsxvqx07ML47xeTonAyaZDIoaw3OFqk2MiElzZ0HxAk+QGX1romEbPv7j
ZXCvokKy/9vbdKryZG7ZAwjWUcJ5Ilml9Xu9HQSXjWv91ujv1UtbS9HQcNxiBc4PXZMESKG76c5n
8Nn/D0FlAzeEZRhIESv8NvCMTwumX+kGzsMzNcSSoyU5KUT05AGCmFXB1QAiLsIY6ISZEx6+j5xb
+3xlz+W/dDZHbuW2e0XxwvuQc1cmiRlFiIF6nrGSW3dagA+7gE+EM0mixh/YxVZR5z3aPcK4iqM/
qWvattHgf95hRza4VBDZcijd+ENwsOuQCDyY70aAxCWR6AVqLiS8yN3USdvtGfMA3iMPKalUWAWD
KAf2zfyhv7Ow+DWWMSrHTHaGSLNZkPb5oicok6btfx1PNuzIQzidj5KOfqEdG2nNgwpLuKHQjeAn
/CQmH5ne9Civ/T9F9+BydR4YksrfFrPYqDhBS1YNtEKJBI09f2+rNIdHuDkKG0NkxLSgDHhr8K6I
L8t6DwpMFL+0THs2OiL+XWNbUGoIfj6Rf536HtiljR1mb4saVWxCjNjKFTbluuB2Tn58TlFVvLu8
QlTbDUct2FHsv6vNl/YinJKmb96n3fk6ksdl1PxrFdTSlQ+jqGnbBCJLFwkvIY4VRKfG79Yi2FEC
OSYUoW2ubU8/E0osvj8PQS57osbr3gOkRIPa+NO7XHKtf235XfsN0bUZEmTT8S66zBhKpi7ZNlj5
a6zaNULdeD/vHK5W/CU79qIPTaK6d0ziQhIZ/k4ttMRdAkzXiId4GUcbp8e2VIg/WW7iL7muiLCm
L2bIzbgR/neVBm4TZUPuojxkBQQkMJeAEkeF+LKuzmWPd+kXyJccgNu8Cfl+83K4Xb7pwLkxdN/c
HaaDQXMBsCJ/nW69pWhnUO9rIqwSYcvNGZldgm+aofl1O7z7w5WlJzI+oi1X/WyO3ocTt+UUzX6f
x19v21lKhMsX1h2U8ZvVwf0uJtjDrb2Og6TAZjNZkWWTO6NRjvaAcy37hYsdbcrR4Y5OEdaeaKCR
joZ5v9S287iDv83BMD1XoZLMlufV34Twh6nx8MawlIW9u/8mTazm0D2BIFZFgtFBYct3KIo9fWRV
WEc1knkLK46RM2Vgwq9qzTrxmU4nYaGXlcMPNEwbGuDjm4gQLifdcgvTSSDgM6l5IA89L1FHEVQ6
boDvDTsgh5rOuGkRpHPtKJAK/Fw8c9igCnlsE0/YkChLRnpHtJe0xhPxBs03uvmctPXR4ijN0aiy
/yPEI0tToFxTzMcs1aw72fpZ2wIuEgxfrzJZmeTEZh4Zcwu7DlWKAq10ivARZ7hT6rSyVW5XLKkq
wxXOxi0jPf41ydTWwthT5Mc96ZhqEkyRp/AioUwml3j5X9Cc/F3lC/Fj4yxi5PZMChU8KUCIiQr5
hn+LHKGW9AKrD832GcXN7EuCpjiTLiScTF7ncotpCgCLkrcVPDv91uX3HpNhgZhYUcpLUJe8MCJg
EKaTITCC2kpv8BfrDWF0M+PNnXxZd4SsHeYnaR3QFfF4pSxpEbqFZipWrpGrndI4IDfCNtcMTuyC
4+mAR0LmEzAlAZPNCq2mj73MtVc5BlSH0nYkmLqTdkvyJFQ/nLFNoJFh7LR5GhZGvCeXjWK46eXQ
bg16ULzhov4qazjaP6f0dkuiPi1AttTPhU3sv/MAJVAuA4mxR5ZWLBilCZQkKNGtsIYfMgxQjpwa
zeocACDoE9ODWSk+LD0/S82HaSY/t07DPPVVn6kEQu/P0e0aZQ38RjfgkUALhSy2knqdPgQDUEHv
JSTpURIkDTVPP4o8vwpF/4hXm4KeOOpvTBZPqex0uQKhIMNpw1z+Y2Ohflm5HrHEiXJcpT3F+W9v
ZreHBhWiCmghmkJwr2Nm0OXHfxfUmGomenXWsXAi+5erHXOhe4I0Pm3+Tyha8AMmJsGsfAzjLVof
1oeIztDP+RYDJ/pmGRagLVhcyLO5ynpA2UYZzkQksJFJ2e6ustFNKu/GhkRDWtQhB7aaYAj0m6Co
nwjARfh2afBJGM0pTze9aWQG8vQNFst//0Mh8YWyxP7QGKRtHmowr0toUPOH8hLue7fWCNExvoVl
AiHG6qH4MsGw9xo3Jx0FnQH98kjfGFcXZpdnxZe5khB2E8YX6WgO9loobIf9SqKGAVhuiwsKRxXa
2lG0xz24UkLY0yWe0mEg83fz3RpOJ8tGOsTSPZ6Y+RoQ7tjDN/rL01VmWL8LLlMtT8AwXUK7xr2T
KAjdIdDbhd7FuCcn3siPkvfh3iWOsh/rzVGdQB0o0ZPwTQ/Hs/avcQyyigq2frUK2TKrSa9L7CZ3
M0F8sB35bPcSia1AGoI3t/BpeZQZcHQJUGmxA4qgvHTVMH6AfYRoXNAnjuuG8ZzAnMMvTKt6Hsx3
IPgkwpgP74VDtStDv0DyJkJ1CdRIfLyFm2NuAO2s+jxnqQJ42aFOAyM5hNEtBCtFLOTGtNmc/Wwj
u2LJ+f1S3QJULAnht7aIKHkvtJwWQ+s7JXlB4bjIZ/4/Mz4TTDKMK0F6bZmf/w5qwNyX4ocIk6sD
bchXpqH9J1QrlPWQ/R37fFwRIn1ID9SRGWfqJWS4en3FXLU401cm9a+jcx7D08NLcx9CL69PzgPi
7i3NcmsOj/pK2FaMRDKxYIA8EpC25UlBu7aHoeKKop2Eb4PHCQSvGfUqMJ/qylELG3DshowgmEag
VRddzCSsbhIM6XHhlDTaaKI0fnoX/bcWXFf4XT5pq9pbjo/gCQNqN8CkFejwEujMR3H45PeEchzh
Ned1zbnugD7HEegThADX/O6uYFQtDgqB4Np4NQmJu4DeJEvYRpDs1WMyb8ym2TRggGp+CFbjPQ2o
gjrbseGkvTJyJ/B8lBc6U5Xk7gTTLpDjktzk2ubdPQA5AZzrryG3F1ev/9oVooZlBrfnGxUuC02l
dsWL76gkRBAjSeIfcpndCnvAkQQA82ZCdDQT1pdGtd+v5rPbdaCQTkqzbffAhmVSiKiCNnOgJAEy
NyskMmBqWbkauEN3YyZ2VkV5rXOSkdZv6pDFnrFrI/luSDxinveMFUfgH8AcphTS+Eqy/Z3aW5GB
SfYyNFFiojXzVEA3K+JkpHACeConVK//7XhH1RAr2W9iOb2bSynTW5xb7rTZ2ufte4JgFPnI70x5
cbPYjKh1P3gDITHLGFbSvE7wrcFFkT0KmKSDH6hJZzSm6gjr0R3P6MJEO+azFsS+qKOj3bGFrf2H
yKM2CKQNdXyfAR4+jNGKuOoMuNV6Oln53dY5W8EIYmeLV7Vq9M/ze8TF8RWw1MqGGX5fE/gz0Ctt
hJCGfHGymxlKHyS9cLwo1IYDGkCNC0iGPQr41wYI1t6a7JDgZw1OEZouM451j8oaEqMD6N+D0zAj
hnyprQS1K9eOxgiY15cbjdOVQEz1KQQqeWBAe7M0tzNgEj7/UI6LFr6BwvvS6ZN8eRfR7WUJpok9
YbBqj5iKksJnbjWJZw6PfQ1OyjSeOtXnVlRASSMacQ94IkxbHZ2KFLben9oZ9YUbX25GQAx726nb
M0SFEx3fEwA/zZyO9LblYZeKu+PGHIrF5hT9H3QstxAA5kWrol80KCY9Kj6rCPlMOFlSWwNHM/B8
v+ZVNeyoHD0QykjKapLtZI8gVcLDDXpwoiKliLpCvFZ4xUULVmT9BfzNSNapeoqS+6TwHpvRVh8B
SlKEmLLTaBagj7EPdvl1E6CGSGzJ3coXazT5BR/pEcOZSCRvj5eOt1/sMNln7+9WQBiCEweMwCpv
9++KNTnE1EZFjFSPtiggD3IW2VcbMVJ5gWrt8G0ksFmoCvQGTdraIMXWVlB2GqYMPgM8prMaRzAO
EdHjXks6Zgn2x4FHSH/oT3KS+YeiKvxGGwkSsjAYrROJh0NsHVeV+Z/ZVBxEO9OygLdHYvDhZTA9
4oiHVWrzgoTVRqSM+oUL2HUQZwNmXK+fWmeEghrj6v0fA5LlkzMGLt3n/gwv7k0fJQbKDQTVLxcG
ThSYUvEha70Fn4s0oRD6SwXg84++cgSOHH9W/3krbjLrF6xQsWqxmOVRKAzsA8bASx5tnUpPVdji
J68skxOO1SlujFueNIfVHj1boOaYXka43KEtvqQrbvIDYh/menjbbjNTf4ax6D24Mk0oTjJagKpJ
M9BrhLD7FaYCJ4ErylVPqA9JL2iSkxwHm9x0bdhvT7Rao0taP6coLpy3ZymmmPBWQL3hYL0QJ8r4
KXM1y9CRAaU8dQxnZDZRA5dDh2VyF7mFY+/qhFDRBq8qcKsB10B4NKUnItxkwvOScP8qTexy5ukD
0R7W3u/PMbyPcmwzQ7qEp7AOktPwMayWvyoQvChqRe2WMTtNaTvIY6+vvm72iESaHRJQsmD5op5n
0C/imgHcSzzWiNk5iZeAylKu9AXLnZOSEKlXYV54ABcqc0OoZfCkjUM3p/WCP3kbVnhmfjcJxWiB
bLrgF5EOJhLqPX/POjjCLOcqNLvL3pX4M6sy4cYVdvkVZ1qKVvvUG9b3UC+4tuLZ3BHRNMfrCCt3
24kl7pGp7Y/UHLMPRV2xFOfqDxwIuuXcHFsK1qmb6+q+fCY5SmAWaQHwCpdY2gwifJr4n3kFJdFm
49Fynsi0oUHwvO6h8Q9AgvTRj4znRUuFf4+osjLpFL8GyE8inK4BjU+r/xncA3ThPvhi5aK72CCq
4Yp+R4jqPGPm3wkwqZECn6S0SQwM/K04PpKDN+xYxlh6F/LR8teBOIFB2HVVnjuy0FxCIkTt9bWM
M11W8rF0POQGKsrA8SS7+g5NPb5Io1HZiv3O8bjTL72EgCNmJYlgd/RCn673MhDj/G5mxGQ6kIya
vfHuMWioLO2B8rw9hNPgLpozRgvE+QdS3fXNF2FaQLYj+SiA7dI1r3l13TAF3Bd3uhoY2uUQnPkW
hwF7TY22dDwa+3UAbkg2NKP5oEi0JTvVqJV6GyTq2Wx2ZzzpF69hFtFDInR8X13XRf/3eTk5uzUA
pleejVBTbunIgkE3Srikf3I1kPI0/7+BH3mLHceqvqg8iebP7cZPFcDzgJn/RSBlEsM1Wl06ohYd
nKrhH+pDUQ7UtdE5Gev8p8qIpAvqSsl8QQLSluEHoLQTlD1xj0R23JE5l5vlXmbnpsKXqZVGJ3pi
UjUJUAIG3SQVICcqTLdrYIX6MfL+nYaatO02F4xlty4yFs/3JCi+NAydPgszf4eh61gcHHYNXxdl
BJZmTnIEZld07ercKhftxKa/+p6oRjDcL9Am1d1dp032DTgCWjBkJ9Ap5c9bstquuec10NJNR++P
R6eY71rhJJrhZur/+QwOAYED7qCa+a7sC5XeMdLfC5j43caWL1BtTgsrfP3+S4z6wy4OZJf1LDNh
5FuKPR1TrRQS+YDyITOY5FbvuwKNR7echyi1BaVKkg69ZUVFvaUb1zhAp1MCudOAd9g/3bgT7SrV
WDfZ4bDRKWu6UK/leNNC82YaNyk2UsfMjbAOMnys9idGvAKnSqx073NQiAsUTWsEIq7/TAdwLUWx
2xNW2y/Z0wnrTzXtQCl92rtcaVPzRN5VGmGZXAdIGMf0m0Ehrculh8T7ixAzJ8UIdAuzESdGIA0i
wvZx5ryoqfIRzh1aR6PeHPZv0qiKy7R8Pm9cDYSHznu6WR6AVy8a/a4pK1kvg7hZ3sQSy4zjDnCG
vgqRJc2lBQB2sZYgGhFUJR4OWHeNX1xMOcbPFsovrgUxsKEwAWsVSu7pkZWJvJg3n4rrFKnjBQAP
r+SXH/nc6MFN2DfUKArmDJBQDws0K0bqm8xCVg8GgQfvMTvQl39eDzOjNG8Y9QwCDlNuy5lHYzJu
iSwl33Gw/lWesG9PxeHj25+aGSj3cOGx4QWbFawmiAkkn6cF8lIRYEJaA/ZWA2xOx55FK1LSJefM
aTo8KTDpaeHzvjY272/primqs813QG38CmE1U8+bb+u6YeodxWCpN9b10LCMK16aR0qbvU+w9Qf7
BD3a+FjyIl3YOAeuECZnh8u0PJI/+/OPt4GMTZKryszt6okQhxLSY1l8bM22oQiHEnA7WghmmhI5
VCR7/6juiPXEtqZi2Wb5m8DNq+10p9/dvr2THXI3ugi/7ko5xbSX4yQflGi2A5CpPYh959L861IP
4lH5Wp2E1OV/RDMSxNCRJeliBrDE+Ym9xna7iRSR6r8W8ERQEa5AQoizpSv+U7STBO8pS/jOLyQK
z5G9AfyG/pUKDolsL8cLOp2nZK6e+/6mMby2dHGYtDxmYILHU9t6hqs691dF2AIoeI8juiCN+1rM
rNA5DlGpo20SRTv7uQCJDGHJrPW5SO/CQNejYvNJevvv7tqeO7LJ2c8PW2n/jWlkJdpcQ7DNhwvx
TYKaCYzGbVVMflJYWl8CzD0C2Sv763tHuiWkxkpVl82AHU+22Kzx9T2VehQLoX29DHlh6TwNFKYW
a6n92Fz0vpe+U3wQpeGqhGMdJ6yhP20urRu7QK80Ici7LSkLOwWig8wfwZi0I6VIy6rFNuT+nbcL
0wZKHpuLtdsJKkF3bULOxZqiotX75VOj4/mizTiaK9GBaKjXh8Dr8LIIFvDFz7PspMk/6LXY8SQH
aMkhCQAs84i3uNb4Fjwt4dc94g66pmg49TVysMBpVoUAPGfwNOiQYrL9EgQrru6XgcY8d0UC05nM
Y5mMFLoEtF8y7QNPw8n9y9rrT/yjlon6L2PRz/hiKPX3VFSmOSzSGelc6uxdqoz5DQh2su7mT97V
Dwq6lP+paaOlnIqoabFRZaUkAqPm+Dye3vokp6lU+kRIQzCgjrhCXYfdAvDmZDJD0Il1ELNMDty+
GNdimVFvtpec+mnbORtYqj8dxGnPRwJ9yRgJ1cOv/9ggt+2ltDgP3peSJQd6vans3lCUAx0uTYA6
dJZ6FFvTvgUhynx6Uh/qdTlgqXckoCTNs0tWVSus5e5MNiKJSNBNqWOJnY93S81rRWNuakgdQEye
w5BXpXQMHlyaoEArb+YYqG0D8JQRRvW5J0W//WyOVN93q1+43MFFfpqiR66mtufbde16aGalDqmF
Ef2HCZAtN1XN251v2lx5roosQ6puxsHKpITliCVrNuhUEFP1/omASTfuRq/2VeC+42XGOddc6foU
oBA2vj9KP9FQuvKWWd52QDzxHwRTPM0LoweqdNrcOjBaeH3QiWlR6sGQz/W0kHktja1eAe+oXE41
cxVsDFJwyFBPsgOLoUfwvLRetMnX9JwUZbycoO+uP67tEDm1VWvNOVi5flrN7py88M7uADSYCBWP
AxnbrLtlhkiXZTVoy4tb2xlBPdqXPgb1fWTfWgSTquGbU3FQbhSC3DwoWxwzz9glWAvJjJ1US24K
AoZhaYBWJdyN8ZUbdXdPoqfER34hjI4jIGQ9L9Of96LnsmAtsTjaLH1NgI7EW40R22w/i+JwZKnv
XBUrF1TvcDBkqLxi8fRIXgufUTHQwr4WjfuvltX12ewsJvzmxN7TaUteO5m8rsq0op1sT3UbYeRU
ppgvnT6gIKFIeuL8/JtXMtm8cJEGpZgh0z1V5l1bNgnwDs1S0PcDqzn8Tv/tHqEbrDTbokrLHlxT
0PrIAW07d1p2YW7M0RVEFEF93ZGmhkdqZrNMQRUxaXoP86xjYHce16N1yiqcdq8JkjCf2n5PSp0g
xOTL4bOlR8VkzEFwGPg+VX9V5SLBcXvr8Ogpfbt2hNbO1gEg1ccivjRtbOIgWqQIvrU+9orHq9SL
ELAs0nnseJs6xB2fFxXv2xK1CMZzBVRkcFpPumUKDh/4U3TVSzs6z7nqZDGxNez0wIxhyiOzrCz2
nVReRbhLdF51MGKxqZM4DmqU6fu22IfrMZB9TEmWZy5/EZbmvh+XF+OCuAa81TmArAXRXl9Dn3DK
KJSBFb+sOkPkUsi6FsMOIxrtfSoSQBIw0dyeVNS/W1H38aSxB7Ju48jssIyk0fzG9TV+1Wte/zUL
xfMr0ahetSpU3wdo7X8YT27OmQ7jLD7qExOTmvzegyJz/VH1YI43stwfjIe4JzmbozsWGQHYJvXL
CsMeDa9WlYnOQQVDqTaXuX/m14bWw+8u3kFy6HRf6wEMnJUcVKWH76mGbPelJt2+95/uyg6DtWa9
AWXnEpd8ycBmX8sH4jGxEgdMUXdvNOAhwpq4WVgjGddUrrVhukV8QhZ3+Zx6Yj2k2o2/c3n+tvHd
1cR/4oyrFsNN04EltL76GQGiW6iGq5C8B15+9n4AQz98Q45Z5m6t1FaUv3quYsAJlo6J7ijWWDM6
wCcS7nZhBbZe5rbDNIYHRKTyPnf4w3Rg4Idhg12jVU9MKiVJqNSh3/S9F9i82UbQPqJm/Foxml9V
RE0sNnDk0ZGWqZr9O2lUhWt66zi37BS/A/Tb5q0kkvXgtQEOeF1CX/uhpMjS3bgM4FgdMO8rGzQx
e3NHpY/21yMOEzCXV8NGSYJ0e3X7eSwol7yn2ROHOu2i5wJJUzrlR12I1VMQC7kOVMD7OchvbqPv
aaWLPhUX9R5opaGxxV0GYLU+CCuYcNakrUXOKaY6LjKINH7cJdiaY+l5HNCCL76GJEtQ0CL5ErfS
KvcXF92PYu/MERW5Y92rP9Dh3VRC2e2znbFERyYY8V5NHIiooBNRgjsCBdQEPNY8w5Lt9nZau+v+
Fd/TUNJ/NGHjrEG3GrpzfkH54aNYLbnWJ+C8IvlA5DEF6WKf9WH0U1p4xH7UKkEzDhNz+r6MgT/O
X5XmdpzaBKx8iG/FQ9roEjWVDbes373HvghzC7ZK7+jp/fa99dg5TpuX093rw/NohOuFlJcKZ35o
IeZPCdUJRRoPn1v1W7SWfg72OSzqDgD4/V6r3EZavs09Bm1MIpxPaE3IgX5gXHa1+XaYlWMZtk9s
fUqbGkh3kErQa4FDO21tWdj8r+msoeurklrz+atZUvEHeVG/6lvfnzwdU0B0QTNKJp714ST41qbR
JcwHk+pBEZc4VCsWGxN4VekA1CnplGCXk7Tb4cU6TenLxihz5PmBeqRgS7mVrmRN3j8ZUJ8I7mwc
w6ReWKCexaE+ds2jrXFmXarMdhjWijzifu6oj9HNlUq6JAV90v+DQByUrm6Wh5PX9VBIkbkxDpa7
OF3v1ktBlFXys85KbN4tchbr+SzE+X+R8EJgHXiMxswu2iRgLV1JvzgBExqV009WJ4HExLGic5R+
uoRxJ3vv2C3iMQcch8ha1RsPRNzDhZg52BTtzSjFVCXn+6K9KA/N72oz5Ff+moTa8XgyjmhHPUla
ZvmvbnN8PqEuisffExk4nLQ8eOk21Lk4syPE1tYDsvAJTCEuQBa1jT6pmsTpCN8zckBRc7aNYliG
AC2Q3fgRNxHUFene+ZOJUmwCab/Zkvx9FeKC7YxG21yiYkZ15VUVAlyudToHLPVFZYEPE3QF0Zw6
4RukAReaiiuhzIl7TmbfNdO0rs0C8Bk9E/qzzodjhK4CTviqm48BLrXvjyKHCxL3pmamZquVy+fm
rBkVjOxt7jVLu177AkNxTKF81L0Qj3JzzlZViyE6RSFIqAYq4cG3HAGXJKbOpNEWux9jsD2zNchj
xwKq4wqFuJVGuIc90wxwfUWInMBIov+AqBZrF4ZroUPOEjr37vmrM9ZabF0cvBhCJvepVLDULG0s
tEksH6gtJk9iV7jxyrSHe49x5wlq5u1IG9I/2+v9OTOhfmwGx8cbhW+2C2K5tBintH3rZ9hSkUEv
80UyYEXBUCgY9yy+67l9SOAEgWEdQQhISXOx2tTVp7yUZJ0LyeR0MpQFJUQrAVff6B0V0rq2gQJo
EPnmRqjSm91s3agcZu0D4TfFjpAXUdD4onFYAD2s5GWMx9UdgyTwFzFbHJt7x0v9kasYvNh6SktE
lRcG217POEXD9HfO56OgvXqwjSTd4QpBxm6sAd4PShObxdU2ffAvtxNTV3TVgEEbz/COT/40SQSV
wEY9LMeP3LiWU0DQUuDD26i+2xnuXW/RAtk/e0g714qh+FNsiuSzILzyjO2oN8dJmnEPE5fnf3uo
fE0KcrDsHnzNeExYpxBCTz4P7LfzitwldRsKRvIsXwEHWxIQc67dJJYCaWkfW0n/WTFBLb4q8K0O
lSVSdPSqQ5hik66pxPEdwKTmmXFgNofBc4kGSTqPBzf7E3TiQYzAUF46Hd07S60RMQCufRpIASru
UzXl0VI08kw1d3GZj6lcMBWtIufT/rkqxGaHpYZKfgDEX+P7lSwZ6rWmSwZGBzFbFTTHEm2e1Z00
kcO7zrtshXBhzrJYqzKdXN+5PFS7SnfLU+pWDl9dBP+RxqYrEDCUrKSE37bgNw6NH/b5FZliYPNQ
AUIA2R4Db71rQ8BbH6VYkDx3YXb1fZM54ZNisbUoAbBCCgHXmkHF7QYfkDXnPRWElIvIy1kVhm0x
SRqqi4MSGIF7y/GK30goRhW4Vde2Lg0jltPMjjqxDUd0wjxtCmVcZhTB3N5Jqec2KCI02JPTaglZ
JGXkPn80RhT/PLXIdXnzMfUIhQe16t7aPzAZMGZwHZAPftXDnqMcR7l9WCq+mGlcgiZmnRlEt2ch
R/VpqmOHFsR1lI0PNnIqUpxlrmzPbuNSo9HuZyfF3hFYr7o83yEiGOE5is/7cLlbf02jw37MiOzf
/FxM/hjVRoLFGam6Q0IZefZ6QLYm4og85PRK36+T5cnWfVssGrU2aE0ocQH9ZzWduy3mOpGkNd5P
Q/woQ5D/F5jzwGwLKn5tC3/hPavvW+5YJJxxOwzbITRKlcZexp6hPXKr6J1BYBkPYYbwHYS6mHBu
QUJwz4sb5kqB+74lUaNufJs8kieA8zA0fHAXMragL5LTgFQkSpin0PdmZPKxoX2QJyaDExtt5Ny+
PzBJAmh/h3n07Iky57bsn5KEuX197MuV5wAfe6kxVHUiUNUtmkCZ/pH2dY7WyyIeRwOvL6LTlWDk
omlBS66tK4U7DgabDTLJUFLocOZwF3ztoJmbsSl/aFl2Bo9xWKfqvqWMgmIlk2VaZpKKXG2eT1G7
DUuw8yFG9RE6RGbIGm9tJ/cvxeFrF8bqdTJQa8/mRkg6prO95MDqoUFCpl7LUvTG63RiEJtAUmZG
1Rpdd0DAmr9Zw7urs96kI9l/dU4za7ZzTZPDNkSjj4C/dW60B8zCOsrBw9sTmVOUmsSYzk/p6J6l
jqlwHQYwMvLUB9e3gZFJs35uGL9Q0OhK/YVabuFot73gZDTXYuDvc87NL5eDpglBPY3+b72OQP4m
7vL8cSp9osYSeE/eB0ET9vi+equDFvzGM4Hkq8RLEOCHDZJNo7f+tAqVNLE0BVRbHbAuC0QHrlRZ
CrgfBFajenN7l39HuB2JhM5mg712zQXVNNoKX3u/Rc/alUkqmRwoJSshplKnn9tdz3sgUTkhb/6K
+Kfm05E6ErNnFFjj+KnrLlWUtQZZe83KTf6Bll0lYn5zbUP91FdA0nyuazCFiC5258wHRVyW2q17
Rz24kQeo2t76ost4jsUvMQUWFkQoq4lcEaK1CeFFGwXGqIDxCA0N/a96R7uMk03kknCBDAIGP74H
QJPStEDTW9gKzAeyqGo1h4nnwTiiah20vBhTZebmqXyVJ6Hg3eMhnaT+Y3xxCDbRFesNmu5ShACY
2IS5Ij4AhsxIBmfcCZ/jSm5/xXYBi8GNUZvJTnroIozt2W+ntfT26GV3t+ozTfzxmRuwcSZ70koC
FBEhumF4H/kqy6UyIgUhdFEcMGa/ttWx+73Rwmdw878FYDAY3POewUwzrBQG1Y45jLV4FTNKwfTX
SzUmbZie2Hannnxdyx+SRSTKGt06qAT//BY2uSCSCV5QnnMofXSUORbiPmuoiFn04N41GBHgucXU
jaLmVJx1Zs0PIPPm3OeySlCI8i8wSAyQKUldGN3OjfX14aN5RSGG0vBm90wA0OZRf1d1htoDM6w4
KISh8kIsVpYOI19UOJ50BwcHYTaDxw6K0FuJlA6vImDKqTZWMgQK4P84hlzAJj/DPgADyyI1BXZ+
jqGMVvHezivVweiAuG/dT+Amg0kfdg8s9HLrgGJgFPQj3B8/XxjhYzvbjRynf0dfSWoy1/2CJSrR
JtXsDIRvdblBxHkgsmaHDInqbF5rErT0YH0X/CTvVNuwU298bgQF6oB+q4Ibx1Own74YvnSgEQC+
06jYLqmd0HREScD3GABQ1lgspfNOJA6ebI4vZ0ohPb/nEE4zFjp+6R6RVDY8aJwXoNXKyXictmvG
AjLyk1iE46WfbCx/8+iAAanmXwqRmxaj7ScIkLdn/E+XQmlzpwzd8mOn0uwlxqfEvv0OPqFqdiUu
FX/7FyMJQhnpHJupbw3YqKd3DZpZmrva75OBglKzeESSQUUhEJ/2c/FdjjEYcKnkwMglNWWlejLt
stFp/RV6OiqrPtuKV5kan7spSf2w/TKV5LnCmsMUmySF/ENMFVGw/1KrB4C+myDdsy9A0H5TZJTW
ovJoV1oYuoPFF/FxS7omv4raDEwb1J5dsf1EVuyXVZCoYl5OuXtJXv+VM8+HilD8U6NEH49LN9lt
fqW7PRkk0PGp+knZlmnHfsD5M81iTl8chPQ62IE3GvIWnzLlg+qN686rCQ2nUTiUIGcOn24s1J/R
9FZmTKhgqPU6oaAEz5vCyrCg8kQogqmRBkjgspDvWmddQwJo60xG1W6i7MoDRt7oQ6cPU5vOMyQj
18SW7n3ZB2yYHK3APL/36I8qjGFyaQj3mPwYGDzYNdH4T3Bs/6sF0r1BbboxFEQ4zym8O/QcZ8co
e08hu4Z7Z7TZ5J1hliC9hDkZyVWGl+Ug7MizurVrQh+xzlssHZvLCsRTsK3LHYDVbqu9AzWwcusJ
iZrzyXdJQ7TQVriexoveWEu2j3wq97DzjOI3u2UgLLtamn30+x1Nr2q9SJnjMPnR5U5Ld0rcQIPk
zUMVtjPtwsQ1hnQHyX0aD8vNdr7ag7TO6JFBybOfig7hOWSUO4tnipGAfK69V4fbV9JWL/7FacWA
ImQElWFNYnEzGndPBZshbrpHt4cpDBDsojpjRl+oSgIxAa996sneQKy3tl6LoIuL9daWZqsDaY1N
AqNpd3O5XwS+YAjoKuOiCf1PkUgMBLuuUKBLAcS5gyG0T33qzOv5A6Islw5r0pWyE7IjkFHMZPjD
mIkoET4xSJ6Zni1XSjxbpvEn1nIeBknzbR7izSJgcdb+DWeGV2qHKhIR/qIqFQ5Zy+v1kSG9elTt
HB1YqiSisgETtAH3QQk2hLdT2wnSbnImm8tSl26Z7ISk2+1jjW4WEyg+L3nUn+TWSQYQJvA6PFHa
NZVC2Z6mq5jeIs/hrobXkz22Gxg8rdbudTOXKEpcvpFZwdCjS/wwUJpTtGypaMmBpapQE1/nWmGk
gEX88c2F4JUONMIPDM1l1aQDKFb7w+ES1DUHUAeYJY7r+DrGPRIxWU6TkisoWCkc+hPf8TiIoP17
1pEOt42hB3KaaaL6J+MXUqP2JlsljHbP6smPOjdjO7G1Q755SF/JMUr2YSX9T9NYu/E/vBnq12ba
uqNeYrPWk+CvtrcAHzsXBAuSNbg99wcK3aHU9d9b6aY4xzsulI0sAD+sfiJACxM9fqeP3rBSnNWC
/knb5p7O0fLElNmyxlQjJgcLI6we+mJ/o+MRE4oqRxAgS6TFLxQqOyHInnyMINmj3D50PIGybzmW
cBFl/XdOnsvWSUd9VB8EZg4AAz2f5Ow2uZRGnCpdgvOD8fB2ZZ4UWf6V+HUU4h/HLdmySRmoH1w4
0U5FD68QJ4WjfaVfue+u/JNrpuL+9Zii9GkCA5a8ynpwem/ccrABkYMm7UKblFi+nOSfhMJ+ygZr
YDC+pW1F4IF1UYXCWekwb3pmmfz17kgI24aSyB0y75gtVaur/Y35HMOnP8qc6567UaUf0SeRKCN9
t6Ryg9lKX26eobZeO7F5c1oc4h25DE8/dDDIOmvP8MrORlyajIauOsPEoCqrU115Wmqc9OiuyI04
mgZKSHOM9ptEZfUEg0bI9o8FCU6J4yd6JeLVvbvJa7Th1/wjbj9R+0UlLWkhomuYEdwL/aZv1P+U
+oLokhFOy+AyUN8IP2YRG/Z4LXaqPj0I0qUg7W8YwKcgDnpWQtFbX4SomcAea5Pv6aT0bvtdtb+s
hNIAxaWBX+qXQgYEh2wUjehM8C/G7zmnueHluplm30bhz/EnGccml8EnJM8cBCAAbIf4Z4/PaQ2T
IqJkdtZee/UBgjEWdtS7hJ2YM49MipFjvqV9pooIKo4kuTUt63JSH9PlPoncnYyb0/27AT8apUSc
XyHsqUjT5Hx1zj/NTVCHeb5ubbM6KveQ7sdVi7dPi9/xNPkNRSYqKBAFcLeQjM7zi191HAc+xF4S
Btvz0+zIPbMG/kCCczWD1bEsS6jWk5xZ4WE4DLRyq+GMuqff/4SmlYeFPInjaep1h5KgZsU/Csm1
zjPGXRLsJc8rYC5Hm/FuBwZZqquUpA+6vOT6eR3Ei5sAapH9SaXWRK8UptafS4wn0Irhc5/sM1N/
sK8Qu5r5a2HuB+6t3pPiUCgW7c0+0sgFdbccqtxEVFV5XXrNkIF99Gmj15ilEoiKU2lBntSizJdI
MLUEVqOXfVMzfa5YrgEbnuiYPKhw1u8ff4emi939vK0sKWJ3UQwm7ZGzvFGboXvNP9J0OeGkiSou
mFBCYjXRA6+1zI+A4wen1cWs3o0tNdGUv31qHVBv1Su5qfwHSML+HrAzn+KKhInICtxNQuVZMYwM
2nNyP9+RQnUedVXNInoFk7cGx5XMbeqRjsHWSxrciEwJXMy6uaPx5kCfKQe5dB5/rS+S8ApRTCLc
djBKO3dIhVccPr6Z9A9UQuk3W8w0Qmf/L8Gxvd5ejbuy6SxrP9/eFoeS1tOV+UMinFAcK/+r7ddw
W5rHBI6fJE8ulic1rO66C7UVmNJCYiiz5UBVc/GkwgUY1cjjhtJcZ46LVlkhC+agofuyncjQXDet
PVLczGE7Cakdi6j107mOGZRueebbc09lvgxOjo7CPUdqVSDII8jPQrPfAWWL1uHD9v9lmMxWUwQA
bBqbm+h5RMcybcSo0JC/iMI+dZYb9ym46zj4oC0+7Obg9ZOMUHhNyUC0QZ71Z5dWM1mP9U729gyr
NQS5tdwK92udCLtFocALXt9p1w9iwKNYx2VZKgKbmRjLFvRQt+vPuHa+lRCED7gU9hKNhylRZ4K9
NXRxyFIAYGYlySzvarmojkFadUb8OzarNu5L90fdm510iOhOHot8m7F/T9VWB6UnJCusx/zX9pm9
r+5IwpjL+HYQr1o9VVbRPtYBy8EXFr8aHPtEF9q1TzjGRJJnEGHDtGx5ZTRsE/h3Qbq+HoziUHPw
w7JATly/Uj9GcCMuqhVLxo6wA9GRZeIR67Zx46SjpLIcD6+AlyyuvVnEz8j7AB3Mw5ZfwUUU2pbi
12vnxk3zcWHu39ARqJomH9LxRdyeDtZd0BxoHbY51eiVtv6yvE4l+pi5NdeQqlkOUS52FDW1+pFf
QiuaFNxrL8PnB73TQtSw2OSSjm8FYSpwrDPlimzEDOcvlpIk4jUe2eo1F6l0my7LnmwtJUa1V4dg
NJ45nAQGss/PRuI5lj358jcJYJGojY5R/nhu7utw4EHVjp4Lr1qXgvAP5GB5i/EA9WWghtzQwah4
ZimiZDZ88Ki+NhGLE/QuLv7bFkd0EjCVafzXeCgDZjGg0DM/lg7Wbn/ExKLh/4EuNMyaFGk1EwbM
bBZWRnukHbo03X3NW/UQyFvUBEtv5Lfqlszk/TDfldozkiJV5OpBFki6hLCp2DtEcyaZphtj0w50
v18gdKRZorSZSw6VPrQcMRTw/32YUZOkKKg2WQoIDnZR8jNDti/6JSaiOEPTOSYA3N6fNYHiXzhe
1xJlKNvSA3lv24QBp3/OLyY+Pf6A9r2DCqXZIjCsMuOwLerqtQjdqlEGX/2KXMB61eiDiXTs3vyx
nsy8l+FxkygkwMLU7mAZkeusvhbTVDameFiZMI8ZqxD0Tk1QSn9Qoim3YcWM52sNlUUFXLQxF8yD
jl3E5sTZ0E2TSadG9OlsjYD1EeEOqBMMFMQBSsmq79W4nU/OxBeDBIY6WagevrQTts+fNCh/nFDr
Qnjvp6sGAW24pMS4zEfINn7bfjRV8YzX9sBe3wBCViAxJGaVf/hRACeUrbCS97urouPvsIkpdftu
JuRl0a/LQDnwEOPNDE3QiGNsDFMlCsFW2DS+sy4XrLtvkEh5iaTouNhShWLCFHtFjH3McU2SZA3X
bS2ts7JeCSX4jcBoUCC+mg5QOawqLf316Apz5VqF4BTAecWy+pq5lalsgIDdQlPoVutvuIQM518Y
UWeJEozpoNKK6sqjoaVG3P5UXPFSHRRsudP3LAg09nNVkyvmKdCtAJFRFykUcxAbJuGljNhv7zPd
x1ni4QhrNbxfZ6eKq0hdQpudcRpeARVVafW7OyiYiN50a52iOZvxChKihlzgHGSm4+7mO7RDAuJd
ZVObrRigF+CZb+K12rkjBpleRJYQ0PCpdMK6vkM2Zxz9elEK2cMyH6zADN1WRsp9rjQuqMh6jpKe
2WevWeNeNS7OO2yZRm7NqCbeRWbswvwQcwHyZWfRJxS0KIy8IkDC3aGbbLv5URNHve+OrzJ+uxUa
ras/2EzAQnUiDyzdopJPhJuJEwufo2iEYcNIf3Ntr4PzmyP9KeDkxdV2hmzCM6if2wJa/WR0UFHA
OmMDJdyf7cLo9L6tI/+pbG4wFEWKCGmiDn/pBQKQAdhP6DJQcIKnQihmRkU1A3XqfPVpeIKkUoL6
+g5BPhY7aPh9fPE0X4LmzKkNeyeRlmUMJPSBZ5HEuuWOWuFEDNlfLGblfYeYr2qR0wccUUDbW8d3
h4zAkFmGT3cY6oU2IicJF5w6Pu8dlpR7Dn7OS6OdcB3rorr159jiP4GX422cIQ6NKgmjVnbHlStj
nDBo6FE2V0zM4n0HX2siKFbr9ii2oUwRw3gFkwZeHXXH52FD+HLc/JzkVGHAbO8JjDuE0qTZ6cxO
w47BAx98CSEasfVGjI2P9Cy/m8QjNnFeqFl4mVOvA7gWJ06T2gMrFF6tCeV5W2c2QRn6wlsQhCdx
PSI9iXlTFVctAZSw2bw7sQqTDIpGk2ivBEbSIWS4ttKmIUKf90HeX0brbyy2W22wP60gsJlh4kHm
X7+WySkS0J8YnzwXLUw4FppRcXAgiio0W5FmKXp8sDRveqNuYgg9+S8cabVCcJ+Vh/PUtuDIYyNM
hA334suEooCL15cEWHFCg1T7hXAbXY5REBXUhV4ZEV+aGDqh9JpoSQBbamE5qYHoE264KDMW4Ytd
ilSbXeUakwnDAPf9jBderrVQMK5PzsudqY5h7OJa5Rceb95MGSzTEh7zCjIZWcJpMwipq9QPxdNi
0nbQ56NMHGYg2iK0L0cfKuDm5pnbL4p7SVZs+lbxgENsP4gXxiEhS+A1sXuj/77dXv//b5DoY6UQ
Pv+ucaG3uQEswdmGeGJYBxoAd50UimGB1x2/Q1kjiDsnVnS615K8JZpHvQB4iWPE3MnlC7ORiEJh
lkPyw3TFCHWpe+yRWVpqRQRJ0ej/bX33Q+U/2Pou+G7sqP6SACAIwGJP8AozQRZFKZzC6wESz9w9
2oKWe6CQi7RTh1Mah7foRA9TXDddyloqsODoBK6RtiGd/HQ1OKVwnePio8cJ9WVRXFD/9zNE01LU
mba2aG3qt+oQriOYmgZGLzrR8l8Xjb9kvskE+gboc6u8PZFy3zdjcfIUfhODaghCqlajjYMcqVzy
jww8Wh4IZ2na7PuxK8jKdhAvocnJf+1wKeRm2+cxjYncmHGiAw4nweBEcQEBBm37XxQl3Flbdoly
HoM+rt6hDfm8Tqv1HGNqlqTw6t7JgcQ5CpkmBqvb4LWnvyq0/JoegWuFt3Q2/jSGnAewcUsNPE9T
PBQY/iJZfXE9WUDS1JZyAsPhcvMeqWtySyrIDPMG/fViueKFtw5kL0cW+OjYOZvYNwH+z8TDb/If
nU+30cs/ViRfSD7k9otlJ/VSPA52rHZv7VoAeLTvbAC/os52xlOyPGXAGm3nsdeJbw+JwuPpU64f
Nddbi0hsgpJchWM/jCdMQlC8yHQumw7CSo3V6Fg4o9B+RCj4yUwqmk+IWBTNWoBvQT3veLBF0a3O
AgEAZsFCXZAJehp+ztUfYVeEj8sk3BCKoMruOQVxpVEEDQoMifRTY0UiFMNUP7alpzmBXjYclFog
de1qONNjkYpc52nHTmLP+6R3jXkGSqJvhMXOip0hgT9rjtWJhT9wKKTVH65YXzOwch5Ef8c5SIY7
tPH3D8ixbjNQk2pHRmXcOffqkECwInl7y3CC1O9jL26nHNw2JtPfEaTMFgWhzTk1e5wABZzlldwY
msWgawvHpPWHSI4oSZlZI5HNfMSnfGHpTeZZjVCuF7p5aG2zK3XLka69IJUijxYpBPFTBaY3PhKp
GM7KdVyeUEP4LuZXY7ey8BOjh7lLdVlTf0/d3EnRY0mPYTROJxcW9HzRre5pPytNenI3idBE18Bc
7e4KJktw0TKEn/GjwmuBJ5Th42U2hFJFL6b9xGu7capLIjTv/HS6xN2tuiN7FRQw1pyk6VY+QJf3
UcY5JRUpLf+5NecIapuLaONXiB7uU8t+c4DoqQV5MBkOmzC3m6TZrDa7174rDQmo+cW1Jfx09A10
ortQkdwFLa1xp6sxmUnv0LbG0iF1Pk5N8qGusU44mp+aA+EH3SBg2TqUNDdJFShMeOHHJfwSjqkQ
hhcOkrTkKbllOHNhcVphFd2jcabstye3ZwSJmG5Y1lDFLKkb5GPsNxICxn6p1OmjLYne8xBPJIBW
aR9JP7jr3b3RYOtmowXFtENtSHa7hIFn9rYjlsPyDEQ8hznlj/4gSxwdVMLVbZWlWiGt8irCAFUH
JrPUdzVaHSwN1Miswc6lhR+RarIEmG4M3EK6+fg173/VScHiza4070y36gvjl/n/0bTQceOQ8XVZ
5vaXvHEPyg5mEGp36Q3E1npUZCRlx4RVqxio2k8kjmbGmB8AnLStJvodr2GnMPYv42hUyYzTWJk5
MM4AxW0pHZm0H9s2ekJQGciLm5iFkjPqOv5Ooc4+2Ew+sG6fVu4UXtu65Y6Y5j78xBBJSwJJWr8n
OBgq515wOO0a9YJJssIqjN6BDW11b7ygKd8UmjYdh35rpDEYjEUdDNaYliwAG21Zl6DDzvlvozpD
X2iqadcoU5OCdf2AHXL5UlIcZ0hQyRm2nE9nD+7lCh0sbLaVlyt427ygXuun0F6JS7W59RFLhQot
DMlFyeY6LiH+Q18yl27qkubyCFTjEttkhQoOM4Uc208pfxhP1uYQXS/EB8KrbvTX50JMackOBsBu
YUcya7Teg7Cu2xqw0+a/Fb1mxmf/ssdhhEfKIlS9VW0bUZJjypAJj6X+NeIKbYvBiThp+V71Q19b
499j9IPqV0yrEGBTwt2Ej9W+zKJXxGMrBjESuRIUp4bywC7zOowiTT85NsllMAz63aAlcRk2FRJF
VCQzndhDvJHYRIXzEPEgNJD3BPLdj15vyvGG8OtUyTPKPSY2fo2eoeSHiwCD4vgjzsDM0sRHPJ9e
4IW7aw1KolBteuvz0fkADaOj+r9o8+U8MevF15MxeULOoNdmX74s02rKf0Odvg//XhRMkI7j4040
vpBfCbh/XU/8ERw0kp3MoHPblHUBc+xzShHGsEWjJt9bdk79yXo3DfDWyGP8WcTL/sux+O5JBvIz
a5ujKPAKFxqTQwoXVlw0gDwwipMhTUsvKtXq2gnfePJaZKYZJGUu+Oes/Sej1QQ8MEXCBW0f1o4W
oScFPv8bIkdT/YXAvXWfSroAhrRbmdges8UtnILaAy2rxv5KydClFACDfcdrc7jgJdP3ecm+rBL8
quWSPhebmohJgV52rU+yO8amqJt+6tS1AHIL3waaOJQpFYoa/bbxeF+GSg35j1oFMliVTE4I32NN
YWOfKebtk0StY4ZxZIYicys6cXvPltt3obIpkGu0cWQKhHPUkHxSp0da8W5XJkiAk+dK/9TgjhLX
cUj9SKFUW70ie02YXDNLwLBeJ+N0nY0VL1BueigDkfvhl589kuQgiTDgcrJkeAtDW5e8YZePDt3j
K8rK5qSedbdejDCC9SHTxjm9nnnLrQlrVMq7UPmGGSApfwSIo2S/hIRzeHDlOQCoeFI6TFHkxg2D
HVjY1TnbijxyFsNrZUYteAW1/Xrgk9/7fr1eIqataSuv+iN9+16j/yQDnBqNicvTYYvlbYQwJAOR
MfVJtuVZjcbdYLJ0GNL3h1Oij1CwCgAyvmzhJnJFTCZz0cJGmboeaZLcTDaScfij+1GfMLW8vsWk
pctgSdedf4OEtBxIc8esiQQ63xMUGspU/wyT/q1PDQTkyoUpZTcFMFPIZ+YAiYtjB/IhLpJXJ42I
XK9aioz2F1SJWqai21b8OynOu+aGFtXmbVIyZdw8Hxoh+b7IyDB+HRKEvp8olCsHor9eO3gAlw9P
9/FffbpBPyndkWvScYnm7I3zSoMCs1ZMRS6xuBTlu4uGWujqM9dpG2KAlLin1CC/TuJqogKjXgzy
E+MBc9LLcTauV58hMfqfyFYaLkZsl3YoQ0nRmo7+6cwovaYH6+YZw2bcHc2GtOmTlPPY9J5JBTUs
8yeOsdhGhZ+CKHBLvhf5pG3j2pQfhAF0Ln1zdLqWW8FAS/X7Jh+v5eC5zwWw0DOgLl5RqlnzZGzN
+13Hs1uE6iHTEfe+Gm9b7nJ/eD4rtnHTDC/PwOKi387ZMH/4OpQ+0RXYsvTkMz/xEDqSQa3MIAoM
/DFP9YhTvur0RA5IBWbM9igqFLSA2S0RYqr2PaI1uNsCjoZpO9DTmg4VX2rtS8GPaE4hpjkjvrVQ
/LQ9nmutrJzhf1XaPKF/JtqmUIbLLTaXs/11gv+rTO/03LAQMoWuWJM38mkCtQsHDBk38Lmd1XxI
dP0SygKvZaGn1ZG/moO4ljF9Oy719xfigBzKdLT8V3auVvpdj4HzrLvzXvGwCuWgP23mmF2H3LCT
PH9ZO5+hIaid/t8TngkNp2OAeIiTkxALjhri5vvGtn+foRx+fZgI8AUzmXxVff1oOj74zM0Ri69p
DGcK9rL4aUEUV48E+XG6vFyjFAvEPooG7mx9+6Xonxm5ti8wY69UVx/otedWwMY8LxvO4lmEqCF5
7C54rBNpc3Bq0EGNY4T2yHSL8TSYtXlKQzx5KzSJr/LxYvTk1Ib/E2+YPzfQc7e132TEQkum0jBv
oDjWVdMHnSBc934LnfftQi5mBVbPB9J8i1MAHZRiV06Vv+r1R/DuyNZU4HNBiiwMqCI2Wjs+Ydku
xvV0m/heCEit6Y23TwoP7iO5nFl6g2z85vVwLY9JliNqCNE1wn802ULQTFObihZjQCs4wTRUgvCD
sH0r0zTSOFcCxjee+CHvKd+7y4pTgKbhz5O9x4A3z9ar2+HftYkie5C6WsKXJbHVgl+Yp+3eY5HS
tEwV7TAgDohUO2pMa1aGkK0cTXwDNdKGsLh2n6O+6jiAElKSkbdF8pidxOyorK4SLCZxDgosYdxm
9GKja4xlTc5JXIsBNbl3hhRW40QAu0Zp5RefP6J3wWJ6jJQBBoYrCZcysW3Bux4sbMKzv0l9//Gc
QgS51JowZhoCFbgEawSI8Sf8AtHUvvnl7jCUhHc4OPXBzyUoQyZPXY72u0WGB0hPuoL4KY8VUrn8
N66g4CgvmwRBJT/5Gv5ssa1xOqbU6HSuKfE12HRL4I+0vllod54C30fE0j5hZfpV0qK80olBfz8e
CzAUEdzNBqHj1+zHeQeEFd7zAOnlGbXTjMxX/Tx5SohNdseU9LIAfwAleAUBm1ekmzvDhEvKScwr
u5cbvML/diupgiG0a3VnolUQXlB73bysBnuBuNtXBBKNxmxFA3bhjSu2/BSb6EG81eFt1nQVzcmt
/BmuN/I/oE8kCxSqZ0N/tdhP/biODBHOdT21PhcTPU+ysD8DGtJZ4tEA8H33DPrzmxTjBDHXICtM
Z5WFDErUiPYYV8CZs9cIpUbTkEUFCl3rOYAHkbzZyZvmbTADloWhtYDjExnK4rRaSjFANW23N9QP
vdloQXbc6lHoKczmtIb9CFxBJQ4eiwPHkJ/pkAx5cbkI3JdnQoKymyDNjuw4h3wvfmtIb+y/s+Yw
1Lun8iWxpebqsJxbaVpCJRRucvNjhtbNzqv5OBqdej174Y5SxjNmq+FP3vTqDzuV75REBvr6Y3kf
ibtrqG1yP4Q4G3h3snuI4pcf2M9wXXH9XTJ/e2+7HVRclBRRi5FngImOmobuUeMVZqKSbm/jwL4J
gDBfuEDuJwPo0GAC8hy4Vd5Bb8PpgXLjbJ6vXbvK6J0CLJXAM34gWzPycb+vvPdbtPuxa4XHyJt3
oYelF9Wx9QXVL3vxjmYP/k48DBIchoLqtkzJpkgjJJhX53qqaaMeNBnfiG2POhEGww7OrHtwPGUO
dCpwxOfCqZX7XB7rPsgsWM3/hKdpMfextT6XFEGMD5eUxAcJBUzZt+ngs/6MpKU++GaeGBLMfPDZ
Rug6X2e9cVU4h5IK//FshJbF7b91XbggYEX6E0VBNgl6FhA/O5FncfoNADYBHwCKVA1+Z3MWoK0M
CIo3adp8JunwZ2soCRnr36s0OXSQTXkkydwmONUG1n33/ITCcjcsQHuY6b2KeiXUkIPNzCp+0+1S
lzXFildWXAOOxju+vlLr97AqqkCpb2QIzaI6GIyaAkGeA4d0yQjc4Wn/e344ReZIDNbCzz/xeLS7
VqopBDDJg0RQK65mdm3MqAXMcNWewXMK5+mw+GOJn1zLcRF8BpaZzCHq0Ycm2TOo5RBmXPNnHn53
DdzszGaztEKNsns3AGgXLFxMxJDQyYpr3XxRDlJ8GCGsG5Gg4qnA3UNLKSdVmxCN6yDvcN+P6WEm
+etsCpK6364YnJvVp8C/sUm8fMdw9Hm844tPVV6SWFaBO2aG3sYPO3Czr0O7hLTx3YqPaGyHiIRy
Kd8Gr8DhedtOFZMfTU80o+KITGBPL8eB0bhgVNPSGAchxrxjuWGz1Z9r7WwCS02SrREqvHrbakj2
xb9sqhab51Z/072fNR7Ejr4aQYk5xH7qp2TgshublHhMlCA8i6kcQ5zzIJjrTnudaohOThV9fvKF
T+3odbd9WYRRjDPPoJwiwrLr1/ssPjBuytOrOONQR6fsscf7MKuXUT9axyrtXufD66fhWPJ5YJ84
V1dSPKYe75x3f9GMZ/kF5H2G1YJodwfa61kxPTB5lulGFMAeXWq5afRiBaeHF4SNVEy/ov26jpMc
gfJBlG8aZDY2ygl77F9BnAqJTyiXXgS5FZLKUuos3dga3MjxETKEWL3LW5V8Xqe+c7OIyGKDRSuH
sgeCiG1rML8htPVjh/jugB8q+LE90rrK6TWAVM5KyLErlmT+bhXWJgXs+sFkswfR+Ra3oUWQ0bJe
XBLEX2Jw8kFLlBuRPOcE/SVnhO+uy3tha/Aq2IafEdV7gXRw1VOOqutXYry5FOGcRwUmEwcq1IRg
OdD8r1Vc0AzCXF7B3To8zX/XF/5sKxynfpol5Q31LdgatC9jBn/RPC1X36+hWMjaVW1eRF3g5VoG
2PjXnYDJiKWQ7pT0pdNq9L4iO0a1XSz/g2O4dIjeAAv7zm+Hjxt8VOMQfjK53uUgQ8pAxvGt3ImL
oPNlLZUjSyndpUBKboLslPHuvzG4XMTpsoQClqkXuoOuX/48rgfaVlXIVyiIXn691IYDUfsnaRZ3
SH8h0a7HnylqJNl+17znFyB57m9/NPGoq3bxVdgt1c5RqTOjfKFh4W7bTXnVoM57Hk1nmzpQtqa8
dSRUGeiSzxi/jWyHkiud4PBLrvEtKVVfFGcMf3327d24P/ryKvrq18cfhi7pqHfpIWDsX+WzrzlJ
a7zuguNJMKPyOt6TLd6XKwjLG59Kk6pHCsBAVOcXOKK74Y8UDi8P7PudGey1KJ9He+DCyLaBJn1t
ZYgqu/KMBxRnULGMhwTLe22bEMb1jiCz7c/FEg6/hRMHfkZWbmwvwjNCYYj/iuaHziv/GVLYeV5I
2p1tW4Wbqk8zJO00UAn2ICvlCc18tkx1FzfszSl86aDiQivPSvh588osNelPhiiktIyOcsrQU71k
pF6algM1iWe94nAi7V7pKyIlsUBQuSNk/Tozwvp7nxe67l97+3Ij4EKcl6DwNC1WJLWbE3bVvdPf
pbbjnqPsNa1v+EA/7Rm71AM1lVzh3QPDqXtHI0b58aVrWr3r3kJHeIINThVD5iwaiuJ7EKJGxWAM
0UFmYmnCrz5MNAV+CF08VlGy8cn8WO5iX5kwz/dZtuHcCqPHhiTg89JnK/HoI7wnvjxEUMNa+pAQ
2aa/WZQdveXZu8JfSV4oMO2YvYcSF+R0qiG3b409tN88r0cshdtxl9IuHpovOA98j2LSsWI+hv2b
isS6Dk1dmH4ZN3duagh6cd+O2bFY1k/ho+5sNwobJ+bUYKCV9Ed5EDKwx7Jw2Qapof3t3vDHQWdC
dDgwK/oXzYZ+wM/ynLl6+lho2+Z0QoxEVziBBVZrHRClJvtQOFX2V1RVZ3AT4xUj9cK0QVEgEP+K
5A/oKeZpNOKSUByL7OOQ8wozSFVcdFPDkwh42EN/RPVBGJXLvNebSYQJp69GWvrzSnGW0vnaiTWd
I7AhGYgTs41IqJ7V5CCVnVylzE1ilFb7t+qxoyrggL3q9Ou60ZePoMxC5RLYzvwPvdazS3AVMpgy
iJcb471LkekufAqTDZnxQh8pAYTMcsO1jR3QIgj5x2XjKlBNU+1isB8PbQAWWBjKj/6gvgV0wBWZ
prX0ZK4O/gp/BeS8uFlDzzKvKU/TLSZDXR5TjoJCHTwcs2gWjinvOLCBexIKhHrXIIxU8Rhq0ekC
e+BXHHtDraA3wha0ZQVWQqgKAIb11DaNRKeTlakFbSva+94kVFTEfWvrx1hcyWP2ZEk5gONyyAQO
6ZHvGBrfV++DCfkwO/Ouy6oKgZJhJ0odytHJjdc1/L8bD9nNYHAWOD12rJe5Ef2OZJ+Xamd1VlH7
Neh+h0+NPW2gi1FYyOcOD+kKfplslk6hkkYX8c6ggcWbfv+ZcM+Jrn1dme6tXrTDuljHzVCsP3uc
/YnYZMNEZYH7Qu/kbUjkCOBQ7XiiJO3FjtHIzbrFT+pXWTP5GykFqwqgB9+cMFKgbOdBBg5l5mly
lgibwR6b+o0199CSj068+TNd54dn6cWHTJysUvdHpg0stptemqCrC9TfITUs6p2ox+uk6HnBxqaq
0JqWQgWWSDGIf2LU6md9BtDB6uB3AyhtLciPoevyZDbct6EXkJwr3aLgsifEJSVl2tK1N6VG8RqA
RiF8W9XE91Kd/TNJwafYkIqNhl0IKBr+7UJ3P82IAYQu+/i0TFYCLxyocj3iQArWY4TENHQwOINn
nBK7CVFWvaeeBMKwWSOMG3XfQHhmXt22p/pTdngcf/D5T0pypbjltYFEc0ak6xa7sbLbQi5NF7P4
CAXKKRZ8atvBwcGKAzp5+NWlOj0G+zsp2lNxWuTJtktaBcDCvWGsMAlM8X+WFLHKBmtV2Em65HIG
zAiufxkaefIL0iQjW+j+AEb/B9KzAISoEzATWaiWPViLcm0r2FpGRJVmKDj3gaBo28GWNi4+4FUe
ZZlOtFXz5MbFNs6BcshRELHF9sLjpVwLsSqi9QmgzD4+lyo3sDxZGTrAZ3VJOc5rvLMSYR3CD00I
UNiRUDEZIBjKlm+meRghzlU8hSmfU2h13c9Lpd2fL5f/96pdwV1zSZMrJ5VI486I1+RN3FEqW3Ea
T5GgQ+TL1QQsf4zYF2xH4rYmdu3NL/HZB8i1lRHJvdYyTnzCjTkGvVDL4Csqr/Oj8KeX5iGZSzeC
qB86ACzS7giaDOGCwhd1BovrCWVdyobGIe+A27KSn3Tj5uVsGcA7GovoeCTv3shwRSqhyOP8Bou6
iSN3jk6OTIssMSveLRf4UYdPOpPF4yfNkDappMQMrNKg+WC+/KSS0dWi2lBVR2BMtnaKSD2jRxVB
GlJgsGIO52VOPLSbo+E/6GuLfPj063VzWafr8EK6L9ufMldjKuqSXQ3hNjA5WXps0hOlsG4Y0nQS
ErP4jaDM7+jSnOxxAEY+yd8EnHkjpSDx1roO5sJ0JkZhvVu/LZprF77oikOman1228nT3BkjsWSP
cyH8kHTJm+fwblx984OQkW0RVj+1s9JqB8xkAGopSNGnyTDO4t7LE4VJ1zp/dagJwpkFM0SgmJbL
sdQYn6RrCNZfYHltgE+ypmYvbW9iTBRyVySVV5qjRpAm8jA+Wpudto4P4s7HgayTDeJF/0obuNqv
uRf10F+8jPEDdqCbMkhBFTIG/4Y1nVIAr90YZDgAN8KaSP/wD+323OVla0LfxgEGXpl9JjRTx8Nl
/IBsppjSQHKfwCdPCZFvKTvskZ+fi2etOQKN2sC0QdyhUYImoZjMy/ZadS5KjA6ad+ylEGzeOvIr
EzDXjWBBx50lF7cPjBKiiPPnqUTrevJ23a2pkrW1LtfvJEh4KJfFV/BsPNDo4mbfgZKf/wqmtIOx
18Z/8dAHWCb70xgiTBwJTOU0z9OdRUJJwbUpSlbi+D/8ktE9oSIxDXrmAWJTuSDjSRjzBXago2UG
Oor4qOZ3zBhKLPP4mexf6qyatIrp5zFcJ8Tk9ARQrBnOFKyjY84xTVShVFkpHSif1LO2PNjDdYQp
P0HZR1jr0OM8DL7huG7ty0z8SHh03SMw0DdtsmgLWFddZkSNHBcbPzqNywZlCCt9nu59V1PCOQ+s
fAiwEI3RuMe8C+fhF9/LL789uCNVNrxkaEjTRPTNABrlwjqL3YzOWxAYmHg4vTf/dteUZyqgxd5Y
v6ZwPhgayUqOk77iv9D1is/xxA0D3L5lPwQUBhoU0AWB2E6ZptZ6vpJE10SGAIz/8lmcWAJ7BB3r
r1ZdWY5SASOKHSZXZcG1Y8zq/Y2ebYAlePRZem8NpoL9w6/issgEeRt5y5kjubFmYi0Xe6+U3sxz
cloZGA8VWRtCc9cUfRsInp3LXcLHDMVh/RThvTnpUhDWpBmHUwTnm+I35lwv6ECI+CfrH/+X0rmg
uddPZ/DJBoxAfnGbn833EKWYhmGeZrAI9K/MHrkrJGCQJtybXOMXq8QPszXvcdtxZV/M/m9MJJIZ
kwmSmvfKswe4wPyt5HU5A6DLRaYy8857qr5Cvz2cFocuUgCkGHsP2t1nVnPmkD0LC1Jqj+C6XLlg
H9RJKZ4IJxfZBdT8tk0KeauuKlE1MQ8vEqcwgYFUBUqrpIFdW8tOb/NMSMDOym47XswmNB1ytmBi
DPqVFokLLjfQRubECtUSk0T4WVU0bo/xdz3VBxwDAAl7APOEPSIsRQkc4ndivAC4jBF88FIcnG1k
nPSsKC5/bYLbMOOfVyiMrhb/zwAHUa+k2yjcgjKE8vGEuIkebznyItMoEV/U8R/IYE8VOLYD2K90
XBzLR0p6IwCMBSIDoCo+wBaCA8psgx2eRd91c1l9SgVvA4O69X8f0lN9i2eMFa5g8epoMXX7Z8sJ
Q8wn0wyhKUgbH3Bp/RuNnL6fzHJKvKpVYQh0KTq/AkmrFwh+rTtqpA2lH2DLGklZ11aMlHc0euAD
Yiep3+NS20uGydZx5h0JnhpVXqQWp9XBXVFN7S0lBYrpcUL2MApngPHd8MeH9p58Dn4zPPtU0Bcn
bf44cKLurI5ECfEa/LJw4ir5ua+9J8UEmLLfNVff4304PoZ3fc+lFPw7wCs6R1faFLUMeJ7mKYKP
+AmhcT2e5qkh12KWIYFBLx+au5mVc1xgISIa7VuIUX8TMSji8bSQ8yvH1LHYGGN4XcXkwzwGgKP5
ZtjXb+eDBHIzfs50A7jYRJISrTnp7jwmvGDLyutZjMGj/k/Ji4ktzTQnYAdhXjJoDJsEFqfZgfOJ
kjYM+Zs9lMDKvGTcMEsqLpTrA1fqrhToCuHJYFOWE95G3ttUyc3Mx5NM/JzHJ/MV1QvDzGNokdaR
S/2PvcbKwXvoEEhw+3ddZhs0/DLHdE7MNMGT1bhm+IjgISt57+NblKrzN9H8FfS8fYekugOQgwbP
x05vDU4oP0wC2XSjA6xCIr0WLUun7uXboaAHDQIsZhGIrAJVaSttnYlCIXtop5fBsqwsfLZzHNhS
DPJYRXsLlibqiXewdD39evVbBtqpOAyEyKgvGbwhbzJ6dwvZWq5cnz56j5N2x0LnUR7QoPVfdcpZ
ITjXBbMTAQPgtGXDxdjZQJtVERnTwaDbU4ygE2iQ1E2pQnDh77mq8s6mvNqhqaeQWpyDAJ3kURx3
tdU9vkXh0Rv7ApW5vAkgmK22ScKnusOpwFA59d5vIp3JEmKJf6r58kPBzqK0/2gQPRkV31fzcQIY
z2muhqPuNqmdK87/O5oo1Ukz+y9CY5u5yk4BdF6CJvvQzqIgWQAPfjpp7WtIfokyV2pCLBn7fikb
B1OVz10DpcqoQ3MsXQ1BdSs7uDZROMOt7jwfRZAwTdrXchgr1ZQ9xnNGG0mHZsKOaAMWzkvpJCkS
dWGNsp9DYqIF+ZY6LElcwh/J1/nWxlWBLbqnU+adzOE/BE5tzDPZ30xu+c4cZvQWHt6YwXD3Y3Y4
jaiinTu5hn1k2Da7XhN2tgRiBis+g3aYenbi4pnIJiQSb4FbsuxLj4XP1KqR5oGiO8tDGAOwY0O2
Elao4xV3zziOcgnTkK7rwFcEBT5rbXGwUbK+mvfLJVIRIUqP5Cty85Q7/48wMmqGKmbGHMqTeeF/
9FcVnhTm7lnXLeBdd85hAmCEQLB1wj7cJs+TIMBqQKS1hjDwxzxtRuK4awSV3TJIQcIXiHVZV5JP
brYunYBOobxhmqGK6Ij/3gQC6qnidOkH73cmTRDn8mTCCJxtr1RzGWV78O2KVd/gMElFNwyLiWhh
USAFM0qkZjrhz0LFVlaXWUhHwBhX4jI7ajNEvl7xslb9YjyZSwJb7rzG89vf/QLV/nGMKgEINdfG
f+iwAb8BoNr73BVfyn7rL+FPB09qp2fMgK1Kxj4q6OAOYYD/eAthH1kgnrBYu0gYZeu9QGgZnu/y
cuUYq3HrijoNYXWWjYGGgb1uGrwx94Z+uGAealF0J5x9RZWSfnuLtXHbjjxRZPaYpylw3cDDinv5
Bh4BBRp9cDQ9rjmvAVSskIhWlHrYnTIiblYSai+6Q3zAfjndu9Ychm9dR/RQwoLoaGgXjR3XqDGV
xjRwo120O/bredYLpr1ABJRifs+fvyfh9Ts6y1ox+wBLDDUTjJ0H/ANQgoMw8gmfI93kJAPSn66L
cnmhJLx8clrTTnGFqbY2TxO0hvgVbfcn54BEcXGkqALO1YyS9IL7xOC04ubeEWW5qnAwP/Wik0a5
lFT9GD2Snj6+dd5ypchad9CvuVvObagKqiPrlzvDzA9w9AD2uzFEGfZJN0AIY6hjcpTKQRf9IutT
QganQxkY668n5pGNKUswhBAUFuED9OZ1N6TiJNaUEDL3vUzDkRnCaMd/gqeKMNdvfgwkO1n9jnXa
Nn3DBAku6jZ2dvgDUDQSBT0+n8FFhuttZwuohewxke0cPk5dv4epMbMOQ/XitRO2074n9oHANTEu
PXxNsacNEgw9h+3s41syCAucRexCwlvfy7nTEYUDqnujzsmlXXcH1ae4J+FMzHLsrEL06j2kd1ko
vOCTHtXkweKr12HmcQVppBsSXyao7SoA4ecCUBPW260MFNELfmO/PeXOkSscBmHw5HYTNVWZjirp
aV9fDdsirHirkq6NcDA950Gry6+f1i768HlvyrkNOVbzUF9xaNOZvExJ6vlNq16eW4RZ9p8z6kjp
J6RmgJT9KPU9Db97QrLVXXEYZ2+wzfkbMktnjnFS0kyP3yGtJCNy3NmHhch21vSOaHdmPIhQAcii
y3REpy6YhcpPNyNC1EGT8aAAmrMp14h/yadjR8MwkJwaZMRc3i/G14TBeqlOkVy184g2d7viqODK
lqRsg9lPkTGXSeA/DJdzM+ndkGOB028uxws0DmefX3UgUbnpP+i8T0Ca/s6rjfcGbH3EcglbldwC
zKlGkUGHctZfYgo1lFxNSSLWWCMmUrXq1vcDfC91J800+oRYO9zo7KH2XFWaGH0gkKuQxOkT1eIU
HXhkUD2hmxEGuhJH9NvTsOF1+/5xZI8mZP+Ibkgf0+d4Z7Lt2mw3fswnJwdc07BQoQwwlxkgvXZk
dbeLKjjxaJ9ZxLVZ432sb2iahNKEMz3BhLbSwSaqKb3jN7k3tgl4t2q6YwKsTaccWQRCrd48fz4t
gb8PXZV1F2Bk72Bq811YY+xKqfqnshD3yfgy7cNr/4uq63uC0L63CjG+Wb+19ErQbqauxaGds+AV
u5AanHkzeoUUeZTmy5jA0HTNHsIyJSNGCwRcBl6pX7qvq1Tr40CIOnZvO6tKLqSs0dCJb1/oJcIG
fS3d4F4M8osu7zbzRIy40fInyTEWz9+B+uiClYR9dFmYUW9nAt4LehC+FeN4P1LAfGfm1tGrYAsB
BsSPOxobQvcJLcbUHr+3URN0s+h5celSfs+KunblbUgvoTLXksy606AW4+qhq9RbRk4qen/pI1Wo
6BJclNeCaH3LYdyHzIMZwZcOV4egfRtLfk1NNa82gN2jjs2GojjYPXVzaKd+BxtpwUI3tYBCsD6h
BAvdPsDayMbdmBSSQ4k7ORnri1T4VrQcxa6TH3xzOHkH9wAbBEquhBbHOiaBxFHpVaonlmKva5NP
83KlJ+ympsWvm3Uy205NAkZbyiTNu+dGkzfsDqZcEVmXiyT/Ij3bvxQo45irYG6B5OitpzvCt6t3
7HaHVZiF54cN2m8INqFmS9uvBtIRDdTDMXgpe+QocsdIjLsgrQomDeEwvjKxl5TSn1ejMYZ1HQ6i
3caXuZvSX7b6ObNCLvE5ZKV2pgcRFjObSThahuWCscW0rJ+oPUwyr4tPKXGEy1qJPrLYfriPXOrd
BhfMpk3qYGqOZVC4FkBYCQA+LUB952g7ZAWgEWLbWKAl1QDu3Jh35erKGJeLdJxIwqwyqkMOaH4V
Ce5VwkxEP15UY+N15dY5AmaTIxHxssVEFpCwke7PqSWp1T2rMssAxudFn9BkdfR6AHO17OBLzxuB
w9YcV/6rZhi3eMLGz6KdiL4AblRiKv7IUgTcBVzQU5VMbC73NE7eGOXTN5EcTBmDbKanmTuGLOeL
twudTIgrk8Xi1i0Ud06jf/qJOyc0L3yfUf4NnQUP/ylXbp1HIDE9BoBIu9qvz+I1hbTcCInqvjow
tgG/a4gUVgBJwvYWhW3Z0yHvtqKDUHFWLJOLeZ+oeX+11GlwA7CismSpzlRJ16Y1mqoe5UD4ByH9
hAwkBLe8zDjQogH0vRfIk4/NW7lCEDPk/v9HnNmJCSOMXuHjD1++dpogD8sqtoSAToSchsordKq2
v9mNdmwmK2SFBZZnpUP8SGEaVGvntJHG16oOtiByP/OufFf4de9eTuXtWyV5s5sMjP8h38hrb/kJ
wCXm2JJMCPBN4iF0I6iBAyKGdwgqD2IUkD27b+c6TQBZJ+MT5s8/KvRZbIx3XxVYKU0tZ8xUFb58
XXaoCNgDEfMboumeG8aOfls2QKPb0tcsIQeuzHmws9yOaIldu4NpqoQZZY1UFCYi8zzOP8T/T37N
kwyj9ShucVkreDNJz0R2gDoyqOgxeZX2xt7y59EX9QEdA6zaAX2H73miGZWxBDETcg21xBnqSLlh
guH9JEkoMs5FBOhqdqi0DxsXOPCzWVb6cZrNpvOchxCBJlCK/T3u/xjC9oXM7tGpZkHNKXJ9kCu7
yN9Igahe4UjE6avHtkkJH0HsnPDAjUMyh4Zz7CKueHIlp//GdtIZVWrBie4bf9y3WH5XSssUmv2o
udpAMXNVDtcSqxYhn7lwyPSNYGPIR9mjkZsBlFEdhx0qzkigcFbHZjTO9Un3viJSQ4gfuzSCzjJE
HL4STUg+awjUHKny8hiMn0qj1E2RzqePdR5ciYHDn7j9eh1HAxBQX55oYwLBhYpIbvDCAaBl0agJ
pdSd5OljwFLqwgfS29o4Zj73Uv+xDKTyyoMLwoH+nQTYnpAGmKZ+Ti7ewsXG7iCNfe1JaXKB6LYc
uNxdcZdreoWw8Anr2oHoDuhb4+JOQN2gNE8XkOZWTjeqK3AdC94Wv4wyNP3aaKdAaX0BIEuEIf2h
nZcTzy4spMR7SfcQhx1PZTBxwdfi8/9JzrTFs2R7dCq9UXLCaJmougvssTKfWUpKY8LeMdokOx9L
6gi+RCzaSYzIHbRvZYHRRcjhpogNQKc2xXVTQ+R1RV/BYqm9v0y2cTTMOm3IKxc5SwewysYVqz8K
8XIQaiTmckQJjXc4nxXARYRTk+e3IIvLDlNUu35zNl2d2FpisVr3n7xpHMIrsAjBVYGDEM7O7CXg
ImjMrBdrbSoqkgWnnax6XXZS8y/E6ycCzhO5X1pXNCik+Hk79ATQMORms4XZ6goEU+xGIOaL2osO
pdJHq4fLrXXXx+hT7nMHz3ekfoRsievRkkWXwFwXg8iBYP5fjnPkH2XZvJESmlCGSQTnQjIYLNYo
yAfI8IJHqjIQeuAH6DTmVV7ZqFq8arJ6+TVFS1f3M9G79wp6ABBsL193iW272k/Aks9+xq7Smk3P
yjFRVL5CP6USx7R+ej8WFGpeGwBhgVX5LTWFsexHQCKadqpXHuQSHQ7dO6YY1B5xZ6PW2nrkG/60
30LguVBlSA/VPVrS968n4KGmche0fx5Sgc5LzWtZNyIIApQLAwuY2H7BcwiaxdrZTIm87QDhhcuf
cnLwZhtVM6sd2On+oyWl9vG116uhtDF2ywSDGpIzlrVNW/akpPFn2igSyEUQHjdM8salQs19kU3u
zN2F7kO7VkfoUF4J73/JSASt0zZxhBV62jYNlAJ6kKSZOu9RP52nbV8mJ3IL3+ch7Z7rtw5pTIAu
X/5Bhw80C2Mt33/p7j+PT7rZAN2eFiNzNl4HafZTYVN+c8f0yecXqMcnVa+Hp3oYBBQLlf4SnOR4
2UTmrx8RjRfIEh5msSkTxWb2KZJ2bIgMEVkfWv52ttMSjR7jVr2Lh4fWXPA7XK69pIzNrPYi+Dok
OAnqjGyGjsQP/Z8Bvr/gSIeRIfBZg24nfqpwFWnHF8WMybcvS1Don7UOTPZSX5IJ/48V7dYM9teX
tzIYMcPVScCbdhdQhqPqEFducDgMOtkLAGWMZDCxZHKdLw61Po6B+V5pgbdpnWC2RoipCbkQ7oy2
FRfIb5rfQjU3kzWJAxQ5WQVSxOkXPW6+ADA4Ai1vTfvz2s5IKHxQTqVNYiTRlJQLn+SsPgF3H7eS
m9y3suOXpMbqdiqx4jwjmZatky6Nxa6Fxt8OBi+jJDOcX8jTQ3+/nnrrM9zpmmCj6cuBiiaZnrxD
pTlF8wshnmnligYSXgwNKIEzs2edw+n59F+oPIqzKiLAR1d5JsERZHBCdkObIZfD+aZVufXUC7De
7JaLVpG4LmCYSe2EK8QLAKhZ1Hu0vlseh6MxeFbD5VTI1u9FUZLAaLDZovzvAyxAsPrpbvkjMGPm
w5Rf+zk4gadmzqD9VP7NVrNOpgovIywBj1rD78Tn5Zp1g4VsUh0/yxzvMziGc6Zy4VgCncZSAFzM
kkMmGJ2cBzG/XqOsz6wtYIFELFugbcZk5EUxrs63zpnB7pC2iCiE/zKUvoTJxxQIoIRmvVmImgYt
ffNQvoY4jYdpIoQT8kw3g24MSjD3pdE8XkANUhkFmp09qRK2+NeGDvpIBbN7piU1i1PRqpsuLRWM
9CCix8TJpFqMDjpE7+7Nq6CnzrDwChmS17jW4blEVFPCadot1gwKBb5qawisGQlhDPRtWuhfoX21
HoAtRMwmyFfwURyZD4eOs16LCuEsTZRZk3H0WK71+Nvx0ALI/7bsMqoVnB7RT++H8bvV2MlOp4rG
Wtjpi3ykeVsOKckFYLQ/UtZH8CPZYmYrjCL8Ik7LwOnKrgRtt8OzQSF5M2NqFHYOypoOJnFeuoy+
OeSd4FNjEUiK84eWORh0QB+l3d5ZX1StlxMV9isdTHVVxwFPIUdF3grTyEmm2PbB1KPLK/NXXNc7
Gk0dPaaaEQmSk3zruwbTVbToizERYcksrkz+uCCN1cwuhp5R6iE4/wWX2BPDpbNeuSBRafr9sX8F
bIwsIyQmr21m2hg81IGh0xHl+dLxea1gTC4JrVLSVZdQjJqeQedZ+ODTVL0/b8BSldJJAZ2p0MqS
MeYJ1fG4Cj8Ulk9DxeBd86G5tO2ba9lYgg1Hm/QwD9ajImPtAY5SzLVYyviTYg/sLaZRzBIiMqJg
+D1ukYEdOPutUEcDjp0a9Fui8ZzvhJ7S32hfHsfKSWH4WN3yaeCBjMDXSb+hMSG3YLiWKxT3G90u
s5+Md4swn4IhyhE70aMoVsYEzcNmPNsQwzJCCRFB4bk95/R3a5MQ9I5YM9ich6+WBgHPzFuxL3uZ
FtzrVcGFS+OgX/MlF6cfZIWTv4EBFDHJadgEOmwLAZYAuwUdqVsGkBJ0P7GXJ97hZT3ISHLemoLS
qdWY2zJFKQE++Zt0eD27H8G0Jx0LbxNQbO5LB06qBA5Cy+8vvTPe3P2Fq4AR4WPcx3uTToqnzU+v
cNnumNuYmOPJdva7STUi9hqzqwWkyiwKC4wwgoOvKlBbPtK1ekUsPgvpFfsDe/c47yRX7TUVj9VQ
zo0ELY+rHbTnZCCkuRIa0dCF4E9RbyhLBpsV6tK26zKTgE1ZB3QlUChoYkGHmwHAmzN8PCudTh7o
VHjFTFVxku/VFVWy2vVySiJl9AqjYpb1x1wBYrRFykrwKyTWU86J5dJI0OB7bnectS6wkliHej7T
TmEVqcH3Xk1a4nuV8c49y8yLjn+FZJhUSaZspmFdHtpJ1yDtybT3Vcbg05JUDhbIHoTOkjJw+zDI
G6lQIgSOPvbO8NbbpurApKQ/V0fRrLkN7NPfGVV4qgzmb7wl0wDP25zJnl8Lfv8xQGGV77l8ekyc
Pd2oM4P9URo08df02VLOR1pCZwP3WYzhzFMQU692PcA5kFinfz8X6QjEtY426IOYGKuTnFkKumZY
M3IkifbNBeOCmlwnBBshiy4ZnV/vzeEe4RPM8lEtwK5F+1YFKzZDInERjy89ORBDtQyUn1XdSltT
Iv/li3R87/VStbGcsbNjNYEv+6xFgDbS5kW/eO0nfxArx5wG+EG5j3I0NLALU6/b2SMKUOjzj8lX
QylrXW4VjTL4eVxKQ7bwSBOckqGEpbLJo0beBHsPt42NBfaOiW8XzXmYR4895aDkqFQxd8MtfGt+
q6oFafWvV6k1HYgYFRdReAqoZPAm9QZL1o8Uqcw9qnLCKJSznmmQMJTjqU99fOty30mizllqF96Y
HsKDOUyfWrSk6sUl//SLQpH9G31Bz4E4TkuNL3t9k5ValdAP6FUs6pP9WnsawfTL3lCh2q0HJQJF
a3KGDtrsacAoxQn8+N7h6k5tXHX7WbF8NSGFax98CP+malMxoQDxfAc3H3ZD8geiNNeAJQF1/Mt9
6445aY8RVfzIAOy2JKNQQVwl+zmu5jlsHwOARK5Gy89oT+47LhfZ68ZEEixrnh6gFvUTS9SKjc+V
8RdEMmZCmvXI0bpDX104yz9j4TwbbKkoky4ZXgxw++A9RWni4XIMzA2S1C59RGLitAvnmguMj+SZ
NcilqKzC6SzxtJPqQsWnxrytMBwRUCvSb6h/7eOg2Z/UoZPa0+Pc8Hn44UHTo5maE3AbTrUUd6qH
9lTZQfS/hX+wbVM3RsRxt2cdbXlhZAPnvgGuIFDchN+c9L15/B99Lv0b7rCOeDgH7PnwUuzjuI+j
UX9ZA1XWwhvy9pbgky11U/5LHKfr+YKHrcqGFe2C63fzjkA2bx3v6FXIGv974NmR3oPwWTjrpDhh
98eYQspu0G4IVLINxxy4FYOKvTOu49gSrVT0OH5AisF9kuNGsTDAiFGGCm134bu6hI9oRohVPNfx
AsrnuqoXOvzi2Zd2nAQpAi+FGm8zvOWQcUvUOBVmF90q8MysrRHF68rXra/5M+KiF1vl5YpNNjog
8Kjhq/kgWHiTZT6GaCKbozIGKATaS4Z8f7aynb8p+O7JLDLhQycVDzsrLhjaUrDLVLuszuTAatVC
iiuRl7WnYPtap2u7DTDLHn4Ixu/P7OV58Adb3Ga/5huPf4jaNTYU6lImxnhTSRQMirWLpZ5lD0VI
pTtTlCsTuv+wWwzon9UJwmpXlhNkUyT2Yd5xIhzYPWn0tYLa0yKFEpHJ8j4rxajtN4b8gGalxmKm
xSLXKMaaXhPGPC9iQWxVlMTiPL9i8VIIBpJtnbR2Q69ayjVapLyK5liJWuD/JBTW+fTTTSlohQwg
5R7U/pLgjajHZ2PwPOzDX+KVp7eIjwA8Y2ptKSW7nZFNpsYRCxaEQWzMqPgL0Q0SKpc/IZ1fzwiq
v42ObENgauOYv6cxA75/7tIqovbE+UczqZxbIuDtmtdqYR2etUGSoChNW7ZoGQmguN8QcrEHX9+t
igfL0hlN9gHq50P07trLfXFo2eChpPafFjobrmXhP32O8SqfnSFh5YWcaE26Z7YsmYI0IZDF53Ag
xgW1WV3/X0hAL5DZv3ufxYRbkG907gWSSBWaW62jC+Tt6v0gqd7cKHh9CLp9bHWeSCesDB5/hQkU
ltoWORIOxmt3p1ger0Fw2u4tZNNidvl2XLzswVorSU2lPoN+TJElfmnR6dEqnvvwWD5rGxeLutZ2
O4qkgjx873cRiFtxy/m+9OVr7wfF2LTQBXrD3ObAdQ8SX/3wvx2zkryQhrW6MEAs3p3QvbqTK+1U
cfAPaIm7TsYC9PEck8VliyIlBEdfc1c82ztpMxMrf3FjVc+wuZIcQPVR9BFrocjdfzsjv0vIEilZ
7pzauxlwZUczce2A4Ipjdu2/pEkUY4w1//u52llGzl9UM5d72tAmW8raFwwSsEVCjq88dkO1hvvb
ftypIcTsfpwte2bP5ZFmaAvc9OXKfVwGClo7SxIde24Au1iFYpffx3OGm4gPuugu9d+IQuQSNRBx
UBT8IsdxkMXczS8VCZalnCop9Le8kfIqK309gQH/zmoOKhrSMlesKyDC3AL8uruf0z+IWjYRQZVT
Koy0Tg5W4vZDDWgRtOnX0NPtvTPKacpcpSY+gRxHUIMsKPjjki0ksKRwtbvsWxZLfFvV51z2YjNJ
omavtK6/mVLBxVEmpERpqnYQ4BpIBrGd1XtertYGx5i2nxMcSWd9UrJk4H4NWxXvKr2tD61NRVvM
IBnuQZibA25BzIE/jgPQXattQi1q/8F1JW76znbQuBAMwWkzwJYaDTYBqS32qO2Eaq8eAh6CxQvZ
GyJBwtlOStKP3QrNuUTuIIet++D4kTsgbSVNiJTiPHMAUqM3j97hQBwjQlSsZUS8KZ+kMOYYb783
Mq4Rm0FNZRHE+/1xMnSHTsJO5ZUbLKIWvXfFGS36szsxzgeVSOlv7D92T67xxSNfpz/GvjE3w/oU
XOrZdw7a4ZKzRR2Xq5/NHweJfWPrRBnxTAeWuy1D36slw7v+IfQ+Me0KELdttYPwL70SQHNc4aRg
+MyWrUJsMG60SMiWd7hgthKOR9kd4OPviAOLOjB83ZEPXusvgsSadSqif9R0xre5eqwGFfSdZyTp
Avf3mQ+LkuwNgqtq2+heCzvyamGPL8XCbSbr45keDK2N6SGq+tYUmvMkE7tveNnklkB/yoEV9WIY
9rWkCahyhWcwCc7fPO7QSZ+t/zuGuAf39brf5NMxG4ZjunpC3Z0laDVQjqlMDITPNJelZIBYgbm4
cUUI0KGfkY8IBS1AFJa9sL4JbsKTRrpzdvYq0xRjszL4JCYU4XWLJejhXYZhEBpGWgve92H24Ln4
69TyP2GMxxDqIYGOVR3fxqBbdtit7Sdev6Pa9hYWztk/icGzvlI0kIZxo4f3btr1P51XKvNG5J61
u5iKujd1JvK16qKhBtff2QdXtGbTT+k6+bYBe57Rt8U4DP9V5AaWWy2FqgIOsNgzztb7lkmMInrs
DbH9M4iVqYE2DjSjAY9ejkGnjPPZTOXO2qggkvOzwX0jrWy5aA8LtTQdZ/wujx6gbKjjF6KN00fp
BB3vr5P76UlqwUyN96zv5CQlQ3VHzK/TmqtRjnGrTXi8Qwf8HBXc4y/djLoHJD8swrrJxmE+8xhA
SbcSeNHIFrmbjJiS3O/UbMwBcRKjS+HaiP1qbiryDD0PuLXDqCCtFEi8EWlHidV9Nnw16yO2cN1Y
zRcZBSvx8aSvSULwKHSq2lp6TgrKUvBR//NbB/78akTDqW3Y3CnJ1ISSLHI912kYMzVem9vBURAl
FKDP3+h8YHqlQmX9pMmCaqwRJCj2CA3Vsg9AXYqHpMm7IgPb5BheLk7/QpjpzEfnZC+f2fRm6gf3
k1YYEl4P4fUlzJ4tF9sKpZV6avEKGVwiVG04jQrdIJ5sXsLrvsL8DBiobxo00QEXSfvvA7rC4B+t
N31a0XR+aLIHjiKfwSN1NWPXxmEB+QxejqSzvJZgacnygiW3Mt5aaqCX7O4fQgnYSYtUVMG2ZSS6
Jpxa2b2FCWiMbQ8XYU6Y5ayf1uijszQJoAY6xHHA8Lt6euqRoNfu0h2orwKMn5Aj2iDCDufcIbus
QlGQgkKc4JG+jnMTSHATNiXWEcOGbrWvrB71mSWjaShncVuaTCearZEChaRq9kGrK9ayjsan5BgW
9+97QSi5ncjPXgOhnGdTy4OLsnbR1el9bnr7bwJHQqawTcuNf0t7pzJ9eBpjzNM71Hd6RKZwAVPm
3AR7HmZhW1/6lqcD9FKIjm4OzVgp72MfB3p5LA+aODbjs6VEZ5ZseB5r9zDtMAvs3RegC42U3zhy
KJtNju/QszAZ4MArF9A2xN6DIHIvzbEGLSmYcLY8W8lP0XFk38VjZn08hcogtgW46E6i4OSm4ztO
Crx8kfIp2CNhxXBxC/+enJwUpaoOVaHZPia7vKOR3YOYxg8tBATww8THW6+Vkxp19OFmKKpQcV8T
jBTkMvHVxTBnyEoIgczgT44Ia6gllc7U6jx0mkuunGtioA8ysw6vLGz1beIknCOj79+qm+taL+1J
oFDWnnMR9nEGwtKWaqlV8DQ98waWpF7OoaVUFVgV96t2SqBRuhrxUOx48NkoH4fmFfR0p9qgVH6e
jk9P09YWVJNq+bqlcMEeZa64IYMPNjVVjLUB4+hrdfLnqCroHiB1FtnRhNYUL+AoHhfOa+d0tHH0
oAh4RGLBDdnejOsUPXBbxr8Qx6EvpPuZPccugt4Lx2kyKsJOOjtqmKDwgP1fkQIm0YY/fk6V5/TH
Ub5Tri6s+VF1Zm/Ie1HZHYdssaaTE8lqWi5hf5w/1zbKAswutxnMlNxdaRfDzERJKAWys7jPt3yz
NTqCjX9YaC/1J8V488G2k15cczH4OriAzZxGW/9aYNEXKzw4TprMAunu1G23tqRFbY0CbyJYKxtm
JoCFtqctAXHkolGWvC5QBKuBUiAg32nXR8FZ79PXfgummJ5rIojxtOaONUtEbdcO6rnuNw6Zq8Xy
/OL+je620KaDuCEJHjjZop2fnI/dT6bpzUNyOkZbHVnmrPZM0+xG74nybp6Ta0nPBLqMFD8s2vzd
01MCDHFZhx1/QLRMBCri4564x8EVkHc7zfl2CMKnvVIsIVgnZe21dSaTD5ccGkWTqtcs/azv+AaR
4geSIGDKbMaPo6lNRitKUOJ2fHFH+5vFsnrh11wtDyJ2L+whS/lCBNlk07QRj8MFPaj8bFIT6Yra
1Krx2RrH22OF5gU/FgtwLH6wy6hqpMRcjFQfEenSGxwvz7cE5TlccyG0vdPpDPPYOuDXWe0+16By
vQtmmrRgRxtLKBpwk1EqQ3piKUCopmUz/hH+e/95zm99b4dijln7aU+F97bIk3yFa+mkTRpTxssW
5QYocsO0EPAiG0b9Prj3Qr72vTtGWzdkSEQ/64uRATYmwL0pYTUl2ApdER+xJWEi3784oCN9NIY+
qr71uFCG/8HTkIoI4xG9gfF53oTbP3Qz/wuEyMSzAZrWfgwnCh+vx7GnEReIqda7ITfPzIXITXol
3l9wsNci79ZohkgVhkpTYQf5G5G0dKNfpqiAuXQScqA+ixK9LYd/goHndCFy8mliRgsvgMHmJC2Q
e/C6zqIcBOKvG8zTj4Iol3VsVaeeXiyRyP6G1ugxSwE3zZZKpZ0YTieZuVMNFm3t/SaEVLRb93Df
2O9wXk+0bBF2wsAdNDMNKQJf+q6Q8ftoUNgaqedhn7IBUv/pTSR0b2fbVZWsNvpqOXVOhRT6nF5o
ncfQkYIGKxwX3Dzp3YDz+HEczudDvSgtReOj6j7UhHK4Oh5kd2LU4hjER6rvFRHfjT4cEMoVOyTq
95CWdMfHRbZSCb+PXiZ0mLm8gcjL0zsEcVe10cp6egsd0NTN3RNSfDoadfGMrBRqYvRayYweDunR
dKDBpDGhBkxd9DvxDkYSMfEDS8SodYOOE7zXJBOIhFfMQHged8EQ/PrRw+XLXo24wb+A8gZqOkQe
A8+SAkpIlMrQEKIa8u8zbWOimrkJJxGW9Ad09KDm1b1cPJcEWxTlsYpLSL+h7rcmEZ3ngGhEARFJ
ghnCrWLKF73SzMmUlK9baPxBxO/KcSwD+Lkdw/Zhlqt+f9oVXgGIqekcyS77yuTQmuAGbNVxoMsC
3CuSEOsXZthumUx0/AYi1bTUTsR3fU0VJbcV6DoAyYUOCCtN0UxNiCGgV0Iu3MeNnhRqR8URTdWV
qcHEs0V5qqiU/xIttKtBj9dtT3p3K3kqWA18EujqErg8XZPN+HL9Je4E2gzTBjA8/v7N+Wm6tAWI
eNj0h5K6yWajXd/irebm9xVRfOGi7UPC0c5oF1OEy90mf1GLsUjRdfZYcfro9L/OBQo0STmoSI+f
ggbjKDSqYYJuNOgkX84ybfL1ZgZ36Br2+eW73WQ9op3ZynoGo2lXW4aSLFy84aho9Xk+ySzfeukp
08MYwdRh6ji/G8hZd216dI3Zs1wzTXKeFkUIQc9FwhuRk7Gry/mRKJFeclsu2SuN3yFpETh6G0s8
L+2dYIs+r7aoFGMyBMizR9sYbLxbnR3+RnNAdmcIEFB5kAGvvCSQliNQTUkQKVA34d67fjSByiHT
IS3t6RQaPcp9i0ODDvsdAQfagp5cl1vwmcHE5su3kXQflZPJn7PT/nlZGxQK3p7EG9KGUY4mdLNu
IE1RTs91wUVlYCgsptuS+CO05d4LLO53izs6WYYBdxJtDB3s5eu5O0aNJAjhAg99lqPrWdxmOS2y
8BSXI+z+kQxmczC0OV0JWIuQZnI7X+3+A28/m2z2M2TGvKY+/fbd+3D0HeI1Ky9wlJ5wVjEHeQVo
Bz6qPua7Q3n1aeKleNyjUNQI+IGLrTHpPCYV24ILbT/oLE3wFtoHIhVudlzckP4DMorO+9xQxbfE
dxcNwBLEJlbuUa6rIXr4a0x3lQcNZp2u4TK5sJDXV8fPhWy7affO5ked79WHcT5jGP3yvQQJLrcu
iPZazwmczYYRZX4/Lj7w4hkNAAa0+0aY/kSlle+cljbmLMBkWMNpC2j8Gk86QqCUQygZ5dpQxm+k
U8PDm5GURn5NeD/OJMJYYzrXuhFhwjOPxpH1S+0sV7id3oo3X1lBXh6FDTAsGj/QGjnvukWlLMgJ
nGoOTqpJfz7rzYZEbP6kdC6iTsaJdRsWxChXV3iTmcBV4FB1mY5SSNAMVYoGLSk+m/wsXbnZhfQF
gvIBmPURlA0oIW33mb5GRpyKYco6KmRVAvlReheY+8NQN2xUfiJENiokqqxwzMDR9E+97a15iHte
8evF47q6A8QDzcvbo3GyKyAk1jYssfWuOLR6eEScWIsRewBbdodffvifldnLOL7uTIkdiDPcA93A
PC6R2UUv5RGoZOnIvIiZNKRXee8sJv5NOjp3BzT4xIRWwQkDRcJ8qZqYFacI/409b/1mxS81swbR
fleu0R32F+lAz6uHa2vEyY8l1cZKeLhIirgdJRsicy3hSuaMYeAGRroiR35EaFr/pOcIAKg9m/+z
skZfTac3TBtoEUM4tCmSq9lubKSR1ct2k0ac8JYREXGFbDRhHMEkrBGUPEgb1D7DuWIPONJpYzCK
sQz262Vg84wLLYJmqPru53P0gggU2vfOXsp2612IZIs5/uB2i02ZZJ/eMKgdgEoAgihPO+y7Yg5e
6OGcGbnwl22Yla8ei9vBpHhilmjaYOp4ZKhrqHeBobzIPOsn5MrikALtoQxX+vyGzGFmed/kMqh4
gJTTFaMZOb1ITmA0ZmisT4kKeNQesSTQd0PNh46nJWmiOjFPedGtD/sWOfKqAAXv11ncFOW1mcuk
nZZVtcz45XhP4352bCRDtcVMJvmMcW0VlJhTtWqtggaao8vmOU/iMtQe/5EIbIaBWD+bnFa2M1if
Fo/kTzk7X1QaGK8EzVnWy8ZPhjsoRqaMzPnJbaxmx2IlVLgIFynlcugYPrE3ypd9xX4CG0T2/ed3
fUj41h3sUD5ANrebyRLTxrF9KjIKrAZynpgiz5EA+ruMgwn5++f1vX3OwqNsDBYbSM4VmhMFVkRL
73PqvEqaDWAebyUnls99Xbgtr/wtbrX9+RzM+O6StKJtx0IlOJGPXR2A7ax7EZ3ytJvqwL1USeFO
ICZIw1eHfuNxQMgH/39pnp9RyxmpRHKm5tyrg+WDp3P1rLymaSEMwNStaCOs8V22oKgnvIgJ7Gul
kH3zVM6UM2koxz7nUTRy48iWGhbyW2JW3GPW9FLCL+MTrP7tvkME3br0bLPWUwY/kRqW0iCFKtuF
Ulz6woK+f5clpzfK/oJ0/1r9O1FPN3YSeUv+szVOjKr1JSZCkryHDr0rYJeKnlmCIvDhWNiEXIBI
YPgvG6dUgNJxmC0BJKvvU2vo2nPgmXnFP0G3ImUgWVbKPr/+ypMDWzTJ+v8DspKTpMa9eEQhj9Ng
VPGPBnmy9CUPHIyi81jEOdBMP5wW0nzQU411LWi2mWq77e1Aaw8GokbZ39CM5GpPC3a9TNWx+9uQ
GyadzXcO6B5Trobonwjph7IzEUujeWmH6wSEYrqFEJtYE2TXJu94mDmkRFK3y9EkZtN0jz7s0qdC
T+wfs9Avc2R1ko7VOBvAhNNjT0zIhjYDO61dLFdLcQkyvwSGsB1ArkoGhfaMcBrn38qEOi87qJy7
8Z/KLBh7AA2aHMjZF7EJc6u7LrB8gH+6FdiGgsAuV8U0fRfZCbrr4ROEiqkIOkCwZxlzK1HVxgu+
iXE7Ox3uq36VTfJXw72QSXNPaxSxx4mvGpMOm4JVPfeNxgUV717y5Wyxd6EJ31rTfAJixaqUjg99
AuRsI4cG0uGPuehSGYmxzO9BgbcHwbSMyF+H+nk6BwXK+NIAi7Eg7BrFlxlYjcWl6nDhEdCMvygY
slVBjZRkY+Qq0Rfs2yNeV5gMu1txh3HgzIBnB9Rn9ljCnHdVZgsgwVq1A5mg3mAfeoXMCoKJODWf
ffr5xW6KWLrnveuMWPkai7xh5zuVcjKAOm2KS8SokCU+cN+wJcHd/40pBkSBI+uCsqKV7r2K9yL7
k59jMQSr9UGP+4mm3F0YX96WYQO0AMCRoIsL1mkZ/BfwSIvkO5I/B9paMJqD7sVfJoo8qgjfriYn
VIvyjDDOfxBFT0g/U86dG0bEgtbkUP/ClstP2KoT7AghWEDjG/UOnof7ntyIjLn4cWgc9zd9MgQv
W06wazNVEiiddVYhxyTX094O596xczj0gHjFf+BDwz3ZHIbmSLUXDkW5ayWfncLtjACQZUSdhu/t
FuQCrXxgVsGFtFtvMAbtGqFGuTrDbs2enMM8yjb9Qg642zUs7TJfQFQe6OnSf0DOt35CcZMFze4t
Z+cfJ5ih6ff0LZabTr0khHnKmDQMY+PfwRBhVXQqDY7TTUOL9aTtx6l4YBFL3fySP9pyqxZ18vJt
0gJ5ay+AbwatQG/4OEApU2wEERut8w2wtxJWCQGwX9Scg248IG32XB82P5piPx+EfKYg8JUXItG8
U49hkYJbaUtBc78PrO5epcvqum8JUU+ZRNtGHOtRJgKqTgPhEj4nWmqfhL/ElB1XmYy81dnfuSlA
DoFkj8L4ha3rr18D7WjIbNOoNxkWmY7Jgr5Lil4BHC7lzLWgaMgBI12n1akibEf+jN7qIG4jSZao
c9z6GDRiaLbZ8mQ1l0Lbjdz7D17/l7M2whmsjRgTmOa7pFOvLPxfmwuFaDorvbc3gLqzwN7r0y6/
TU0QqoijhYC4as86OqJPjMMeKg3rxeCUoXcO3zfNb24UqBQdboyCRa4mQObrSPtioyR3lOqANlIL
asMuI+9q01InMMjGObZIy/2FThrAvu62CwF40JcMX6azkpQWNocH6gnE1cltdwNCfvyRVBsApTPP
fUBX1WBE/hf2vs4kLzKv/A+9mq9ZXIbYXvtrIGhhTR/BwhOtm5A/2CO+tjkREIV0ipHTrOZA162n
MEO+4NY20P8U8jdHBGMp+Hsi633THLewAiRNBLogq+Q8abZNXY/qiqw8rHFJjgZrbjbBJ6Ccxkrt
ArescMtMuumanrZrd+AoeQxrk9d02wmo5DIOwlNBlUuGUa4YcMCjR1GJ2GNJsE1TMhb/mcMy+F60
Y14++N4zTI39z/bHw9xZgXf5uzVRklbOurqt0xDTDbqqJ2dfAiF0rvmDqUp0oWGxw0QBB593rum4
tR5LVFseS5etdb1UqscQSdQIG3128/OJk9Zn5TTQuqqk00zbN/uMib2dKRv4wbZdMJX2KLdYUaFK
elJqtWql/P2If7SQZTn3VCOJPoRgyGdhSJEI6OlP96noyQh7THpy/bq/6zHk6XZu+wBxHYXF2xIB
lJSQYG/UdS7fa4+uoTq2xeCSRUjNoW0n44fGiYMSTERvStRkrunAD/f+5MalM94bzg0zfRWjq1LL
/pUMAbMs+zk/tDLoGiBCTMV5RsEReOmSeYbY1/hV0+W086umRONrA6C3V+1WLOr94luFuUVST2VO
BnR2bs2o+Xsk/ToHAIeDEbpmq8XA4YJxNFSYbVbplwG+T6YlFbn97jX8O7i4llebs/wbe+XuPMb8
znIvmGx78eSaSzApWSOAzOHiIgTqiB1uDYFJtXfEz9Aa99ORcBChZ8NAqRO66rSnBLCrwqmZr9uw
nMFrac4C2rUmxQRyf6gk1Dle5a26cowrzXfEOubGJEd9jY7Ng6fLBQWUqi08b96cc1dyvcQ4PsYi
RAOJXK+Q19+eYMpJ9hU1ZIpe+pEEcww14USszM/mMe+j+22DVFXWFJZh+/aK+U4EtbGFIIN4u4b+
qFD6sHAIZU8E1BTW6hVU4S5305c+PMu2jXoxRLCF8XgKi9nYNlF1rAz74RHTFxQgYfOkcU424F7C
bZZ96gjpfRFUVNrB0yS51R2lRmnhc1gXQMb/FHFdG5owgraejZs6ux4iUeOyoHUG+T7IinU4zHhX
aVmD9zxt8wviwLEDcjJckLrZLjw9VDsZRh4rlyNszZcyiN+eA7xWpT8H+nQwnbBp3CauwuLg4MlA
eTWS8s556/GTh9rB7N2wZ7L6DS/aqjXbMn5ft7m4jq13253J/t2G1i5VSq5sl1Cn/ju7CKs+Oo//
kmgDarbYCgGWnXUhBkoTbwUXM7yPpKYnHL6vb3lQNySGIhFkRFPTQa/mGwU+CdeFKPdsy5qjMlqu
g43ZYlqXpESA/ggAVQ6JDR6F0DFM2hP07LwwANalViq2HLA+fwHBU0zttEs2WaKCLCQnlTCbcjgz
pcJyXDlYo40KD1EIQOnhQMeomViKyh6qlvrno649vcqTmIs8Xwb6bNVwxwiO70NbClGwtz2TRhVf
RZuhqkWhp2Ahx9eZGLX8yjj4bIxHs2OHvW90kvgQx6nWARDDuQkxUOLCj2GMqcssPhmNzeICDr8Q
tT8m4mVpVoDzQJk2D0N7805oC7tRLpEwJWej4rcfnfKRKZdHAliPD+3CGW1GlknHQUyEu8o8cqbp
i2ikbEJRG57B3n0NTynBhgJXYqV9Y27YQC3uPwUsCvTZPT74xhksqJU2sJ8a+eO0hvLRhi4XTt0t
9XImi+aj3DT4adOV5YVIl/va6gWryFFxYZppAgXTDel4tYCCQ3hORfxWW/NCrk5uBPtrdaWLc6gT
hQ7MDui6W5qGpcKfafVWbJ1rWZMBKjWzJ/SZx0kkKm8B5/c0QF8yXR1y6OHuKT/ZzCLFAK4xFwny
hBWAyf78Hhmn42QhLVYrSfs6xxfdr99yv4KRr37Nc3Qz00+GGde3xDIYsp4351WpSequMgtMhqkP
H+f0KGTEureKEn1CqJBEYCAvQvbyoClAq8tcULetbehJNgubGeEqJmV9rdEkfldo1fxKtw2na4RR
XxzD94DEJsOp0z/cRSo7qjVecrIO8dmNkh3yLErQOnlXzLtvOQA4ceKdgg1mueTJyEMDwbL7R4WK
bavwifwyt3kiO2OcnxU3Zz/HPlBKIE93f2Ja2cmymBCwcQaGB5tOmQuB/iaXEI9XRzp5A4ilv8y5
okIlp5iHaKvaI1OVzA/IMnNlNti9vhnhcGG6AUJ7Y3rc1DA7BXu7hYxDFl9dCyDMY7Fn5Oz8BjB0
75sFGIfXzWcS7WGDOQb1L5s2rYJgb56ZYwrlnuG+fiBUsidbf4F64Ipo6Vc1cVfstTSZCu8Dl/qW
mKTfzdv69FoiSlR0tujUi3iQXqt1Sp/Mz/xw12yj0SSWhb82IouFnQbPBNzanhx8bClyfmrHZeID
jMU2e0o3miHgPjqb9nXxlJq4eKRAmG8Q+l3/2Xz5o6pncHh7LWLoRFd6xMe3KV/qfjVgKp3F4iBt
5XUg1BPIINb2qqtAjHUrbWtTHjC/qmEugZ5unXRkjdB+Ztkkj/t2GBDyiOoCwxzdZKzXglknUyhz
DBao9QX6zv4v2KYSqafyxtyR/wp+JoF7+pw4YhgdBllhfJYlxTBoISbGWc3hj+pB9EQE8dcMJoe7
w/HC8w8jmqldBuIBq3WcK344bscWKhxeaT8Le86r05KtKEBRyDvtpW7ek4hYEQeTdqGi8xB29IqS
Pf+IMuxsz+3QGS0MtKN4LUYw0NnCz7JR20udE1kuyzeeI4W8iIzj0w1A4cwWRZcJN9U738GOMm83
GiClIyGGvWIlorRMh/q8D8wRFhClng67MzB3QoWMYhWdfHRsJExY/NRxLwityRlGfiYh1rtqFYa6
ClXfVhsMXFD9gSokbewNGmTOkNxE+LZIgHvhF4viTNZehmafmgzwQvsWdR/CLssgmfRuLNvNvrQ0
ssQDcTjnP3DtQuukw7m1spI11dYCjByGfswCRrGNG9VgvhwVSFZqPY5+BpRIusctYQlo9xDue9rS
TN4SVgPeaR77IWozo3h95SpAUjZvxfPHTyh992/y+rigQ3Z3f9ftKTJo7UyVCW2iLxp9ylLBCOks
6UXjfyqTGvyLERDE3NIwt+RxsraPyjOMQr6abNXlmezDNBKa0KTHZMN6UZ9PowLnBRrdLkq7wdBf
N2V8iNJi7xfQx2UTPM5YRKIs5EOl4WWMT21KgOXaRT5Sa9wuUg9kiaCjWg0t3121PpGA4I00hnvj
i9kSKwg8tdWdxraIMrJn3bzh818S8abVo5hxXCys5ehSI5YMJNNwtF8lY8XDC+FZrXaCnRW3BuIU
jVEy0oYnkOqXgrkgdtsohbgBpJAK8QRSY7ywUXwIb2ze94xM8yXHAkHZFo6pBvvWGESkqg/pJSez
EJ9ht1pcYVTrhr/u5H1LdHOiHe5zY86AfjONNa/REBCHME2QEiui8aTRFE/2la6LmUkx3irxOVPm
Ho/WfJ5F0dgqecxzQ8rEE520eETnxvOVSQ9sGuPnWaphT/Mnq4kl4kJMANDBvOaUm60HzJc6nS2E
/hiOgVh5wzZ5+zf4Gk14NkKBypKAFyLjMMtirLQAJ6Wps3VPcDK1zqXNOF8ecE9CicUVUOPmuaes
LcyEpbck5HE425DX6qxEFi3AhI2vcOxCe+HNPRytiS7naSQplPZ7wU4LPHf0DqdeUm2rdWp7G/t5
ZMTIf02sTJTqrYDcK1P36KyQNBboKb+63xvYeD6QziTgFJmYapkMa6jgyT/zw40bNG6xQ3PIZuAr
eUwEK8Ytf2/S6lU7Q18fGbmU3TIPt4ZnONs21UEI93muXSf8p6WGKHXDznAfGcZkCOkWTVeKtbgj
/Qfj8vdQrcLgXe5CzvHGh5SixUuLaLGi0/hEsGP+yVwJmfWOUeijgPq20MEKpj6oC1hRWc5xzCr8
kbUwsY7ivtqz1kK3fERVmDI1YmeqXCj3nZrUqYss9apyETn1Za00fBup00X2fgy+QnK6rVEVmGZF
7gYNW6QSaUQrForNuYfrciRLa1QM68xA/MYAWlTZw5TuAIg93riYF78TzDdcA/OK4I/KkS91/ytA
KkEBTNNYlpK3n6PTBW0jQXeS4kr7J+4mvd7em9iRKmidqZNak+/7ZRKUIWTNTq0KBzMrZW9W9DD6
vuUwKKKrVyXcY4hfAQIpE3nRtc7qf7Eu6umuARx0MdECS5TJyA+LimOM7Tl0bbv7b04cS8lK5Csw
mVWtDLkskXN/6kdVRy3t/1DBefJRn10U5WsFlEJM4BTHownPdXH6rxt1ZXY/dzjvMeGVlOQVbCFv
KczC67CE0gj2CZgII3VDz4CrablSvSxWxaxa0Gj/FLQ/lAJWRKdpYZv6/qGljsTNVLUBCkZi0x3t
cucd43PMENGKr7MjF/INk3ynQL/bJ/c9e8xV5zE7p5ur19Pvo7xG62ToMGacYqNwiqn+vLffBvEj
deXqy8QKeyLFvChe9Mq++qMWkJPcKAj4NBy5eAf+i3+7SlYpzrHexAUF27yIylQOWpBTx2iNTa9a
cOK5Xy9y3etKggiV+APj0MEyaHGcPdYOLd5/xMAOdev6N1Xhf4BcrRlQifDuOwhnVA8A+xpIzHKw
j9cEe7w00KTDA5OUHlbx8lRo1cTU3nLh0nUyaWwlUiZ45tS9t2OUMIl2wEQsRQzPowN53sYb/WTS
DM8e/k+Ke99eo3GpIesdqkgA6q2hbxi+JY0AIl6BzHGPDv574dToEX1j+tZrjWwlW34TRrLuI66q
DpDVbpchLqCbDR3KHeRQbMamR7R4B5tGPTBn33bCKhybcBNSI352RFJgdRf2bKrD0yhDojapLdQo
pnrbvHWiQlHHgODQh/CbrSkWIlSXMdTF8UUy6PN2/5Qr/7s6MQYNBgxUwcZPnxcETUv0CyEKqPj7
0UJxhWeLP8/L+IbmXle6bN7GIJ8HhXZxYCU3+1jIiPrQh2e6JsPrXtCQ1dy5GnsNPg70oS9Yu6m9
I0LMi5Cf6gHuKdYax0Upeje6iRyYRFG6Pb7YeCqxq5Eb7PFSKC+49LrRj2xxZ73YjBXJBfj4WIf+
cGV7LXuzrTGYI2WLsAHnCWKMDfBus80H2ng2Dp56KmdgoCQCfBhZcMk6nz5X4cSfu2/OXTA01d/a
VlBymGTYm8lu6QlO6UmrtsAjNMUioYwnQF7rs1YE+Vw8wx414PJCmMHSEXHGJHn6UhAQ4TCffLo1
JasiUeb3gQoco3BWfuiJtXTr8PNkPdb5Pspz5sOeDeplpLzn22MQ1I2zAPHdMvq0mK9ulbXHx+E0
ur+AtkJgTKPDp7QrXHGVJeDF1MBM1UFIbTQpIAhyJsgxVWhZYq4TlpAyrygnExYAenWXbOjDUbwu
mc8ZzttJW2tHC4Oi/sNZhVRw8IyfHi7MEnJJPvHDBjl/Mzzp7YmE8Dil+3yp0nxEE7lsolTQ5kMr
VDMEG9wc0yipnptg7cKBrZo/he8toSpxkes+YDbH9LBT7RpYs3gF64etv/C+3hXCZCaNTOlYOZSa
1avhcUffbepqlzW1jXY5R979JvCi1Kt6pogS4qK7fM4IRDQhBPNJhFMyF7dtco9GcTQXj490dE+T
R5RJLlq2iTTBxoCENlgEb8z6SBxqqBIB5odrrEwzMIscaAwFk53WUIPZgFbWgHtQFipXx0PPx44D
kZVPbe7OOj8kkfBserifXJSNULyeWgRVQ6KiOkvj3Uw4efTG+hCt29kf8uj1fPFzV+EDoe4GRg+u
ebkj48JZv152XhrOz/UawHraObz38hLBbRy70s39KFmVVeZ3uJGnMrj/QYG8tA+f5yIBDshBUr5K
C4cSkGZyvSuY8Z/pj6/91YabgCVs4eLTA/nQDFcBdETVLM5/OsqtWDs0ANLaaDJgHWpuXdeecBuq
0AAbvnYlUYJLXZ4J0cCym8+mU/APXSsr85zlD8K1+00LKtoiROM3B4clf3vMTuE8tYnKtrHixNf9
OhzZnKaPjP0BhV5hv/ozP8hlM8T/zGkkYcI331UflZvh1wS9WfWbFNRtNilt5TAd7dAAGr6PvCWr
KITOEbZAcubnfxGYhq6T4YMWsuiPYPuPHy4Rid6A4QsKzGAOxL1xJa6S3ZCZ/bWtZ9eWw49LmBx1
ksib2RdX6sRk8T/HrpwmLRASbTMNU9U0MK00SmPe4h4GP+88S1JuwGCDPski6JVbT5fs6pT9eURk
Otwf/+yPcg5C2WbK+DH54X5LGhIkBZHD3c7ry7W/rYOyxgZ5BkC/kNIlDoRfA4qXnL0cN9e0phhq
AsgekTPwEvaXgqud9j3mHupMM17FyB+YsKn4lA01kpD9UFr8SvYd8vFDOfNLZ+fqiX6yMET5zkCX
nbUPXi2g/ep4+TI9KXkO6qOEG0PaJX6naoDtEvywwVcf2Qwb+/V5sjnt1FRH8OM6acrthiGzhufo
QTHUS9/3/XSdaOYGqwjb9/BXMxnTZtmv2BQYpT5t7qlz+DtYnHJzTxC3XFTEjLCdlqEpCNl4AEmK
BYrMwBaOJ8uuLwXQk6bn/hYFdXxIoFtO28Mqr1afQjbE10u7oODAEUr+AhwTeFTlz1qY+hJBKcDc
AToT3OBTB+M6cXZV4tFKtBBZdN3C10pOtlF1wbKeFKu7tysz8t5GU8+LPMUWLCFLyXsQj4TPagkD
g30l2J+GZp6+T60JT4uhH7CmSvwxoKbXr530XtlJ2D/VeGbwVvFyrqSMkiACqDvqdL6lS0Hhz798
Mhs6yURkMsyPfr7+e1WVjtADVx+KCVayOA9HS+t6xuNslURjHKaqATnqUP31p0hHQMDMYRIS9S6G
8QanRQwn33CCSkdjkUqdw2DGRvGRDEuSIEYqMrLoeYYFPxbLgLPk10rIyKwTYNTmXtlXxcIhv+68
TgsXnKb3FBgDg9GJx1FlB4/2Fi0LseGbKUuxZsM6GdpqqEWoTE/dM6mzLyYn846CdvKiC+SyV0BQ
Akl7uJMtZQ3VY8nIHbHWZumV7FQIY9V9V84Nlk2PNh09ppLXhqCIHNaguICoDIEWQ7SzaMC+eNFj
hPTck7beBUhXbKTJw1F50qKUybFCKlN3zf6tn408JgmoY3xHZfhNDwIfh63nGxCJJLvtF2uJEgnA
EicgZ3/O6EznExQoR8Zya+wBoPMtNvapBVVZd5YLxN4vppDK7O7SNR+y1kmYqAnWi3SUfBFc4DrJ
O4125DMaLN02YwT0qmhmOuqSt1ARQAj3F4av9q65JFDdKAO3QA0O8mQWTg03YbKcbfeWhC3smI79
WRTGjxh2Yp+DwkeytciK55WjuMQaPzMNk2kYlEHXGeFaJyXorfl5RCWP2IYSDlVSuXbLVdmXSiTm
f6mvmJCzLhd9Dfn5AZnCtoNPCVPZbOJw+aKU456rpKijm/2uIckohljlgjHwBaKLoi7LjWO3yOaB
YcIsLrCCFJ3gEYybXd53CyVlN5WxflJdrnEtl4QYFnmKj3emibH/kqlKc6CFUbB+vPv9Ad47IDdA
VKNoToYz2rJtJta4PLCX+Q4zVDwy4B9KTx1n1ZMVHJFnqv3DzBFDzO5hZtfD7qTuJ7PHQFkI8B2t
f39obD8HEtFJHT1FqbEhTfMTTJYUe9VZDMBF8H1KXxoam5DTHK2aPlZpokA41+mNgsRSV/m6eNuj
3FT9Vv1aQaJCEF9acFggiFdrXwcS5vnEMVRlWm1ivfQCoNcXJmu7PGmBLOVx00W43tuJUZ5Pwzzb
FlToF490N5+gbqyCu/HdWU2llW760+N3tPYQYG+3w3YHjkhc9Y6MUxMoREPILQOlI+udwC7o28qH
bsXHsne6bw4/0SIkbARZw2CXDEEm2QuEifqwjWLA2k7kFcfzXOacZb18Xm+ztJQs4FwbFpctyVbp
Js/ueGCVYWyj2h6uqfQeEeQnUw58VGu3wHGtAz7ywyyca/Q0GbhzhVE/Exsbl7f9/SXqPqlGLm3q
1EOmA0/SSnFFNccFkOiWi8TMAjI8YjihTcM4zKSL9HzQEK916GhZayjavOqB6NIrhueKYdwh+/dA
pWT5e1/GpAQ1SHVhd9E2H9KQn0WaUV2xQsI8YKPMrIR67NcOR5D8a1rfCzoBrA3zrS18mHHNQ7lT
Ef4LIO1v3dVMnrlVmT8iDdO9s1aWoeGKghQaBA2okYWWRMZGNdKm3fXuG2GJor+asC/Pg6JKDiUV
acQC/Osxhkw8LwyPhkUzS/rzECEvQ3sxUpzYydjn/6D395qePyKGaT/3XAbEALXXMaTKIgX7hw2q
OKWwD4rH/826xw9nsjaDcI/+CTXLB8Z20oGHIk4poXfMn+7u3Ij9lWfDiEVUYfQufPp1DXMbRqAh
MKM5q6fCYuvgzK5qlEBczhEvFBFBxIZ+w7ZHgSWzDaRgNdgEFfeGq1Hknig7/fzWHkntmuC/P6mJ
46MrzZqAMqAbAZyMua0ia7DJCd/MhRfgl6c1StkEQous3QmBJjl05kdt8/Vd15PSQ118BLNH/tgk
hqclDQgLsyAVHj+h+RnOS8Ag/bgJDNtx3MvjJeXhr39+Z2tJPOUshB3yfvzwo1bq8dYe2MwWC6h3
unxuO2OhGE4fJiuS+QCIQQQ9a8rtcJzJPVu+aGe2rCuFZROvlFAgBCq4cd6T1RXZmqfoD6IGhg9p
FusaBOTmx0jfngkfrIj5Pvp6Ucu3QVs9s92dvrgfZ/b2Q9h39iE4j9kxeNZLXyu2aX9L3SYPkE0r
tP25+gxDrOCeFfOhpruETrBXSt+o3V1UhPtXvtFuWpx7T1XAjAemZnJ1zFYnyQlJMiI2F0UgeBzc
hruUX/kacOUQgF+hIaL22rXy0xQA9LIvJh1+jOdxhtrwe51myds0qe62KV++hW/SxAQGj9YZ/1p3
gzdVtoxeG9YyX2jfJydWsVV26GGsyrkDrlWTjhZQevD9bdKOt2dXJaOPVX53+1LRLarKFHpRyoM8
ZuuweZObK5dltCzv2hrvwk1tutaEXVMQPdlebBvTPWt89S5Y9Vj31MPlhcy4rBASxR76j3eSNR+0
fHy2SMkZpsOZlEQazPFvWgW50/Y0Cres0n1ZjdsLwmD3vgb7SODlpasr2KS2VviAt/zXIk5tsp1k
BbvRTMgKzIuNz3WE7UFKWO5coNrkhtmBL5p13ix6Y02YVMLuc+64TE/0Yq5t73OSDmi+GgzcYwxx
177CgFelpKzvDli2VuSThUo583WD7zJ98pWONxh4/26xd5PT/+3Y5lPPK9uoOWctMxpDAfhZgQPi
rp/ssEsB9xISJnx8N5QR1pgYspoSIPN6cmVj27sFNNhoYfQt8cjhG/Ps2NHW8eSAuP42vqfOwE1m
3C/CY/8vmC2QE6QLUoSwciTVuSPJRFS+sTiXHYsqB4xLKzhlrL5YEJZUEi4puvUnRQHzzKdHk+pQ
wrnqIo+GPXLNst1DQ+PTsSlaPzW0kFa4eTOWx8tw7AnjGHlmcttGny5NdfNCBXOGpVQdAA6RzvdC
FkmEMdqMnepGy532lewSDQq/O55NVlYGJcU8LtTSKDH6vQl0FLgP0//J8oTfllq2p0kdBIzwQAaL
drsrlF1Q6cFHhM/Vn3165eKBDf6gBFJqhRfY6N4gUglErwig4TVMU1SqODijvd4xuJnPUOKkeuFl
3vJxE/rt5KZHK57HWPG9UhEgy5//0YL0/9gH22kZC0+aH693C2JTOAXnXTg7igNr9uSBEBy9EDPu
PYPe3SJtNvOJjn3O2NcBYWEIylY68+q+v5UOOBMtjDtB0IU2ndcbVoMZS80o0f6txY2Kp+IZ6iL/
MYdjt2+HO77ZdRF68Uw+/8UrXgIZxPh4VOSpEPpp06YsFpgGAXG6FEPMgvyM+mhYCUK0GI8uPQzm
VQktGEoesrFpYjyIRSHlvXJwC7rXjk5jZ0Cr+LqkL4ClA2DtkJRmmPQhSiRVZomZkcUqH5R3go6u
MAUI0S6HCoN3BoVnsvoqUkUzVdrSd+KYkDJmx3iRVZ7jntzK1F8Y/S7C6ossK02V+S8TKFCFZVww
rB8+bHKmz8KJiUVeYe9Uyo9jrns75R9ynwlgi4uoWNRoRgtdTqMeDN7WueDMQjObOnTjvphxc16/
1VsNftKoesc1307mIHvY9mAZGAswSg9dAPlHPjuxOyyf3bRikRNBGFOM2LKV4KjaXOpMmHfxnjg4
rQePekGnzdDRIa9ROKA5/pKZeRT1UW0+TlnMPHYgNB5jhwHyuUHFDktCK0YjXaeZsI44wU8ZuIVo
ON99VEdi4ptMcbvmClJ4VQ4w6+Z4WiyLQvbqe/TEUD49RuutiAm3wLiwxCi4XO47FCU0CZtcW0uf
9BCYbnLJM3BHaUnVF5XT8CWalW5CcO7a8Koeh9H8/4TzUYqpHDqaTcJVcsZASzswH3HZC+6IoHKI
B5jqIUtrkMgRUE2M9dq5fOso9Elgv/Ehi1d7bRRnfDN3sBjy0XL2v080yU8YS1vC2mt3J5Bfsml6
3t/Ev0n7GO8CM1hZWRNrpBUvLWbk3nkfVJ8TP4+etIlDLbVJIhMI73JQWbkffHxj/IK9g1e/Eh4A
mfCF5n+fYTyhVke3ENznmeAtOVkGTBnGY1Hg+lxxLMwmRde57fVaaIVZLWHP1YwxfYuHhG/m7iaA
7mRR33HruoImNpWy8+dPEF3vRDQKOnaNW+Onm2kJ9kJ4zDEJh7I/S8i4i6c3hR34VQAz4oZobJFV
nTwvfXoJ9p6PGE/3ZpBcWSWSB4dE4USCwhaoE/MsaTZlsbE7LUSpTEtXYK9lpcK5LXCk0fhZqyEd
XRzfwRlLV0therrLZF8ZEb6LvaIyDZ72AJKgwqhD0fh7EAbBq6JWjLSfv25gYkiprtEZBEVeg1kQ
fAph5T3e5QnMm+Y+SMeZFmnrrDfKGKQAghHrz12rKrxH2m38yl7MD5a6nM7uo1VztfYJBI99zCCi
l3DE+LaLFDy+OVThvMQWD8BG58ulTAFUgg1g+xJSMTlURsrS5I9V7HO3XH3r7C1tH2EJE3NocngJ
HStrqRtJGp1AzM5+2HL+EVlkNkDwik1Pje9QMvNBU1tqojSGK1sK/9EKxsor1S0VlsrY53/e9Y7c
r4lckUH+S4L5ZkxObOR3fHPpOHkKL+tdIT2Z7tX4xo9DSoslHF2LBWaUiUwP3DGjBWN+jtPzRGkS
C2GAxJL73MzsH2L6OT3vZHJfJo0rxHijhzFu5QY68UYE3X5OMRWswtVb9k2QyZQ/lZEWoaDjrVbH
2Tu0EOxGJg8e50MoNiGjktQMX0qwq3H+A7JfMJdTqEYJyI9QVUow8Q4fLqeeHtsDcJzGVVUljoD7
ecbWvnbFX48ysihVuh4sWWNSkVxv6t8v5nNZ7Uw48uEbE8QslxmjoXe3uGJ1VBp2lWpTo0H7hazy
l/rG0o9qeDyvzWwUMqw60kOIwo6aHudibstbK/K/6SNkD9dz6CP2sPOq5m1te5TKmDkxMiYqgxz8
KsRg/gHheRCiYMlhDOqOOfV9tEpUytyYw7XjBUd5Q7mRyV+q37XSSmIWdJJ8uVFYSaZLEN5VYbwe
dJSPsijpVR0CuiKmQpywi7bhzmGHOHAERZ9ot2Dd5qKiZMDaTiqsSruG2fOqlCtYiNnyaASB9Q2Y
mXk1wX4ze3yMbIe3UkJhgUQ962vy3kcWlyl6+AkOh4Ds8AGDjpXR2BUClh1tflqCFAEtO5pW0Vec
MWTCOpb1mh6Ia+QlD2xr1TU1OerWBnkI73yWWswPr33c7bO/iQiBOt34k3Jx3SPHnZYQpsyV8yKJ
NxbTr9r2NCAHOJ0/IIP7JsEM6H+M1ekOm0GDsygBMKnAJEoOg+4dzq3kJRDP/Fmk54tq8wnhWk3q
3ziPsNoTSEyUNKeWXnBSVHZsheYZp1Fb/blMpb3g8t2mOz92TJf5xy/P7BCNqDtjeEV+8jT3JXWx
dzz+rVUsUUX5pkYDlWLof8RpKVF6rKdM4qHTAs1BaI9K6KzV+CDkc3VyCU9wXXYiGsmGIw8Zovfv
UOUisWh7JQmSg6RscmAXtL6ggcGtFnPJcmTLfcKuQgU09yJCBT+1o+t5vaxz7O/p0/xl3RROlIiA
mj4zJKYNCvOrP/mMJSvhIqYb8q5ggiBIfCorclLR1uFN8EU9lB04x5lBMduSpd/IbPrY/E8obDet
UI5X094y81dnsDz8v65GPxG6HjmMxarCi6MX6ixG4Y1EOJeL8ncrC/yWLtoLp1TubJOlPPg/PeaJ
rvHk2swUwttM7u0ZCG4UYdqKgoJSLtgYRN+QBUfReCUiqITIGw/N3O0j+xdLZyMNoHkoPBDa/gZv
NiW5orBFgoaoJjsiSDCccoCWpITftLNhymU6F/8wuYzWB6Fu+9HPZhvgvsBaFBMX2t58pT+IXSP7
ZfG8ovK1vgd7VeiQTFG8TdoSwSVzoo6Z4KkYZQ6A83AyWdN3EItDnTCB7dvbpdtycyn3PhZ+GAkC
GNV4rR1F7klxuvQF9Yzu8TGDIlGr4B6y+5wW8rZ0XcMdMOMrKEj6po+Lqg1RLA/20QPwrhqZqji7
uenEfLRINpQpwhh7p+9agEplzfrCKQVzIOocdFJom5bxbnBOVArk9xo+HpjhI0g7mN36eyKFpUHc
02P+CtHUI8mCMqiJyIJ9TP9Sgdp93DbsYbqT0RONG1u/OXEfBQEcnIjjMhk7zmYJABjyqasAhw8E
/pyZmWyc7tDA9ASLAAQq2w+36blDcJNQA2hjnqf8l4ehMNV00grrDO3lyjIASe2UrItuL/F3VpQ+
BVVHn5mte1tjSoBluMUY2HGdkxxQOcHKxW6kESburL81wYQEJsTjuVNU6HfwBma/0Ua59FxHi7++
Fo7rm54hd/ZHRqNaOOfJ8qq6IaKEV2RE4DTYpQQL8yA2fObNZhXNW9STRLPgS0iufbWsVIMciU8u
AepTPx/iheczj/LW6lEykQQzET8rgnkBzGISxAh0dAOBFp+ACbggqrHbycaZm3KRC1lyP49qDIEd
6v81CwugeMoG1jhF1AYCLai9V/tEQUwwReuUoqRwjZpWXXNMDeozbYRR6pHKjTRjEb3Zjg0qDiPm
9KqauZ0Us9Xd+LhmG0wCv5lttRJz3m8pGa4OsFxG7tjB/dVSwU5GwcvSpxI4VrFISNMt/yEWO8c3
CWTBWcdBwxLUi3vuZ+HNNhqPiTNxEdTHMfukVp54Y9X2pxxes9HHc1DEeIo6yEJpBiqOoYi8T/BV
mWnST7DBVMBzbL/7mZw1MCSctoOKlcp0VxOYP1Ub09zXvt+WC5eGOKRKfMJPSF3bzCfKjJloJSRk
rhKundrWXZJNn7cMHhZFHohk+I0KCOSwHQBt7CeFESB4dG6qAeqjEzRkjbiHuU/L8ng1l5cJd6WK
ydi5wec1tZJ/z3JGzwreXx+uA7kjAmNzcvYopKUR8uql0qJZYFbWc4MSG9TpLw/2QM+bKcGBYqXy
/mfp3dvSbJQHkoAZLP8ICdK/4oQ5kde4fmHNMnbvvP2K9LzKVxpB6JH9VNJo1/xDBaRFWJILi4kw
mlI4+yTOqKKJFA9nZh0InDI2HMt5jetdOkcY2lmSwtcqEHAYVRK2yZ9KyMTDxa2pklVEsSPcofcO
+DYdX3qEcr8uMdf5146vnJu3fiQJ2oBVBqMaNipglyH5e7Nrsdka1BkoBlIKKHnZcs40VdijuDpt
p+6mOrVwxAuES46XkD7tNGIv+iVc6nUedHpQuw1rfInR0u/DcK4kqtpbxonqwx/4oavXn5yXPWQF
0NlsBFLZR8GVhfPmCgN0+W/wyQdbuMm1kHRtJogmKULIu4L/94HqdtpMVlBQVdBwFC186i9e8RVE
Ha/3en77IcgS9b2pnxP4R/VoEtCk/IzOYk2wJyx7rwgPqJeknxZ1ZmKQwywdErYx5fI53gDVII2H
/AmPYSTrc57+uDhOvTCIdd57gjX6dRC/jGfhDb8mK5TQkfZ8Yde6kTpTQZMEvmF/7hJccoROipHn
CovqlgxRAAniJhEib4rdLX1oMjSqnyX/eQPVZJhQ2AaBsXNkgniLlO3cj9rhvRsFUWpJj3HjobWN
YGicjzsZTodZ+btP4UpqrDKh/ZbZc9H1cPwG5MCzKxqyYu5tJqY5SSmzOErlqOaE8r7nCCRxETZO
1ugksduyD6Ny/ZuOQUJ5OtkuX0zjGOQHDvWVnDSqDchdOkpTC7SUsqebozunebht/h9UJODA0VaI
gNT0G+LADB/xKk2HaxXXFPrvEN5WezZNQ4w2PqRQPpM7wt3lfeiN/IfS4tVSRDy/5HO81tUYmMWg
UPCmAMOopSSAKX+/DS5qZoX3mEWMHrN3iQTjKpKj8kwxfJjbvCoibbsrfW3z6NXUB7hzi+8akES+
/8VZy5gOO1nsZ89JLYe5cqaqGXNGhh0xZk14nPSx9EhrAaIcTtlfSKyTaTaZ945nKdXlweN/MCeu
hZE7y+zWEpbBjeS0hcap+K0uS4DIHbG2wttuxOkJIsW6tAuCPUZh2/JFaYSV4Lmiy1SiaQzczK08
3jisEGdmwMUv5qSjENxxVZyyfVIcgC5yKGIvGZkhkEXlXmkcxSZ6pGpCNrikAqYzXRYDeoiIhLpa
An5drbLTGym9OOVLL3FYFUcqoaLr0LYfOZm8FX7Upb5zVtVnlrFXuukvki1OCeOfVUFimI8j84Ic
AoTm5QgcHuZibc6CCsSTL3a4LHL+38IlOT8uDPA4bpqy5nH+i4hZq81hKLHNEEXssvQeXGol8MnL
YfdTcpltFYaB76TXg7SttOjfumMfeYVwekzSLY/GOFUFq+Xtbbn0Sz5HIU9upMTYrixLNfOJ0ms0
FED3CVTrgI5+yj05SYme6XTCMi5IHdXgVq02VmjBq2hhr44jxf1ry97Q1pI8+wFqNRXPSueqpRgy
Q4wnc4ieM+s5mGKgBuB++MfDIim9UVBjEQxo8gE6P8dQ0NZLpLy13rk+YXaXwqpsIFGirtejUpPv
fnjex+aOIZxpUXKbTFxzv3Qv/aPEYd8ksl2z7Rg9mSshKkI79dIbEEOhyMkDT7x6pQQd6PA5Hx0k
MEaI6Uu5FOQWeH7/OFw4+JU042yBDWL+2iWdDdVHsw+0io/PT2rZ6taH74b2R1HEmAU/UxGotIg3
QGW2EDArVrpxj3NW6wSZAz64XDGURrbMbnbCl+CSGxipgk2N6HlZ3jyCH/lwYDyay6rHy01vHObj
iUw2Vl4hp0F64sjDktsxtbFHra4RPtg74+f78mrL6Y48TLVbq9YJ0EaJJaQoqImaxbbd6irtSkcS
VGXXS79jvc7NVN2EqF7yaErNzHjy2PgT/147AL6LAtdVDuB9pGQLHj6owbNNc9byvctIRAbGufiN
JO/qZNIPYgvOqPMlzCitiyvbcx2rXG2hQZj+51O8P7+8ZkTPqGPHYgzTsYNeFSSLaFvw2cHGioKZ
YRwoBORKsIXLs05AlHIdP+Lj/UB+oBmJHcZFANBKxGRnwlQpIoxUdkB3sf0dDUdIueZBWr8cIBo/
9Fu1FNmF2lrZiPrzuWVHgI8V8bxLIEX5sezuM1SaRuNby8TM5rhIl8/UUR2fyuZjVdbNMbLtbEHI
MSvG1ohNh+YDV52gqi3jF9P7yWCRxkv6/KxboY49VbcTbU1F4cH068ruynG89w3Hm5Xm/4SZZYT1
4ReEPyRlJTHS0vfCzDWe5BjD/NNJ7mNKHPf4cb5Gtf0nneQ/Ldzpn9Cn1eGcclQdLSH0RuLxpvN0
IUh7V5wbQ9nU04/WJ/9Siq8QE2jc+CGEUGqmeBEIfKw8vDM+NTE0dbDboEPXA6MCubWgbblzmoAx
33Lajtp5AWZIYl/i6atP8/72Kc1SYstYM7B3X7+SaPnVBkNcHZK/mA7eNs3e+1g2v09ZRCuaiRCe
zloEifQYUV0Yn/DxJVjODOAsbGeiTb5fmiyGV198G8G4fYtRCWqcE9coqQqdupSuXLdy0DwAUrYC
UhhJoOAHGQBbiFJ69TRD643aYpr9WylJzjTDjYYbiNXHhPAcsviZI02jFts0wwQbl22fboAST+Mp
3an/uNbTS/jUqLbYD/V7wi5G3ksHWXojyB3LQzw9cyMIcJgZK4VPIEbuRI4CoOPriPUS0MLiFgwU
1QjXVj3SfqLHjRV9yoGh/lUFlpCiQotMKl7uqSWhXGmLPvft0OuExb8RkZfeV7ImzjB3UFvBfMac
72PPyi+W/knqiKaX7rQ8j2fY1EjPK95UKsYSMpQSKxQ74IUTLMXK7fzgsNp0c7FI+gTnnKCJX1up
F5CiFrwPdoJsP7XUZXmy+YdXlioWZ9fM/B2Gku6cvZpy4eaMSu9skr74VZ7lv2inuNP+IzPBoupE
Fs3QUU9fVkMV7DfBE7vxG20HaxcxwgfcxMiLcHBCz7jRfy/aYOs8tnqNi1lFvjbaJIpbJvD/AOni
Eav3j8DBU6eSlzuzQUn6EPKQtLEmvt9exuPKUv9j+BCq6nX1qDBZiGzgBhh7NEDZaJJqe0aR3arp
glpG9M2IgXSWr2uxH6c/8iuC6iRbrwnVTi54VyI29U/MU3wU1BtZGkL9hbfsOPJAvqGgEVuE5PaI
PsO4GSRl2H8pojWfv6tgborhuyYmTohqTsQa/bgvx0uhvtU5S8fpPRpXATmGJSz+7nKvT7wxIJ4a
E/LGufUfqPjTjlbT4IBTbzCAXw3FzI+ASFxMimXEnShb5PtwKEWqOaoO8x7eYuMTBQgqq0JEsPoR
GFmFjCslZq251bSVElpF9PKP1+ZmUVZKzVkb3A/Qv5C/+x46KUDIvfg1jq0cQuc9TW4AHwOLCAL/
sjqZEJpfSK2Lx7TynVVuZi4YdYa3UsfHPJgC6h7+9SHgI2/Wp5ET+Lz3x3JTFicRFNwF7K3Vgu70
3x6O5mHTh+V7lhe5wgeeN62SKziXonoBUanipJSGA/Hk+1q+S97iGasuTKvWQDbDof3np4DH3Sp/
8Zz6nPJaRXGkbSCqmrLIHHBEuMl3RLnPAgqcJU/Jp8TcmrGTWBlaARTRREVHkCWPk2UZnl2F6+/p
Zo95HXk+28dMcVowb7whrKRHu66MHoSVfzQ//8AAlV5nTJhAvd0C71qs7Eilb8VUMB8RKbsLOPsD
xPYTZQwje4c+nP0IPjz58gIVLZaS8TiqysOIXdNID4YQROPzdP5Nanp5aTF8kMTPtkons40JFC0w
akpQtHto1YGVaURfOOnXJL7374S19v585OenfIOaiIpNhxgWbf8wQh95D6STq00NspOfDqNOxnuY
6ZyRGrrZNKp+hNYpEQ7NjW9mAoqGwjbnwT4qV2OBZ3Gel4wBRXkYFVvbRLDrvzmmHUPfGHT3jJDv
It9/HBmg7esHVWA6SS8Xdcdgqnu5jOU+W0IUF6HBKNpJ8pmjBPojy+vxj38kFkE5ruffoZucl1ND
aw+CM/n78BNKqVwP7S6mOAghJSEuRBf4wI7v2+wXG77H65zodOE7qg4kh0nG2eWFXLeI8Zr+RNVH
z9gi/W2D3HnOK1D1pSidX3KuyxS/OPgJrlHizwHO96IU/WVUJqP2T9i4Q1xWQkz/KswbUR6Hot7k
nV9A4pM2LRz9odUxovzTwx36dTcr3qSW5rhKkkORVupzzyQY0ZjErojTz0UPpsAGQt97zvwHP2Ec
OyTeDqnHLx+aNE5fAAqEae2eSSuAvh0CJJWkgy1MD9Z7qEqRH6kF4ero4cytoYy0nz58X5ma0nwy
QcT4B1GvGsLiq//5Et51CU2QV3DtkOHkhJIexnyKpcQvRJvlHbs/ik92PkuyCvs3JzwWa5TarH0V
0Gk34LpehdtetLV/2/Lyb/wIGm79fW8C6Spw37y2r2MSf46t/FHnX3jhbSDxCUiOH7pvrmn0PPdk
O9dVahCOKKqGUq/UiML8mmP+ynNSLSRnKOh7bWbWup6OEu0TGa1zVVQTEUtq4ve4fSVPgnoGEsry
dD+n32ELciRdCIX5LpPaRvhz8528MqylhYWxAea/eMScSqTWbiM7sdJdwjbrWkGsS76mHo/q6If9
TTBrBmdatd51nnokid7X1uUN+xxBGVf7aQglhEl5cV87maWyivdd5f5O3WQQXyIU/nC+f1zrhstc
KQy3VTlZ8FW0mVA+iC0Dde/UxRBusUPfUHN/6RZbwTIWwrrezSOSit08lti9EHLMLmekm1qOFFlA
msOIBwzzd4dT8iY27yR6zcBdrsfa5eQVJANq4O/GdPsMB/9rh+YQs3dPHU2W86Qo5kN6XDTTqclp
xkDVdjIUDQTrEuZiUMJyLJzN9tzu4ls9xjrJy2507XAWSVYl3g9ucxDSDadvKvcDXLjHhT4hJ7oS
UKVzMeuK73GtTw8tL5myKF0FXk9I1AuLEcjo9Zzea96c1GyTXo2MHKMdFmunLul1jNi7HF0N0mTB
Gy2ASGXBALouw2atC2tUxy4TSiAaxAR1eziwXde3RFpG+IpGGUEPeRzJ44hsp2oWfetBx/mvyFDd
woaqFkuYH+jmARW4Q3uBFBytpG939kqMt2RHvYdaeIBfbI0HO6NMXvzmBhG2LAuFwlS9c3JVVtfm
xUSRvKAw+mwk/UIy1B7FUvTNeoKVpxRkydjcYEj+a+LqleRmh8ShIVt5niwuRgUWHNdvP+h8bGo9
4nvzHNqTKSb8RWMby2yQDsjX0ou2FCq7GEQImrN9dCgpchF+rbzlGMpIVhmkvQnT5vcal1mSrd6P
BnVu9CJ4qnocVyeY6eQBYrrfbJ4ZqqWMRgKwG44BUG5OlVZwcG3rwfxx11xuEzuIMtFt5oyWmgJF
dMyJ88lfUacblbSJUwSi+c/5GQgZZdbexKnv+kOfh9TfamsUQ/k7fgBeY/Bn3wxH9tNMGPhAgrtj
kGqKxDC1np1ZXkMXQLcmshE4ERgv4/kml6s1DLtJYnF8DPEUghHJNpmGf3UdZASB8zfTlCzcjK1I
jowMn8az0O8w0ItG8VfB4mkDoXmTtGrEFXMn6rHuzTSP5CWSHCJZFSIkF1HHSZ9titdP9o8jXqbP
JsWq0Jzm5qV0Y4kcFvX2IxYWfl6nft+2knrEK+Vq+mTW1yyhEfSDYhpQTvdnjJUJ4JgtGTlsR9hi
Xp7aXycErtB5FkWW6gzviVC7lzwGCWN5qHZR2N/iIR59J8Z0pmJwz/cn5I8FH2fqtyoyIljchBUE
B9qQvBzz/5UCFr75G9/HFURbgSsMpR4vWX8n4rIjKCDqowjvx+G1O/GH4/oruGa7gMJNg14usWCn
zzAFQA/b0eZB+eCmJdiQkuyBvHSiygG/6RERgUPWSrCCn8r/nf9aKv6/XYG/1+zk1Iy6K6BSrbT+
Mbgggo1989hEaYF7xw2l2A9C8nKdGtyO5nNssJ8YgNENSD81jyAd47L1zzxhzd4rUp3CNnJdzBCW
UZuPUqFdrckdPvuCQOp5v6TVhmliBQtw8SnEKv6+8pMF0c/OTYAvX1eMcpEkZljzH+OGGrjqZksD
LWCtqeJTYJrvCPDnmrKoqqbcffsDORVito0ORF/ckOwrJpn1cuZFaYzfdPtA6muldsF5/GSTd4Fh
bjhFPtTbw9/khwZh5+DeIBRdTsG6Hqy196OyT9lBPAjMGjfqsfdKRKrI16i0svKP7ZmlHE976JVA
pqCnWGJ7AmYn3blUmjmN/CATo7Qnk8qo4Il2JBhG3yIsdhSXpzU2wiOJk+f/4qYcfxsEA5D3wynp
Oa+CqJmjNYOtHXQ38DCbDv6lz1ZrxWwuNamAVJhNJcV4T3mcwV4f3Hyacd/1aQNNw05+lerDvGyV
QFNs125lEc1tA1g7w4AShSsRuWmDIHWkZwAT9YjYAJTmVMQgZJO9e6uNRTS/PTqASMRok54QVGEi
Jmr/XVRiv3AUYpQl8ytB8s4Zn0YIzXff7/h3NtBsK3ThcQsgQBfm12a7D8AeGzXwmHCZj0Lo6Qld
C3TyWu8BvtQKBqnwxJ9mv4B6MhAmGUAr+bNR9IMEOOy/6EO/zdWIP0vf3NCCTCyT1tTQ/Xgu38qe
MgG4g7Kv5Byr0YieHG0zQBsLoPwfwR1R9HATm4F5G1guVm7iw/chCV9Ci2TNdAN8t4+uNKIXDYXZ
s7D3NbQUWWfW3RpiskR3x7utd2aplsOwaK8J6TYv3MmXtPzXyj5hyn9tJVdTEiVKLLMJOJncuQ3J
Upz3Fds7S6EbsJqycva4/5rSWIqmod0pg2xe0d9bwQthD5NdPoEKGMjdejrdYDSVdM5TUe+zjEc1
QCCCRi74uzaOW2/Z9Ka0AWMTlodA3Rkyj3WBK83Grq7wXRMLeGRH2TTIVkSchsAVkrOVU3G4cLD2
/n76WPyEsnPAlazcg+yE5B3KLBLS1j+lxK5FWsyuSDIQuTy/VIMLRewqE6Mfti4qnG3Kf1AZk+tv
pRxUcDvTmYYAr0ar9ECSaGRdZsnAwTX7IhD0oy7Ax3DPTkPPaICIsiMNH42ug31PzvJg39hzOxk9
38VXxCR38NVnzcHtGgwsT1gxxp5ODRNQ6ocztVUod1cESDzZpprrKOjucp8JRjfCq/W5KuWVdJqv
8livbjpyLI6lCzeUMFLmLYLEzq2rsX1L1fZklJ1QXdby3IAie2LrUbnHKB+qQm/Q/PkKoa50Dk9X
LPMmcpt1Ud2HOeON83fmcguELRlIWbpMLZsAs0xnXyU3A9oS7HDhs8rB2jpF5hxRmHXEAStSnvfs
cAziK85hcJnesh8rng9lOMGwetg0oAZLOSJPX6hJKWTS4cQZbvdN9dcLNJq8OTIncsMtba5dWXjH
uX5YqP/bwn1dFJAksa9F4AO4zPRrWc+0KNDjSFKU6wI6hzO3xBYGZyubreXrIM7EeD/K1EKN0fBS
LzuNQKy5flSZdrygUIk9v3D6aL4hlVkwKSaaU2UJIzj9PLb9x3OtgF9amo0x33ck5QrbIhKXy0fH
xTltbyYf+Z3KtumfsxUIbY0H6flibBTGrqod0p6KTuCyqYuXE8L3hBI8jcp4QmondMDWblhOXMEP
F4+tjcENNquy2Iq4WAM952jFW4qolz9o9dxJ25X1yGUE/C+uJPO4S7dWJveZliBGkQ0miwdLPW9m
Dmy1iyEISJqS+tavKJRUA9rJzKecK71jtWdS2s+BOB64mpNDcJzFdVB9V5f+rm0woA75YHbn8rsx
kbpB2zVr5Hmz1juOfoiQMzBZQosmvYrPiYmqA8xzLjzTn2o82KqYV4Rdok1QTE0RRyNWpUrA9xrr
LH8RfAjoZrHKrTcIzrxWsxEAtK6D1Tmts6aa9jR+7da2mFEB6r7E15pBBXwolhlzHX3Wp8b2Ux70
3yyHoV4OTMgU8LCCN7mNDBG+GiFdEiB/Vw52tPDZyxSiwqHpvHMn1zVqFq/6xVqhgwBBtoUPjS8e
RN5zPET7bsyrJih8Fc9TBeP0GPjYpHHQvKimSIn4lU12G+FdQeX7AZ98KCP2vC4QIvkVEIpb61FC
q9kTuB7bhEIVb2Ra5FjTy/4dN6QmgDtWkZWg/u6BtZXQFm/tmRwI7g4A/QdlNXuktvyZpH+au+sq
pDDq+Vf/o4k/TuWetfIj35FjEtu++kqu9pmaFu2v2UCtKRcoO0pQzeDrGLnJnoGl6ADTVjF/mi0q
X5MUyiDeu28MPn+9aAMajrb0zm496dEomWJZurfyiKM+e5wpgGwK3YW8gzzgTZBSKwa3WUl5Iopg
ZXpDer9DLvouo/ONFiKc7Z/Bkpo7U9kukoRSUpwRjfwUyAycpjSmeWbeaJP6UmfOYO2fn9FSsf3S
e1dazsStXRhE7w7ehpUhIfgFJFwrd+Wwk39Zx1EVZzpUGE3hisJQr6MEgR08pCh1k0sKUvSMs3u7
c9WmiyLAiSF3CeAENNLx/kXdd640NDgSPGK/X6detjhiHAbcnFbuBQ/MqqOrUkP+S8fW3K2SfjHX
qqNmuy7coZqOg6Yq4WiTLkizJ3T5yQIOEuja8CNfAuPQaKs9u+N5hKJdGMqVXqP5OIBDrXSudJTu
XW+lUkVn64RcBcSOIGiRAj0XztVf0B63eBfVVacN2R30GYYf9E2Pnuf8cpqmSrY42goBiyYAYrB4
jtiJZa3LrukhD0TAw6KP/Dqy7+Y6DfAMEPU7FpxFyEg0CRKC8+yYvjAZI2AfwVfoBwTsNbNKgDy8
fgLsuGnYw2X+MKL+2i8bU6CVgJYMNFs2ebArBCHSBakEW9pCblnVJMnUjVyawK8qsfZHajwqGjD5
V4yR2fzJvpwO1pFZxIRiC+t5jLK7OHaJdJM6vTZAyvrUrIOmvEkB3JF+GFTkSajaaOLBJkRxjTXg
VnXIUiiLb+q+lu7/T37pGmLppO8VDVQERPLqsHPowQmyb64chxN2AdT0JW/IaizAbfezGYnDMMsF
0zi4nrxWAibI91oU7WELaXdIIQgtc1cdV2P+zZC0VfjDWNUefqhccWtrk/cjVPJqtV9EQDHAhiiw
uRtUpkoCmu8UhiwEdPlDfsJGLqQi6DpMwSLUdLlMpTBXNS2pLE0SrOEz89YsZ1wI00f1mLpOYkhj
UuoLL/zFd06j8LTZpEZsKfoTgfjUt/B+xyepNm5o6XCohRpdRov8ywo4YeI4Ze3A9elNdFA6QsF9
yC/2ZyEu4chrF0L82hk1f04L3K71k+EW5kDwVRrOigeADA/xJWU2ZsbAONnc40rmNoWUQrvwEjkF
L2yA9KHomD7SKDMwIZL63/utO/x193rzaym2gYXiFbHP+sYPoMKFEzplr2n4weQe9Rq36gUJO9kI
Kff1T2phZE/zdh2avSozXm+wWyuyIKyRX1l81seENr0jsTD24Qdm8Fb33Tmbnw3jivj+YD82zcCz
qBwUooUi7NHWcPVWGDEBz67LmuYFU8G1MKVMAB5JljughGbGIUMG40Z1U3Zy43vBfBfBENiKeTn6
NwBvtXxZ9EZr15DVe/yT6In+UMaEg28GhJjgZPeq11RxcohEZcymxjHS8RoxZGQFEhm9AUOD4Csp
2jW6qx2VpzfCWv1ulh5aYNNeJ1cjAd5ubQkJv1U7EYXYQTSjuQt00S+RhQA6slqwCcXAFI0GwpUY
XQVzbqMWPsNghUFG50D5J7jQJLBtlUeP+qIh11VOirirSzSfVmAJ82bD1GMZ9xD2yTMN1+hFLxne
DgsyyqUkUggBBCuf5pD0raVck5gD0iFG+m/xADNwz6xUVMkWNE88pGT+m2zZJSxXqN0rV8TSf84s
OFhdljT79sA/+EvQRv+TLRzsA227rLQk3fYQd1/RYwNvzCXmWFNivvnnR0NfB9xzvB8TtON4sBKm
tNJazPQ1+5Z1FCz5sBa2lrmuRMn4iFaVSzoYxOPct5eJa60FzCZ7jKF4KqfhWNticprnSjMjAGiO
f3p8n7g8GzLI4M62vF0sDi/UfKzNGKfmnpBynBXf1d9lYO0GlEXcssaDIFB6VestJZOIEXh3V+VO
aIf1BNJylkoe6NSMj/9b9WJHS6KOUX8ctGmu0NukoShA82cR8hBxj2EmHHnlQRZmrVL/yMAed3r0
TiNCGrRz0St71bXwh+ug3Lui2xS03flBtKJlJ3rLzKpGN7VxmU2j5ul/Wpurgxx8Pv3XG4JYmdYK
v0kluk9WJBm4KGGVlCH+1iYG/EQqXemyzK1icwLwnm8Bt2zGu9IDm9JV69wFFCbYgL4UhtskecF7
RWKIW8AxX71NSZ++kjD6kPQaTlXI6d46pcBg4SngMEfBULKXjvlmyC5+nyxBpVL5i27hpySnkyyq
EkBasiFBAmG/fnx46ecMxgvKr1T2dTkmlxsif8MVr6Qfbom1Z/QmoAd+0R5Jfl8DpaNt3hTZovfv
Q/7uU5XmkMRSjQREbp2bxqOBQWBsQU4kl6e9dY2JDw26sMur7rksyzKOUMZ9JDEUNsOvRmbHmwFy
mHpG2UqbausRNwjcJ794wm61iYB221ornE/9rahvbpdsMv9E3XkEMqGMTh6pR1oeKYhjOgEDrOvf
6sdHiPqMgyFQTdgC8r0msakH4zBgIkgoqibPSwSZ/TX1UQzGjL14pRqWQGGhNWosKI20PKcTuSSj
0mh+OZhXUssNDf/oFUMlNvDLrMoBMLx8HsKvlXHTIRJ0DfXYCtmUjuMD5WAWRfomVe37G4p8etOV
Yl73W5ZobPBu6jpqbYgnFtewA+0HWitC4swM/4MTFGgdcJqcjuQ2Hcmc4ENnnDEfbrHr7HhYMd9B
8sS0D4cePI3QnpmSdBNDymDLa2qmUVYE0Uj2KW8YIU1O3cv800WIJMdFK8WZWb7rrZFHZ/5Qa4ic
o6rUHhE4RlkApkhQ9j8csiXEFnFT9myrfXYGTphBMWQTF+9uin7+BEIR5Wsn8LLEaGDo4Lf8Z+ZH
mc6pLAgnLXEOmCcxo7k5bv9qoiSuQpA2Gz2jFjk73pbVUG59nokM+/g9HPapEBqZSDdxMgW3r1DO
R4WNVXlnLvahXk8qP6pKBLlbz17E7wzNP9Vozu957wUo2fVI/ah0VOpCltVc1aXriagmXxZZ+c8Y
XQ/HnuBpBonWZKD3zu03xi8QiOLJrCTvGaBcdhEKYrnJt+vAv5t+qgqGUK/UK3QXCVdzTb5KyXsI
6htbCDU6exgr6qolE+W0Qp1p23IzmLPO7ODZ7wvGe3/KLZIckO059TfJWu5zN1imQTMNmIk8WagL
2Ev/3O9JznAObt8jMauv49Wi1iZAbdx/h9x1lfMNcGqcKWODxD7g/9xGxavnZgP9TET51Mh3VcAD
HNGXL+iXr0mVoxnIhzaPuyJFZDXKOP19kD5uQHv43sqKurItCPbhbhhAqOis6MnC4bbkc4r0DOzY
mW4QI/tJm2+QLEFHSptAxyDbWKq6codtj3gfvHSu6u7Nos2q/OnZWLbBql+YqJgF0jMLqPTlpEli
n2k1omitUopSSsyaFw+fMuLIpZicZVNJTLCmUZ2D1T67zynKhBcSAD2PmxX0eZX87jK2/fpPa1Lx
qY5LZayaHpeE3JqXZQxV3mrQP9V8EXPSWvSM/9zWrIF/NiPb1eZVPy0SHvvkJ9hNhEA31wqGAY2Z
JCI+cQXiemjsmc9Aol4t/WYn/h+EGm3dRsSRPE59qUSMVJ2XoCTzKextMfZsiDfrhwZk4Jw9E9XZ
e/uV+0p1xWlMprAvjbt9t9D+pHNhV9tdWn5ew6s8GdUnAx2sQyB6X2iW4G+JA6uVJLyPDlDQM37+
wQ/LTZRqBtMjWxJWqE12K1v2LGQFoNLJizVp8nUmxZPKKViIRE561FmQiBAPHmrR7Gd9r6qsIFp1
IJ4yHaKtUEt+gKAFuEaDaCHdNuQePcfU/GKAtkWrTdyRDON1g0GwsbFiCJcDOkQ20Gz41iyITntq
PwMHkx8bCjMdEhJjVb+j4QCEm5bZXfRcO7jXXV4M6hy1n17c1ipTqyoAS7l+VLPo9aOYzqxSgj5T
04B2uEcuoeXt0Su8DAtbKw3SU/mMjW/eB0Be5T1Ypszn/EExjSWeMbQpWgicdZLZ/YSGhxOVsZEt
Vtw6gUVHHINneUHHKjP25a3iSBI6CscbmLWdcZagcZfoMvjooar2hEddgBPC1smhxr3QFTw/Orrs
+8HU+uUj5Kt1eertol9S6W12kT7pXBkkzwZT1QgNZ91JQzGErC/8FS9Klnyf5GpVroSt3gndlj+8
exBif5E3yIxQa+z9a99txBzDr06j/GYjvnAPoOifn0es2KsqG9c1f0rHFKT0eP1MylYbSPnouc4c
b2A4cariKaSTyua5lL7BlvasqxNgaRwSviHdvMaAk5DK3UzQaSzQ9RIN7QRfXhYRMZhSvKT6Xw0Z
QAFVpgP5u86gwuHyFlawm0BDy2lGNSCFWOJjtQFL+odeyu4xY30ZbUGK//FgJoadXP/fMn6ySV5y
b5QioTyKDaBJ+aOcV84Xkj9UwWtVtY6vwaFBAfq0lDSXl/EiLLpGzDoRkelriKsaDFr50EzRMKfd
WIyBzvscBdLSQUVe6ZS+4w9Neo+BgGxryKQ7qHdB0bTw3xPZaRc2OmadSbHQLGIuOyIecVUPv+O1
qs9EB1vCaPrc+jw0abD3f2R19UkfkUhuTTaKWaCiqgr4cAJK4wmRlfQkZ2YNzFbRFZkmwcLLWn/0
rS/KbaTp5pPPR+uxRoA0JQvSXwSr/wgHXh2M0aFpEhnMCNe+pamfePSpCxwOJNZyGGxc7UcY+9HJ
rpnXtpbKZZORFvo8GL0+YLn6AEng+z4l6n0bQMCNNRxAb0Y4ckcjzo4CwLaKFcpsgJ0tyC3E0wku
bjDTbzagWrpNiIVuSb6hWh8Al1P6iimSRuF+TmRDmEzSSveXtQlIuXM0UXsIa3zOdBmpG9Qb9Lcp
ZMPY3fCJed/X7DBt6cbVsK62johaI5A2wg2Kiv76wDRNk5KBn886DTWpkLirtPKNOFLwqT2JhEJh
qR2Spw05C4kYdq8coqmUEhhOzsIzbSKZzfmX/5t/Ao5/lvZ5h6fSEBFQnjUn6E0zZ3zb9uAG6ucz
St9OP5RPeUuZOsRAq0Y5HwmXwc+UR4xlwYlNd9fRhu/entOAreJEXpVjYNgiiDghq6mFHPXr+PWi
BuY6PP+VZRvJ5wA2QTEHeYOXAwsgq4Nt4H80MZs9Eqd2z6sZExmwLUqYKqpMod6dKERtHtpMRUgj
XFm880NXknpF+U2iKjST/y2wDpXaAs2JMo4j0yggZRzDM8alM/KE7QRRgKS/A7CIWP+32WD1/ntX
E0A6i0BIdxEHcXsTzpEeTIiLr+ps6UILe1CV0qKxqm1i9MzAMN4uLz7JCVo0s1MDWXuky+fFv41Q
Q9fK7yNlO7ke2Q8rLiOpvYGxRHMAV7+1+/EqCM787Ih/HYjwGQZeQm4MXEy27kigxkGD2v6mJUzG
0KcixsWHZr0kxB/t7277QD0ddccHPn0lkCnfoie6o6nuzrG6gM9xXc5qsXLwiL/R/fRwrqIoEIT9
QHIX9nrNIKvz4YvJZTR15rtLSYzLSIxkU0byVxPJlTOLDtSWXoB7XzgEFWI3CeJ3hf7Z4snXhSgr
Fwt1rrgCJRDE0f2J9g4pqFupgIMNiXvC8k1DEBANJkUfHH8Mfxv+gK5NSmGMRu5zTpgMkEwZfwXU
KbEVFXyEjIAQ0br78ByVNfT38z8ZaJrNHkLs+1iQtpN636YhHUU2FUCd1vUFSX685vsx7+SlCkgp
GeggERE2+umJnwzMKnNIO+B4+iT4D3PaQNex2T84tV1JxpbR7fDS15MUc2nh1+yqhuztz4cVsw6m
uvl2L2yK5kWpOFpq+BaO8hSqugLSNlHUMBIlJXBBrjo+ieZdjF6k164YQOAIlMpQ/lncx0HkX7Xw
AIEGI0CYjpxu4M/1kY++2e5aZJkjl5Mq8QBJYo+I64DLZRmN8mld/5KakwojVPyOFMjNuNU0pBS3
mhdTP2qLieEsWtj91mxi/i3U83HffeVg/WptDUi37S6i5BcpE5Jcot9GA9Ed/nXvGj1W06zcZpbu
e6cIczLglY056sqOOQsyh5hlctsvFG5NX/H/FfMIIwipkiS/dfK2elVvzj1Nc/z36HB8S8oXERzR
OU9HBclXb6Ozp0W9bX26DgE2h3Kq1GaKcSQIl6DEE4RVQCIcK1bArdlGkQ6EyYr+A1PwaBvNALBv
EnsWqwPuToRsHmvDB+REKGCAF/n1Uttdx1tqF0bU2u8flzLxm0Yvl3K7B31z68hcpVsvZxd9r6kt
RPaZsCaM1UnBWA1IkFU8cD/nC5i+JzpYnSYNfmzNVDqyeQvdxdrFVSaWUQlwWVwWrJ82jj6iD2Co
vYAWaN5xF+PzPiSwFm6yebWH56ZepopIJClX3aFHOXTYtuQEUdQvhxBRSJk6FVwrby3NMSQJ6DN6
6v1giWCxffTwLjWEUgWyX9H5AVcxufeEVnSGhgfmJVi0JBNCNPmjwrbmx0oEAvY6a6hMLLAbyWzl
VUFpUq4mRtnc6dsYXL6ObJjfOBIzJfHRVJXXG0PXwe7hdl3O7XaJg7626hQRqvROmYWghC33z/Lb
y8t/PNzgx4MU8wSAd36MO3dhNgfSexV0Zbq//UfH0YbGXPnj2QdNGBKxil9agGGNKTj9RZJJsp3N
COrlkdB1Iu5l7JJvAefAh/H+vXt8+wbje3R226KiG9IDQbZcE8oRPDVmfq28r6AVTncFFnj+2bFY
l2h/7rHgV4W0HU2bITcMQTwqI20Bkc7cSTYqua6U84VKqbgqAMexZ7MjYovNS8tA6MpucVTE1o+q
K9UlJSKczjYrkx+LTfQdkRKTFmV2UF5Iexh8jSL/zLOs1cVWzUcFcPOzIyfs583LgS8EhHpBUdGx
ivZEqMsgzE34JArjfJwgz6MSt7LotYuzrTivuDuPvlLEphundy8yvszcwbQfwrhjYYCQkr0Tc6+w
mEIky5Kub4QTWNf3kJS5euklhIKMKmsOfnPa+soYuzHe+6ZMKpGJBUyi4jzjJ4frT/Ox4uo07ViR
6bEB7IPEXsOuhiFAuUaFtLmT2VKK17yWmA6FNbtmWbBxY2Wsu/aE7PPudeN5epgHEGhSsoO5Vx3v
ID32EyAXH5s2KNAXdT/h3d9se+hqWSV1wNwFWybvRXyxN3zGt6z8iCY8vv5eHJvlYEHPbY5k0HkD
YFN0B7SdnYGvAau4gMy5Coq/gBHqW7L+7fQreSvo8M3a50Htwx8timFn+vuU94ev8HgIZjENB5qz
ahqrAxSk/HBrtdSYe5B34Ua6cam6VuqfAT3+NlgN4TU549NLVeqM+rCiSE9Gk7JdV+gB/cMg6fh5
JTFHPjThaQRc0AVQvMEO0MY6dX98ayES+kvnjqoLszeqG/7Y9mBXmx6j7A/Qhago+8m/HC+HSO8E
X3lgBtgi8OzZ/X92Z35cKTRiEW3lRsSE9x53J19eqzyz8Th60xnrv9Cvk90R49yJudyQXmNUiYbY
z6CmEvwHVXK/n9pgOQh7++k8ZYL4EuwunL9/e4uJX5CSyV5Tay9h15oBYyJMviypHK1p6EGBBNGx
vUJwWfhlTOY2c2dPYd2kYqECaa8ToBeR8pY2S6svx93wZtIcbNWjBFavMv7HTkszpNjFXrvO1Yv2
loHvW3n7nnFWouOeQyQ3kjLQJIMDsW9NlgSx/btsIHstOB74MYbHPUSwsLlNMJJow3V6eI0r/8h3
toXBe07nM3WopB8H7un15EPrj5j4GppUlnpbECAUWB7aEq2IXT7nneb5YRu1/xJvCnTkeY2M63kV
jVt09SG/g0QwHx4z7w5Yg5Ir3Iovkuek5Fy8dYu6IDOdWSu5VXaRCXTdw3lnyUutBdiMP6cGNSl1
6Ykr6TTuvnSjAvGXfhobjsDkDZpCZiTp3Dv3uemAJMine5IIdqtFSbanhpIVNJyfAyGRwlHJwz2S
/APQVbvprM7qCEgks3qpU6UsWv05su+Mvs4RvcHvQWltQhsx8l4ChD9Kpv/YRcwlcAorjMHHdogA
61kIDovrCSwZ9DLnR76dHWfptxscDV0hhvq9VPFy7dWoWbQHYJJ99ndNDgoybVEyLW7gSzAt9qEr
IjObnM0N9nQuchAcCtSYTACjS2k2dDPCeEWFGzxY5PbZATZIQSz9VL0Rc03Tz5H9LXcp50O8rezi
59uEI5/wczhn8Bya11lfLTjD0lVLyKcPZ8uELPswEo5ZQSpOisTYRDt5nyrQqrVj99s+d02iVPTO
iGs5NgmtHz1me4LrvmsC3t30ZzHjep+UUl6lLo/3CZyw3ynfFTDBn0dFwFo99PkdmxF99X3hlTcJ
ZuoQ9gFE37Z//qMIiUWF0zz+xnaMknXZkC03lpqsEJDRxxtZrlYiD8RCGtiTryYAXvBJupnj/Wko
ImNHUfCW+c/BYLLPhI2RgPMD84LJqJjLCt5yS24KqONt6+IOvfNIKuYmOfq4mUDNDQD1m+JP4byy
jREyZkedx6Yk3zZLYQfiXouM/Q9oxYXjZOy26eztBXwHuJHlllnwG/OPla31T676mhdgJUNw38Cw
K2D7iTG3ubk6XrcENrO/kgJiEaP7Eyz3dLul/zt1HdHTUyPbz6EPbulCmPa9rr8VMi9NnQ7j+euq
ISzxuSI4fQcRw43/vIqUuwOb08/wJJ/sDNMXZg9X4vZiLXNsdzwcwFDP5EQknTLIWT9L/z/J58uT
wq0NZSQbhT+oRdbhL7QqAd1Yc39wVR1W1BJ4HcbkCCG/0S0V1sbEJ+6OUzBDmW9dyszyVibB0Py2
tIYVOIQQhk5tfeMLlr55CKb7qsvnmT6umoR2JxOtgyg8cEEU/nlZOOkcaFrE8YuLQDh7tVRnodm3
WdrVymKN3JOcfSgbf7m/AlSYJTpz+Oc+LUci+lO1DEnvwQ7idcdW4eDg+8d/f4sFNVzXdW0Q1HHb
1ZMpkqXmnSIdlcDvx/oxVr6jzVYMpdsbfuGdPIp+CCBCUaEcz5hRG0e75OO5NoPL48HrYuFKADoF
2MDbySG/01YSFsKVW1B/Ama9zEZAFLlHI36Rr66tYyWi30tzE2+YA6//4kKslgH6ciZ9yoECvWv0
Cbdbqlre80CRo71rTwPrHDYuobp/Wlw2Xtg2WofIj7oclVzp54D2ZI30Phz0EbCQ0N6jnd0gU95q
frkmPG0tQwWFRHMBNm1aM17BC9gK0TYS7SOEngqv+CCjnilk97Z7r6MDEI6e6Ll00rkoJBMV7XgR
3S90KZDd4wPEBcpkm4WcPGzx1jV5dkZ88TFfQHk8sX6ROEqGBMhEvUONxCJm71ni94IUkOks44RV
FMdWaJyoxCXditHJiyXcCyjwPPVYyX7GllxOdKewcGEY2SHFPUu4sTF+6Sy69NRmswBw5RRjOfA0
I+YnleONfUo7TxDGkyBq5tGmSmRWuh1PnyGlWnTEZWQ45Rax53d2WR+PQ/W41TEk1HaZV/JUJvjc
Vo3u6BFxN+w+E4wDHCwZCbXpfDL5ZhEEwL0iRTA5qhvfVhWbMqTIyWbUnuJ5VfI788xN8XbauJtp
h8tOjUZK5pjj5AuKMmo0VXKUEF1GXqvmiKSD+/VjBA41uVMUzkBgsVAk8VFqqgglKp7o/YarzOjl
v+dNgBdOejpHUH0lyBECW0pjZv3p76k4dvzcPTm/L1OqVdxRE82ElxnGW+WBmlyzeE1e/KAuXbvK
BdHCYftQnpktILTo34LNwQw03bRvSckayof/+55gJtqRT7MwEGo2lGlWdRAHZBTjYoMGkdEUUcZV
BY/m53HP/Jj1CNU/Xsbuiq3n4JjsRhcIq6J1QaRTuXvGzjqk41Bd/L4AxvaNjYY/0t4yK1/qehEv
nHGBoqAR5krp730rlBFs48s2WEGrOUW6k3GMaAz6mmMUnHyb9rzJ9ty7m2fltDFKq36IJmviYlBe
bYqSCFPeXsOppMf950OhxNDtMCHo7GcKFcdGS4oXbHcqoGGMTypYDy5L9jF9cjCKXYWLRRd2fruq
J/xxz1QbC0Tha1kAvge9qbhEzUO4lHxgTLF3856ln+tHx0CNIaebmgnl08dh+KbKgy9xbdRIuiBB
vcuGH1szimqJZaGvZwi/KcICJM7XPKHW5bHQb/voEdrMcR0KOaAT+Bf+t7gvdS21f8FHFlBidKYr
uiJ75bkKHQmhArGbGrI4F2AExxg0UmLmOcdYEMBHEJgzvY20mX9X3qI6rxlc+RL+h5YqAtMV1GFZ
yPGBVusBHpYuXPjasUHnEingdUg8YDVzUfSS3jBTGZuy/uXo5qbdqMSI4Q7EI4VNM7efS3vZ0HLS
yJhnWZ5baxyO1mSIG2/T1+g/FNPioYXLbzvPPpBU3f9Yvrrrz8+PuOUpPMiiLIVfb6lwmrdyHAFI
S9j77LERu45r5M9h2ueu25gGiLFmel9wbji0gXITiIoitvMRidiqssCsRGcRZYmSw271xKhd5cBw
XtwHE2iHxNGqPRc2hA/pQgr/6ZG9IYbZuhAImfpyXrYb3SAmfzMXpB1GxrfaPQKot766p/HiYwhE
jmZJjXS6jXiT55S2tnXTurANl/k7CP0dlO/PlhjgV11wlI30uiRH4sBFWyt+WJCAUKLbifDWJGXC
SfO7r7Kx+HXO4XMNOz1XKG+sX/14Sdpve8zfyW17UdgTRgHU/p2AmLLu0EN1mH+S1aFwOj+SmXx3
eCnPzmaAt92AIiqbskseh4PFxkxKJr/qnDBxXMWzmfWAIGM5jXDeL0QbdRN64IyDi2ClHMCMwFtY
pU/Er1LKn03TjSxn6h6YtowRWO4uK6FSruPp79JAiZVE81vyDp8zQhWEfjTENvSvuT3IXz0dgXiB
Z4kw3MIF3wAxxc9ySCD492gvcBEQlryneopXncr5fRBYnPSnoWmh4wjtIWbLTu5OWlv33Hmd4Tjq
OK0LYWSG3zkVM3qTels6YSD7y4NQsAEkkzJUqNar4+DwHo0h5JT2E6J1ChVjfpRx4kZQ2YNzlAPR
+yay0o9JLtHQmbqHfTOr6Nl1A7j6Svh1cuOJrk0qJMtD59DtobkVI+No6pQwuZAeqpPPOOEZj1og
quVwI7tZ2ARzn0OYroH1hraKEAA4KBZf04yDIBtbMeE/BQpn5Vjei1kWYNdaMcF7mF/oEQk5XnLm
EDUOB2/7Io2EiZIK8bsoqamWMc69bhd0RqaAu4HQPlfspNEm+tqJBNNhCz3XKHDailnvUVrHLtAt
aoPhEIximoDHZXUqryxTYvfqw2UUJhfq756TfTMFvBFbiwn9FUsfF3tN2kzRkYetMtE4mY5VPQrK
FKFSeCYa3cdLFS4YvEGs/0YSoztTIlNKi8mETIlmZ5wmtoSip/hreT5rEb4AqknsWzTp3ShD8YOp
NICT7Uwf2z8jXqmjwmMahOOv5xo366vUuPbMb9ZrnudmDoamwa9gWekuSffkg0/rS8U+1aQRprPV
Nft9aB/7D8H7ka56Jk3FmCI7pSq2dJdpWJNo0SmSKPjlAu7JbMZ/V8fLP8NX4ors0r6wH/yfmE4O
w/FRrYLMZ2ulbkB02p9ErxUb5uU78erE2Tx4BSkelTY/JZgUCkgbI04ubKzOHIhXX4781LB0jbbi
xLe/akvt3x/4wefkv3NIk/Ken1j9RIUmhWyFErhA3yPybbaIiRrEfQorRi9Hx3lMlMzrOePS31a0
RJW0DFaqp83rQVwPH6zCrvGGIrZhk6H/HbfEyAem0okted7UqVzzZ3Ts6xWx4tLgPmsCd/XWi/WH
kUEM0RyR/6MaQoJ+mWjOMTT7tR3ae/0AJoErFqJUs5SyNVSrvWFImMOMPdIx5FwpUGwUgvQ8a8zb
3+4liDmblEU22qkAxT2OsDN2gAveAuFlZT3J2kOuMNp62PrqqqCZgo0RjW3JX1RwBeKnUvaDo/mq
Cqm+aG7fTcxMcd7AnJg3v3SBBjLv/sECe0qAmJY3Z/Iy8s3zRTk4bIzMVW6YlY66qiYRGEGAy5er
dcgT7OTxdMlZctOH+uEW/nk9dU5Dhjmu9iGBDKR6HNb2ZXv+bWv+6L5cl2gS+qSpLa3+jEgU0bkY
LaiRBjMUTtqShw5hA5G3YamgTDDcW0b7Eoo1rH88IRu+gFXT8j2ool7q+6jyBHYmC1qniQsT9Gw9
yEMjUoTDnMrOa5B6Itt1jljWLFDPGTaI6694zLI1KK6YrRsHKxnpe5dyeRRNQDeh4bqwknNJqu9Q
nev79yTUm01gX3qMmRwtBs04RflxzXi1dUEcWbpEF7DHZ9PLuEziuBqV+jat06U7n7gDGAwbo9Mg
yJifWCQjxUyL2tYw3LstULvY/sZ2jF+kLSJCl/jUblSBGXtciRz0N8BRdK4BswraQt1u5rfB8AKW
iyL/yw+Bnoqk1tKr/ydTsolA3/ANmOOgpTrmpvzZ9+07rCU6QT3cVLeSZO308Id8tDTF0AIW/iWO
kqB1+X76y4vf9S+YoEw+jJYzkwXaQG8MCoCehXhP28hwqAnyEXE4apf+FmIVzSF+Xnb8YG14+58s
E8AZcx9TElfIoANLootstR9VLzTHvQkMOnTpDOwE4AZIJ920zJ2st7HV5gvm6/VulbwlH92B2mDA
ObRlm7wwcA3Dkt3R4AuzZwljvusMCPIFDoMC9JbmIRL+SZczXO5N0Vxt2AB8qkuYJ5hwfh9SK6mS
HB/WhKZezw0zYyoJUjOa90A0OHR8h8iZzb7zIqGmvAVXtibQ2P8HEJ7uCummE4IVg1JRNSl5PBE4
xcWcBytsgLemv8m5pidweMv2TpHARrh2dWDUfZW0hK3Ry3+dOzyGaccgGDcQqEQquW4ODQOxf6d8
1tyv1uBOhS/AX5e+fHWgqsBkeQ0C3v7Ums2dRco5bRX2SqZ0p3XZzVzWu7bdq0Ygd9pqw++AFtCu
TEXsykd7NXY+qPwJmyvoCXHNjf7QHsBsAGNiffNqA0QOJr+nirwmCbRPI2+xdbV326dZ8Ytr5Qje
NlaLJBPmLGHNBMMe832WSDrdyCTLYB6NbMKfGHc7qXl7Wx4b+LZCAWO173jQe78XDD+qcRUn2+h/
L1TbFGa281UNgjsnaGfh5oz93Y5Kp8dNXU1of7aGDlKM3Gv0LdcnZ1jQDovQnMMeaVdSVf2nar+J
Ene4o2926hdupIqYszgIheCSpH1f4lVLjDGLbZdNhEO9F3ULx5i3d+Z1jaqAQlcicIv7P6DsK4NO
ZPlmFzUP2IRe2AyPb0LQsvESUoHTPaNhqE/faViIWBxSH0kYHetbG0ZPGGLU23PpOEukBFZUux/Z
APgCnUeJ29bow9HwKYMywKnjpjPhkWo0r9a1OmFP0zZf3NAHxVqbAXImfT1yPpuCgvwYQPROEhD4
xtY9NUqpL67FjJlHJZUucJ2XGxNhK51QCx2JV7VRX/3Wj8yPixuKzPSHxlJ/jx9/4F4l2EAC+Blj
AWiCvomZEADK7ebpyZjBDJOezbgvti/6/Fde8jsVlTiG/YbiA4aRJps2ANPOk6DJEsPypcX/4gJ6
jnE24sBt9PVYJjiik/i+DCON0cJHy6SnDK/n+B93Qy8n0z3Ty+4f0uj4sh+9zcA3+v8cXZerLlk0
ykftJC3bHdarSTZ5+s8O1wGHIyYQhXmEHTwa1whh6C8SKECNJN/9dVxV0bzxrQUVpsb4MQhHA8wC
BnVxf74K+56NVXZVOJCfZV8iK/QrhL+rzWyfzcQ61QlfF+4jPVuhwd/qmDb9bXPFM+pLCyxuUSnL
g6QGEvLddJYqD/e6G7BC+OEIQQjsVSJb9Rd1s3PpKUXc4iSowLQ8rbcuaPvBuJ3PbNs/IfryO9f+
WSe9SMP6t3ONAl79hXCJV7ObPxOj70NfVxH29KlQhmsK81dBv0dlo5of2mIvMmJkp7Jkfmu5WaaB
Dj2fCh/iF3xN9XfPpYslh5SUE+rIMcscN880jzaGzwQq/wwzLMpHfOillRa0DmqGuKfqGewDxHZS
vMplnf3KAdXXsa0eekTrC7p15U+aOpXznMF9gPqICLbO0JO9tusRRrcnBCSYBmADcgTW9UdE4THW
OFpSAScluPdwjqGW93PYNvbSwoUQdsL4oVMOHRqnlqpF0Vazy54sDNGuBUZYda9W4nZaSBfVX5/e
laz8Jx14/fGvhYpb5sA72UakePxW9gl3EQ7qcRE8MQi9MohW3soHyZJvHr9akhqDYaibh66HCabo
SV5YVq94xc95YKQQ2EWWKuWTSzxe9dePdvMvD3b7eBcVPT29mCEWi8io34HXgsdWUHs8MBfmJT0p
3WPz1aP1GxJeWpyHaDetEbiJpnss9JD/zeTres6eW/oAEe4ThT8gejIYLIpMBwf/lWCU3GRjZyyX
A78sm39smph0LQArHHgMUFi2BMaB0WbA2WfzgB4awqFWZbAuR8WHL9y4F+fEmC7eMEvcRq0eul0V
7ibFcw5VbNtJOAH1LU/PP8Vwwbagb7eECRN6xW8CUbUzrqOKT5fk5+fpYyi4XZJQWg2wjatbPzbN
SP/TvU4z4pxg3UGTheqOT+tGvd4HrXG82kHpDSFccs7EpcKh4HKzcFPwynrPnrBhSKiqmxohKLp4
lYjkwITWdQ4esAthoXjJNmQVDT6sZ+kERmESHSYy1ln/oStoRE9J+/2OJ97migbrYQKaKJan7edh
CrUzfQqrXMBHHVTdX3Txnh7T2d4yDn+27kHYWmv3sJAgC8caAzwqLmn+pdGrGa3Ry0qjlQDkgfEM
KaPsssaPJhfBm2ctvBRt3GE0X8mR7CnrbeKQaLWQp2MV+5sjcjV4dOvyY1lZPnC0hiXR5S8U/wMk
cfdTMj+svfsTOeFRDGMg1UXSjN4Pboh/9R0NdcRKjVhz8YII/0nDsA7d0oFM1fwL4w2djIHfVSbJ
e/Js1gGcfnIPMs06BdjRNaCQ0+XWyDJbWHMLYHmVImB5o8hr8zbKGScb6N4WhwbLw9O+FYwOEdGT
fnP4yISMEImew1cU1AMNVgxf/qhWBSGN324SjrRVrKet2H3QQR51UHghhTSkJPQcW8hE3dd4bwB/
e7fWdBO6kvPicLZ5eVmR8CXts76N6WItsyIjAg9T188sHi8sPsB62XFthtt+3sDELaEsPz8ihMf1
fZGM9IX1UcmVn/ff6PLAGQxlnEQIXiuMNbRrLzSq1JgCEr8+V1MEfWiHZFWdd+nL8AcgOX2ndicB
zAfrtZyywFeMHbCeK/Hd8O0Kldln0oqiFD/0rfX0zNJ4BfewGYi33bXyrHTmSkPcDfYScCJGynvC
+REkOmyz3P7LFISQa4Ix8lEcPxb5XCTEQUlemGO2ZpRVDBc/ryFfRpek+HgNtDMWQPLGYqecZn+d
Q80XH4ffbfVlUSN28nJL9JltxA9gWMbgBIwOHfnlhQNV/2wOKc8G7p6684hBtc70UBo8KLbBJ3ED
nxpVic41YsRO4nZrS2b7cZmdjCw0k+cOAAlEzzcXjpRWWSMMcntHsSYRpjD37+fk0wx/BjQ2ekyx
M9Go+anaTtXl3dL3ZY89/ExK5Us4VhtR1GcINgl2fLk1dXDfiRdYzPUauTLxOxgqpV6yjpBjMIfP
6Xob3ALRRuTID1XSoByST8V/YmQe5kBIfZ5lw7lgOvlFlP0AxQGAVZA+2cfRtdIdKkH62mwhKI0J
K18lwEGLN/WAgykiDvahb9A/hQ9ivuKWNkvycJ1hOz0yf4IRlRlXKabpXz+EweAFy1sk0JOCU1BO
zmm7NtdLfB6gJJY7cNtamJSCr84s3IY1YMius7pvIRHqkp4ffSBhgq677rtgqfQ+v6RH1PH6x8BB
s8doW4m9SXXMLAgSedwmBfympjoIdJQ72NvtCQRRNzo4j9Hg+gt5ColQ9jvjUXAYONy5r46jxQCJ
+E+DMJEIt/EMYYw+mYg7q0ttegVojiiXGzrz/tohfKO5+UJ0F//jnsiJNb57CnjRWK+Pqmomkl/Z
8pX+pUlPK39IQwtTBZciJ4uBDhwngMgulkokDogJ6OeE5GHDwwZm0/DeRjvePZcXoCZfXg+yNfto
5PAUaaJiSBsCgQuYtHcXnSicBN5azjoHk9YFbZLfceJw/MNg/mqaAxiBB9BRwk6HUbvk5+hl9Pxp
kxS1eRck4EmAWbztOWbfRfzsYdMnRq/5VkuRjWoBaeAfSA+R96XZMH+GsiWhu5AtRfgiG8LlupsA
Xdfi3l0iaZ7IeMBiAm/FUS8ovCGHY+F0R/DJ49zVtO6QG/V8l0X24jN6Q6sq6yKNOESWHi8NYaDv
Mi/TDpBhAm0BzFC7DQ53y9Z0aR7jWaoL/8a3jXqNJLilWlloZW+L/4mCjFdm4/0J6CQZNWbmVxvU
VPoWdBQwLxTLXRm3wjprDvzgBfsnv5cDfiaC+35JWvolmvZ/Iwl+k8nqUJDLiizBdup/WtaxBaKs
1lJQadUsue/sQ9CiuLuZ52JtU++S7SyB6tZyOlQeF3Y0g0wIjPYbZ2/u12X0Txd80pMeMsm2scgX
TDDCyqhYYOUIh0Ug8OsulafzVu+qbIOBIZYI4NCttCNxdOtPwvg/ze7ySDnJf8qbfl7uDjjxuVCz
dTKGL4etESNQqmqgvUz9PSSoGGPzDH+rWzkuqhxwwsi7dRmoSJ8cpOxestFMRtZnyNSNtVk0Q6Lc
UHe48dPmu9SsiNQjWpyah8oDKK4Y8T7K34KiTX/baPq4PWhJaw+w5zZ0d3oJyfmuQXj0oSEh+1qY
m8ud05kh7RG3zk0QyOd/DJ1H9g8OXBNp3wAlw1o7u1/zw1ivViQvLMZq85bvWyH6F5BK5mssqc9c
UjSl4yhCeplzBNUcpkpMYka4iXh5h3VAPtTTEZGn/G/y9BH1kPOxo1dzg8w8Lmulo5Gf6FSRPygk
dlX06Ui1mzzfULcMIojwxBXJge7vXdIQ4VmXycrBwTJzWjBMQ1m6VIf8OakL024YTX7HmqXfbu3p
cUCrjgv2a5g/8Dj2+PdJfmI3Dn251xNRJi8zjzk43yMegUQaFIqZKTo2eQ0ofiQ6wE9ztlQw34Mv
wfl41JS+C6g2D5NN9fj9HsVfxrr9TfI3U342cwLqj+hImytXa8unsbXOFH2ZOlLB3BL6mQdTqeix
ad9gj23lG9d0JAa/9nXoZlcCTe8RqgbZOWec3JBopYllQ4SL9shFO6tDtrG/0joise9vaO3YYtqk
7hHyezfQeYAAaln3c0KZg5cxGqr7Nv/RvbMIqcxE5EpLMj8WuJy0ntJ480z6THZ8whyOxGu2fSvj
DyPFI6JnGg5vdsMwmwpppNai0QQuc11cld466CD81KChaW/jphPPy7r3JqvvvgQB/ZOL43rp5wjb
22gnv71pJiOF3aVEEXWzVVMquVxCDKhdQZWOZ6HOk7mFzFqf2BzjM/sFbMTQKAaa2w5gqEueRcqm
3x8nqjU4WjFz+eWglpcAoQswyY3cuH46fIy5TC56TXRegbN/N4QMnpHdbwWUeMLocxTlO+zOmsgq
Bl9o9dnevWZfSfk0wwL2WmMiQcLKUHRhgo+/M82ifsHlETNhUvllcMisby+bErGLb9O/be4ewah6
IyJ9twmKNkl3Pxlug1nASCt7Ek4J3kJ4WkfGCOn3gQGF2RLQ8Lf+VaAOTZ4mqo4otTalszQmv3BW
uiHdILMj3PZ4vB4Zlt0BiYDj1WRpCUgLrSHFRNS5dUwpmSSZaSZ6H9K7Z+1cZI0FL41AIw93Dgbe
iuq5+eGPF7Eyd1atR+9SpuFEaRmfavWdTWP8WP7csRYRlxe9TwAI6leuPy9gixOqb6EHKhGMTFYp
DYjaOhiTn0qgayJ4BOW6jTzln6Ey9VmzzIKKG9/dSOh1Nwxkpzm573aleAuksCV3mmufDj3kFD1/
IhrGOco5FHm5Q9WhigAF5WLlE9oNGO/227L5KfdnEDfNV5/QLldEvz/jEvXahMSWbr2HjL5RU1hG
2Td79epd/e65NFnqharunTWE/Zgs3sjB8ByWiOZq3+gkopJom9p1P7J7msHyr3/5ZxozzeyDfrS4
OT/6S0s5Ksf+REXHu7gahf3P0RL2/udO1hfNlOoYQM0vCXwtNWb70eBJpaVxWzL6Z7857vAPboZF
ZV6LGj1PAcsI4acIh3CIJW7CY+ZJthyU5hl6f2fqZp+ImINUfUkJiz/8gO7yc1ES0fOa5Oo/8oog
z9N448p5Xe1sN/fBDvPO0dLqZCnB02syQOeXUn9cDcfH9Hv6ZFw1DAtPC9DVlgsc8ycRmMfc+Htg
Vd5VLFyU7y2DguywbpeGMeLy2Vsv5P6xzrBDFsOmF0R9uggPGgBckHboZ5vW5WdqEIwruwe+awDJ
ypJmQtOEX9gGQF1cgBLR/2izp0t7V9TyvAZrcVT/ztNEzN0IVtIV/v9yJfcoXecfs+5etGBAGQf6
Gd64e3D0Af+jWcWndRSF2RU8f4GdUgchz3o/3AlrXXYSSw9waYZWGY/wO0ZNFKXXOdikwCUmvMKn
ubMqNfdtA3WFHEmK0nmv3/vwR34aSInOkGVSF+jCXh0cL9wR+obJDlRBqMD2pYtTXXOznQ5N9fIX
znVrRFkNVPMdTxgNiCYWfRgwnA8xFW0t4JGJkdDK8LYHjg9jdzDwgFRI7xNyfoZ4NBuLwW+r20PO
0EdeGa8XHjkFpw2EypDr9cwIwMYyXqrRxfh81UC0uUaXhM7LUTor0d2BXocVeupb+jjN5Fc/p5Et
qdmU0BP27mjw6cIFZ0ArUKDUPOjoor+V4BD2ya7F3aDXfg79fLnOYbJGo4f++537yl+x3ztu3JtF
MDkEU2lV+ZxsXORDzpoO7WKfzSHtOgC/rCVGdDMh28EHamNZGLXSnInXrDE2WRSF9PrEjEUknHv4
2X/JhAD4sS/ttHy5VDIGrf4HA9yGP2i26ObY9HkkBAJYiDOCz/KFClgnoDqF9LFEMgSdXX378t4f
bAZf2WT8PgkxKC2I8I900uIltBmwKDsi0Lss6EVVs+1BJTkeqVfltlJ3FtS53/PnsmZbR1lKF61+
5UCoVVCzNVRfo/wIx1pKFWt/gtCvdiLDhrb4g6dahXdXrZtLigdt3j2bylenFqbD/lVpXeRg907r
4WF9tY1wn1f6Fa30zdciu7EM4BHMHLSCkZk99N8Cx+nc5MI6MydzbDE35+nISkRmGQS/b8nC9Yt9
wEPdKUo2sPlnuWABE588LwdQoBGfwhgKnZqn/vHQ5XJXH1KfOtJt67WQYoICUkgcwo6C4Q0FCX6D
bYiKhH7pBV9FDUO0El8fCKxDdKIV8U+2DzfnxMSKG1BUUoL+1NEvlvJfLZ+MVoCSJutkThEKi1+q
SJCIR8GpTOx+bVzLPMf+3fOa1w+wRaLa8wQKrbc7cC8pgbAo26OiT4wzTMZXACRtDFcUTS20ZjmS
komdyqF/mnZvIWmIaDIAKq3z5DC+7kQYmyBP5fn7PFAbHCxXN9yz2CUldYv2/AWuT2WwqRTVECZZ
XbbeCUgw7WjEyzQ2kmq0frt011FyIEvVMWmv0CwDu8ZDvDihgqMb9HXV7FqCRvnqKnyiMrvbWqPh
/raGFxGDTh1Mu/Z4CJRwIuchgHzgJh3HumvsZJ+Uw0t0y4+g1rrKDkFKeCxt9DEpjwjJdSaRhgk5
Fxz+59NnVLmKnxNPGxe+2Fif3zjOWBFORfPm2pMjeGZKXmDU6cfVZ4F5MBym32r2sh+mXvYz7c0w
VQY2T83n6K/mnLwBU5RbXmknHgX31q1cD10gAR08ROmoYWzCVKSaOZ0LFsKy39jtmf0CZ4urIeGX
JJ6dRvtL5hQ9pMFJ0khD1+pvxhppHhbZ6WTXVjY4ojJ/KfwZpK6IsX+rDTTzpaeo6Rp6xZOQRRqD
5jOIEZGHEsZERoVVPcUz9FhWopXWnYhajt5M5fstKYsYDuM1ZiwV7v+P8L4GkxtfCYZiLj4ABvKs
dJuqn/wKOui5ElCLgU4BSJcyNjWcxQGwjEUJS9X0JG0N39EvTj0048ID1mPoGm3lAwN0RFtlauLl
ntR8pHwi92ko0L54IDg0W5LTDgwjgqTyp/a29ih5rsMgsIVoB4bT3VUKwGtwBHg2X+34fxK75zCv
a3AeMe3dztcdenKkf52Zvkr8fznmyB+i4US7EJibTes9GJmU3SF+eVIkMtlcrQQ0zMS1S27Eap0T
/OGYfnQ4s6E4fWExM/Od1ivefKxChQK37359QkMgfljTa27kq/WXAehFJDolOy3CoPJNzHGHLVnR
rSKpg+jO2dos73abVWKQl7IO6+iDXDt1IBLOnifSIlPMHHTggHOIQs8vXSN6Q1cZIGqme5CcHjkY
Oqane5IkULhSk/eed/tJWvXX+rAHuNviHFc2Rj9SV1ke4KCuVFFRfmcu3kwUydQadr/AuzWBMuGb
Fr4Yxs+IRqXbkZFxSKzqhKkq/UZzHACeyaH1h3TD4r0DixWNQxDVdnQH6/AMTSe8Bo+B0a0NTi7M
tjMJIkmEwLCq9d3cq6Nu5mli7nCuCdFjed5MCvaUrCm4OdI5WYOrARsI0tix6Wam/dFhJ4RqCIXl
hBHqzTp63nakvbLvcELF0/Id1RQ9C6zTXbczItumNpEEpEwco0XSO7EBuCfdqsypUspVYNKWusLS
e8PFmrrdj6JU1VDq1s7epmpBs+NU1CQwW7pCpPoGObBpOySblDZJ5cCYjELVschl4T177ntqzgN0
i975mkITro6unAktbgCbXk+Pp4w9GhvaG82IGedKBGCVaxTZugkw15uSbKqRkZho5vyjWZ3d/dLs
K7Ow0MACej6IaUKWiCG2IOFdVZQcc6aJFhEo4235PiKFlfBzXvBH1raLAo68Pit8amZjv5d3WFZc
tYpL7hWYw5JwfKpNTX9k3DFmncn3pDPTsZTOK61S06oeHkH0rEZRMN5pnc6bhJAFy6jnLATcNMjJ
4GXmhEUkkPf7fnuUrfagrksnmWeA2izmOeAT/ao6Uzkyy+ey2Y1qzuiniXA5nUhuMOXImM7a8PIi
0W3f19p/TJE6EZS5llSixU0m7wF8UoPTgPjSVzpe3HYdIrybngKRCMmIyA8vQUPhKOpjc7QW/zgs
LsJeUwTzPcWkxuGoxb5YmuDb5KJpkFDnuUTKkOd/KJeubhAU0Lb/xmqyU4E41FplWnsyyxkUpqyB
lhdbO88NIgxz5f60+/srgR65rkg51v52G2MdgFWdaal3RHlCnmoxnKeswSQh7DtP8lDsdWB2SgTL
1aoBfDLQTR20kYGn1tmuXytd4scAV40xLhQBNDa2bRPvtPH1f9AwzWKV7hsSUjMpBjw0yZmCDYlh
aT68JF5OO5lZ5Vlo++nH+3ngkhwLWtYBPXtB2BTBDYv/LGTMDBa8/8iYXOvLQuQl4/2W2Y/slgUh
U5+eO1XPNODHGz8ZkcQS5QXfi954KH7CqypiNcqlP41W70vgU+0ospbP1a3m3FDheUh/7v8G0SIw
vxkvpDOuxiUqEiqli6CTnC+kPf5b+OjlVZVWmSWyMvQ1hnGHysdYAhb/UbiZtZI5qB5cxJdhjLO/
YlsRc37oi+IUdoHzl4yirgpKhazBQ3xewIPnZKHzHuMOmjkQFi/eGlfOuso30qpFxC+BG52ZZxb+
Nay5k/xAR1z3g+kioG2ZcouLx/0gHDiaJkvGS0IDh5wWB6SlhNEjj/nO3pGQkVQbxTRb8cK8BqUF
PzR9gIpMFBRIDugLtWtTCpMmsiR7PgbYE9CSsuoTY+KScoiCrrpn2Ol+aZlvCJB6g2Q7yDKawho4
8eSdg1ZYcuicrKXUh13Pc3dKBx1wDC2Q+uIRpkW62ZUUf7LWzPszXgdVVrvIlUvEoDLIUaUSDhW4
8fBrniqeGlmfyIZMVR25wgWWLiQtXHUjGsyuhMDrD7VwbIWnT3LvcLMD/EQhrrka+Pm5BUoEx9g8
n8BO4iy2UCe9wW6+7D6j3LL3xWJhvfjcmp9cwg/odzEbQaaRF45cJjpHsX/7UR+za7H6OFHaUVKi
yozfzNmCiTfsMn/yGdDyxsTr4n1cmFv8YFRAlIgyqE+hjT/ukmmJ276U1TjO7FmpdJrhIuDrxahg
/+/rvJps4JFq3IU6VmjjtAB1ZGurAXuZnqO0vHYtxsRTkzDP5s7n32ugePm34sMJKY9p+YNS5wZr
TKzrVmbUOP8/Zdq4u79B4aAHQSx7uAWzp4G+JyeRs9CCs4auKmOWqMaRZLRtJE2crnG+bc/BEwFL
uoAVsUQP9AFt1bvHJwyPI84+3W/zzuPi3H2bPwOr4lGJwkTJwMfFAOyRjbHRqB11FVgYL+UC2iaq
v0n+TfKh/ZK0lteMmft/oJXa+1QE2zwddOMKHcivewG9e0CXscZTBS0RHKtKUZZ8h1eaFNykYI8M
sInqFXdLQNCLrHXAULN+aKbAfcTWjQdMh9T/b7VvPsG0CV4+gPOlJGTzUlbvufvz6sT65ouj8dqF
dMAxWwM5xmfCkTU4HsPbftwiZmNswGhoD4j8gc7mPmXhB+icMhrwVE+JDrL24TDYgIH7kz08C9uH
GVJRuruBCEfoWPLfYiAn7QPmE+Hh1C3+VKAfMfYVmH+KDEuop3VSuVYyKxFJ+P27AYW42r+SycuX
SLsE/o79ZFj6PmU2Dpb5M+0OaXLTY1RRWArJFOdwhrTTUHoU83AXWxk+ijGD13/BRZzUFIelzPaH
+NWD5QVcxtWUURi3pdslNbV4Ia2imKCSQVcvPr31qbMl9wNM0u1ielsCBxMaJSi9FqhLwTElSTsG
6mDz4O4r5MPl+DRNj82AhAzjUyO6W7DpXQSl1g4hOyGYZiJ8rnKU6Vwnb7MB4ub/kVpK7ul+2fKc
gWIY0JmUWmvXn6eArFnGdbNIGrwDXFPyCXEJulcyrYA66AxfskROEiJ54qrOthepVCEFKtoEQuL5
Wp5hM/58S3XK3B5WEvVVuGrpPDsyTQpJ75B2kHkuMBj1S2zLA6gUvZCzS6sWO1Bx73wGBaFaZCOj
W6n62o7teNxUWnKCkJkdNaAA47jr+pxEUQ7TTv3lCNVRQfU6vhQ/kS3p2aKOHfi8/JdFk0tjbuWJ
a/hODW2QcRGrcezUClU4OQbFppmHIuC+Nws4kf+p127eyJd1fBB92IihOtt4SJ/lqnyDdcBjfaTT
ubxKdPM+uneVa7jqZ7HkRBuYxmGK8UtgMSVKaVG6YYFQBFYgCpFyRR4A+zca1RmJhmZmdcqR0p76
A1eOqpbBdZGc9SKCZk+TYMY7uakrllAmLR8MxmJRjFJLGLy1i6ajWqVGZZlo4y0UvTMTPxrbBdxD
RdxH9xNmlmCAph53qcSQo9UvcT/BY5evtBdSogGNaEE+64dqVW2PNvuzGs8Yr7EYka0+1f6CNw+w
LZCOLK8V4OuhbrRJcvabKoIIgzoc4U9jdEaER0EpatcgH5k8BV5kX6MYqsmf49rbUonU62U3jFVc
YOi/39RGLB0zdR8Y6ekS23KaJF6WIo9mVbgMRm16QMSnN8Kirp2GIkmN7WNsEu6VOUBDRHq56d8t
m43iISJEtFkANoFopt84vwi4LNvNd0gtKdZTbqigTXRyO3/tTjcxhWQRXttNXI6zxpO4x1Ws3aKA
VU9wqDHmMy8fYnIhUx7DAjxdHAFbSj8ThgFnehBEyYcZW4BIJhpUezlTKBaa1q4l81zrtjHBjbyD
WI42UlWqUJx+cD4kiFiDn0uhnQziCpG3F0FnVzK5WLyPkQ7ZNeUaGiYi3jt/i4gRSGvktXXFyUDr
lMbg/RXHGzug6iq4pW6ir7AnMfnAG6wf0VFg8E2pkEVwDagw83m7rFr9CTrEOCmz+EqeZqlZuoIp
WY3oMMxkua4+QHBMwovv+v7v+7mjVheWdcA7KEljideKLY+w55nZ4HTqzhopwgAremJVa6zEDYB3
a9JRgsxZsITk1xKGeOrNS09+VjUfOwSvZR38ymFOw3ttPb03qwj1dAXL00QQtab85XuH7dOlfXkD
pF/A8ivtZj9iMFpg7uCAAAksU5b6i2fD0H8eMIjz1/hPgBbi97nE4GfnHq1XalSjwGTslhW5pBN4
HUCFGnX9V5IJabDXZymyhWo6vE8F/bHIBvNOl+gp38Ka0txPvKyuIHK76ssthyPEz6rRCLAXuLe+
bRO7oc6JvuQ0OMPVUNpLbBKmWhM+E0EVg+Qm8N+B3+c2JAeLPacICGRTVdFOupoFoBmTarVyXE2D
N92pYotRzRISayDe1NacyfzEyf/PlFLx94/Mlnm1Oby/0Qcctuj7B1YoXBr++95zxnw904Y/qg8M
kFg/NevMokqZoCioUPjEPpaynqhQZalW3y91cerGG4l/Rvt/D48PV875Urxv6JORfFK7MvkZWFxx
2nXulT4IPT2Xh+zcA6SwumgAcpZ08dZoJ5H0/R3a9K7F9oB8GVulgB4iIYNWnl0mF505HyeBd4U0
o84ZC7fUuQHIkNhUSdwRa/33hKZnKtV18P4pfysDBInhnG18vnUZazoeB8jSSXBnqdrtHxUCe689
8InWx+O3ByyIrMmS26Hs0hiHVxNe54hRug+JGjXsNdeS8KkKecI7uYXo2qAqfbVyCmLe87X3xdUY
aQEIKwFJywIf0he0ltdPOk2/84qcAh54FTrjhSi4JRpRVD37BnWDi4IaNU3JdlriTKCw+C48eEYC
//UCayvY6SLGCGl5uEv5w7zfoD7d+0o7VrGBZRts+Gp1V4IdGPJTCbGiX9fKCSJXT+c1pYNkAL85
hy4q3bzT5K8XDpCm/DAXKIPQX6dwM+FbZvs9HfitBIBoU6qJtPXEcxtfNwwq0h5pU2bWmFHWISLm
QaWpbSrpqTfy5I0CT5YTaCrEmlX27bnoGMa3W1gMNiQ8WvL++UqL+ftypT2nbJboYvt0p4/9oV0n
kQO75R14tLwDKnPIyBdGn0qOpZh+yQ7FKiR1KJrkwZcIGhQ2twaboaf2KVDrXpui+wk8hy45FQT7
8e+qktWKpREwqrv1L6kFdw3EjjvqA/4e/bzgcoEQtE7AZAAGhlIzCKmFhvsYJM02wyn+nA36yKGU
6vUBZ++2MjT7a5cBl0cHFTODLfU4LP0+1nel7M1bRYX5ZQFzigEKUivrA3/I8c66YPBSTqbwGy5h
E9FWcay/qodbG6FrTBPALmDX0aB6IaGSE4JSlq1J0d6tYQNGhxKfyYVOrELwNeQs2MSKE1n71Uz+
dQAysku60STipKRq9i2WZYJp37jouG3cgccWjOWIqq8dmobWyMioI2YEyORRsJUyrzJUNltgGsof
tqZA3qmNa1P8lHwd7xneXSWQEUcN8Vnby4o7AwHKEEZJait1jpWwD2H/mF1+zEAiLeCeYWvTNF9X
nptF3witFG+WanpMvSSu57Tdr2TK7ug6QyfFRDxGl5hBSN1KTc6OQ0ZoSISo3f/p+CBETXCQCS2y
Jh+/YvLux7neZIFtXQcjJoh/X+9q6O9orriewxRZwewomoMGE/b3VITxp+xmxJY0ykc/o0K6e7T8
k0CjcJ+Q3CQfE8PjfKbSg3YC2Lsyl/dWOZ2fBn7//QJp7ghfwLFVGJKgLBDq7sn+PWbZVVoLBfEr
OMBTPVcuQRW9BxpZIX6jHM+cIMCLF0j8xDimvoITOXRPhsGSJeOrziUUwFeS075apDEwMPiRaChC
8uutCoWXfcQPdvid2jzbrAFyhGnLp7YKcfn/axyUV5QEXGX7Z5cR9womT39Ktlr70UjMMHTUXlkD
nV1ZZcCEg03sB4b2DJHk/Dibgnan0UJPUic79bnRSDa8dW5swCEbNRJn4AWKmNy9U2u4eP38bWCt
FYHTjWFCF7Eq+lr4FjU5PBk4BrfZgjNs37fghBvBrXtLoFlIJhVz4tI7yZ1Qr6ZcC/C1U+nyuDh2
svzLiGKd6O9y9xHDnGs38ycFbi1HoA0V2MJdR6lAvtwz1e9JXsPdBke0Qdi1QLPnpa0TN4OyLl0i
BTvc0eMDHpUpwCvpf+qdRufN26w02qG8JjgOrZJTH67i04dH3pMFf2j/jsj9b2HW8jTIe/QrB2mM
jYeLy8tlMqbfGJtFSzAcgvmBug2qCe3vTxLTUVPvQebRsI6GdBA0NbS29ABqIaPHfiBKXV7Lkcf5
/meTcahv2pA3rTFugMp2AyPsmsiFfnSwjPuG08H7x/nrixy1acbpbBINAEvMo1KU3O9NEbsaVrMJ
+D+/KmAseCvlF3MHi7Vfo8uBp9HXlAowSy/cgoC0bPVPUnXD79nNNRCk1CkKbIfOBjGK5otfrvb6
ZTsgCmZzeelJYnQXy4oOpJNZV1+NPA3PBPSylfklYQoaEa+LD+1QbuQd4T2BfbDHMNcERnA7Pfph
nrY2l5HEBXa5Hr17Vi33jfGf0J0iuQ+7RQ+8Xs+5eDmk0Hx2LcYO9BaV++ZXBLxHHn/+UtQSfJO2
ahg5oyBPaoNL0R9KQLV6l+hJm6nn7tkbvhC+3Nliw1kDDVC6mNpOptcHbSA0eHJg0oDkSLgYKORL
EplD5ryOGio5w0Ibo1c5H9bGzWKBi4r4mVqj2UqOBOPW8eN1L4a/wrGny8euzbtE5HA+g7BIPHJK
O9jP0Ls/Ayr7V58p6TDotciS1ej98O0suuyxxZBXQZaAnzApytyeR4ygkR9gi8zXMJ0rcMK8wivC
zgPShvtaLyNdi8Er+bveb6pvPZmwQbuCL+V9113Q+0vwXXDgiULTqlZJqZZxggvmtTBJvZFfs1VP
WsWfJ9eE3m8GRQN8FIB3SR70TrX0Mq8x1nNy0I77u2NBEbcw6wvW0B9S9D5lZiR3ZKHGq96gsV6J
yyfPy6/qL1B5XlsfuWQzKCUCgRBgzGR+SRk4cDTqUcbu4Ox6aw80wPwWawudSdI6O8ZmW5oAg/tQ
HsCaauFj0lCP7nzgsykQUBxduYnstElJmdI8MHsIvocxWfddJjD3rief3v//JidmDBusHkCVlnU2
BqXh82u0/RTn2kDKAnV3VYQabD0Vg0vD/5P4RqDBLsnWZbnBNfVY+gdAhkO6MdJS6OsTt0KqD1oV
Km0BZ4vGNE7sglnwxs5w+Q7eAxFe6WnZUP+3ItmVzyrQDB5Nh6TXhWFPSKraFg4pQyWGZzA7OF8F
Cv3hSuNNmg0CxlWujmvg8h6o2sADY3VVneUDQJqfvkUcT31Gr66EPTe6wwlABosOQvwCXKvNP7Lr
9Wrhk4TuXuckrh/2ZOa8z2pgfa7YP5YAci3iEcMdTT4dSfxD/ewv+xge0GEzjxXSsT/RQOsk+VCl
9kg+pVsEYHiP+FXqdahccjRURvPAuvjrIS9JR7IBUpK3cdkMMLnHko1NGMgU3Qflhi/O4ytZdaNI
YEn1DNWXeLWPRegzWNVuVgoXNNU3LGSGi56dk5mm6ByhTYJrujclVoHlqgN4c4VWmylT+z+vR9+r
pm6hrmXzQtLmSvNKwkb8zTqRNlFchFHn6Y9mHVp0zR2j2cRNYUdCXbHJ2QMGi+oGsdgwpLRfhWxq
VW8fvlCHqMePUewupZtGWejOWUSjPn2uhIIeJ/qLTsmyz2+FdMYjQ/u5ti2J60DUXZuibpcy7oOK
DwMLWUvZcknk7FwKxyiUaqXttxqAITz4IJVT2D8E7vj2TukslmlvTUSaJZZNKAY62wO3TQ8kJBee
ZZkn4dVbtGwJlSGBB0luDWvS6s3rFizn/HCTpiMUQBcguTZkrQUU5S8ksStg6bdVHxE1PASViqTu
GMOjsZzNiTrIgAk0qBjgO++871I1QwhQJLEdy+GvtcKKHTy6zqiOQS5igByBUyWKCmcpl94iXlIB
ioAIbmtDGpEdnIlzczL4ccgXpKV9OgJrlzjvpSD+JlmCzzfpTolSo2Rza8/1+lgxyAJFPqwo672l
+UuI9sKLLSvfT3V0C/w5SzatoEiWsOwZhTh6A2c/OsTBuHFH+USQVPu25sqdXilZC7ydxxfkmXSZ
VDZclQQHXNr+22BTi3/eRA3nwZEr9aC38FPC16w9Pu6UUZvydwXetDa9gNJz66joMnFfqSShJICu
N7OygQOQzD1mykiEF3fcZ5KeJ+XsrjeFTgTMnSG4AWweLvZxUb4U6VASxdlh9wOUGpLA0xRocOQk
b4yMBivQehZ2LLaC2O/9MrCuUs0/mtTZPCDKwtRC4GY6bur+IineKeZBGAb4BXrP1Q2BoDc9q3ds
J0qlGXFLvkb9ruu+c4d56pEfKEf7RYyq/Kl7B8w+Yt6VHMZC1HPH0A3TuExRH24ybUxMdQUt/meL
eDNWVfbs+ewxQChUIsVV48dDNBCDSYujZHFG9AlChM5K8mToXcZoKblXoYvpQWYnZ+WXuWw8cMC0
AD3ClxX6VIVsQyBDslIa9bWl8s41PJiws4dnloKDOrbOzJp6avuFdW9r+Y5M7A+rfJkuPynKZd9R
cpsa8dMD4VaDKO1K34umvDkax6FREymupmPJXKNebUbLi8oYz8XiZS2Ap/+urOKUYzZ400L5pgtZ
GfwOxRT2R6PeaNHKMdccLnHxtkP0T4mdf6efcJkYtdixBPoIUN5ylvK1ZI+Z0Pzq/DHfkZeheKo9
eZEypZYTvs31S7eruk3+E52LO1uaitARHWOTYB8Dv+nu8Yg4s0ZbcxtwRCZGSa13iLlnD56gaMg2
I93WMKtyAeN58XA1NaCwTfNh8MWLxb1m9qhYh3HvssetrdssQIJa1ZlNqSs+Yg3cWaJ70v9rnGZZ
YS4bXvemG3fkFH1UKJgsWNVlblOhbJhPr+yUTxvzMbZjb+o+MtaGK9hDebJR0zd7voFp8tYp/Olb
w2F8BKrJBCrs+vqQ31L6yfHBcpnMf58N02N3ybodJNYaFlazCqbGDj67Cf+8fCVcxiHXg5OlIY6/
iJnROBt7iSzzlbJ28s+cMCWaCA68+7qdjZqDHa08l5MMA69XfEtToeg80uEibEvgYVYN7MC7bX4o
UKJz9fIexDgon9vkzgnnIZ0I6HUAWsGelfSGwdK/kssEVPJ72+atVMAR+3Sru3FqA3XgPG1YBQPp
0x0Z/OamXgVnskqJDbMzw50j9SKnxSqAOb2UT2C3zx1QsHfTz+awzciRaT6boxB/c5CfV1dAaw8q
fwTV0XbdFQkERXfJCOO9TQ2DgS/lkGXI8DAkZenddZvVkX9AYkf7fBAK20oL9xwiJlmuZbP1v5c7
xf4pKsaMyh+rxvQZ2WaS6Wd7eEesgaxUqXU07DErFRdNoMBt914lL0e4hC+V88/jDHrGy3SD8fxR
HSmQOBjh+58EO3/Eubn4cSSFLya4uoFfSaiaQHvjT6QfNTI+QkiYvGyZjJ97zSiaagWUEMLyxhG3
CbAD8Uffdet4cdhim2OgxEowM0/2v1x81Wqz6srtlDqx90cI7OwLeb9MDutmr12j1tQ8TpXCa7Yu
oIEW7dGDEt8cqMh9taQLeioJOJZXYvW0yrZMNUtK/M7pKRvfZHg8Yyr3HGpVyaKcsXJ76d8dLzBa
6V+lpYxOcWVPP9g/2AuKUt3YHKQ3Dk1/e0nH1RUivtlw2hqEF9xhPan29+qCXUDo7SPXktLQQ2A/
RYkuSgHhoIGoUAefxm+PHFrDGed6SwSAISrJW5yectSdAlYQyQ2FLNZIRvcl3ipKBbQfRXPPnJra
b5X8vraHPhNcCXg6lehvjtD2TDhqD5qHBiwOaZIHjohyN6PnGKprNpKFpBOzsEvcK3wD4jndaJJb
+uBhx+deEOwR07krFpkP8o7K0UikR9qidhcAJxV36pzaDF0p6NAf1nAwmAXpBEaENbJUxPSFYN00
0D+wHCIEMQv52MWqjgyNPqnZ7DsZ8//xMIGuOE50YOJfXVP0OYNt+2zJzMSe8NBdkFfNj22ptdvD
3YcW9RBtHWELuoZSeVNtHdWOKaJUV7P98LkZSmg9oC3yrq5k54s4ZtkoBSDV3ZFa+ppNgNahRsYm
uTlTNuAfwCugvGg2+UtYUmMDysGlblNudyNdAPN1Fqxt2x25rsBcgeQpI9Uwp9iegv0FRhxzhkQv
IdpXPPxqZ3x4gdLV4F0QTmZzjnW+XYuQTZccxkstgW3S5CxC5v92xmhq3cuxXAWdGnyWW0ncmUHc
2nO2bMSWAHX2ywqs5O73xkxYHlVKr/7LjhWddUrJyCVR4t8BmKI4BZDG8AyXXAFQCewmOWQ1CPQl
7RnTI3vNFgUdHSLvSjfWsQyYey8A5Q/nuO1CY8aKzRriIrvBYndyEviie/34ypbYMEft6Pef5h3M
2lQ1AyUGIyhNISNIIf8r1Qf0Va4QwVsNrQbMVJ4ESS6HBpBPk+ZEA+8fSNYo9yUNfEent0U+qdz6
acgd+l3vVxqWuVRuaBv4YrbWEIaW1s9FQKGL8Ytw+4JHSQeYxoSdYa3fGe4+kZMfiRKsrYDBNjht
cq72RtCCDFQi/VjLy4rultj1lmGEiykXdivb9MRzsi4rVfivVyVq93eiQaj+rVVQ2Bpsf1BYXhdx
t44tTT/0y9Ey+yoL5mWablcl4hGMf6tIZblBw5TUpS1dl6Ogs0dbGGgqp4nqZoX+lwgC4JZkFHBM
l8aOB4JFzBqfS0RQxBdNqN1EqEF57uwZsyrb7zIcEz/JwpE8XDR4yaFmlJoN6hjTyaridHkSUUMt
Th2V7g/olwETrtz5dr7ooXM5kN3uxYZ1xfcNERPCUYglebcx9XC1Kb87m715jt99qUuhzRzEqaLh
AORpYg3NJIQBqqvqgL8OtNpB18j2CAm3b/f6TC+/jlBRy6B87ncnF9pLppxofry2uC45tNIJD+eF
yirPU84DAQ/qpn0CF+RA6cDDVtK/u/xf+VEvE2URFygbz3JcQG1cuIJM4gdPzyqOojo2dGMteA0V
EQv+t5W4uEv0bGDVt2tT6n8PQdLLiuKFaFCZzTav072o4W2gK+h0TnZZdjev7NmeKNDyOwVabNqS
tWBeLQdOxaVdbe69N1cvxP23x7R7ysYlPabkIQkM0eTWsXTVnZe1/8sXkOdD+xH+841rLG1SnHj0
kdqgnrOv4jahS2dDqTA2zibNbqq8Ezw9hEFqomdWakH/BL3YdabJPisMJ8tgNY4ZncI+DRzWxTvZ
2IsbMDdoW5Q6VWtuiZBSmz54UcR+a+jywM0ciam7tRL6AWAsFoXufg2dKATy//mhhjZDSKf+uGMn
XqKnXXOCYPpXAYf4Z65rTgVLNMl6yve/k2v3pzkfbn1jsar4G1JAoBhHPPkeFqYKn2WT6It4k8Al
QaI21itZ/Tnbu71yZen6/4ExvbYrPNX2FZIaUyygjSxLCRX7/ao20gY2GSLF/HSG2nGmIVDHyH9b
zHr1P8mr4ZxpmSu+kZyYDDL8bfb86O0QtUbD8eQCuA7XMO1XZMoJD3RIK41PRq91a2mHyIIx08RQ
YVCJTUjL8EGZ8QbhBzR41X8MmK0My7g26F5kjm2bS4egTZv1304V6yUIwCkn7exdRgQ54VgksvJw
CUoKTEnTnzDpodT/xbz3rDATk2u3ldtxSDWcTLd16zgH9Lb8jvvFbmLRtJefdZv3tM6RA8jbN3TZ
KicBxirSht8cfSJjnpX73iW7bhzVmi4aUE92LkbQiuzH96L9HEWqS2JSthS0jDAITae4gJfdT5Tb
Bvp6WgEAGbaCYNCelk88bEpuyFifvZCWLVEClCVWI3I7vDAvFECV/bc8UN6s8AZQd8oOi84actTx
4bGEaZWD1rBtOZ4nJs0ZX2v9BtzsAJ1PVKLNio6J7eWcqg1hi0MNBR6hJx0EQADF9Crqvc6sNHW9
8mn035bsN5Ataa7HHnW5K2Vb8k28THpBoKyBeLMpL3COvz0qCNZEpZdsubad1CwWyf2dP7CKGt4n
NT+0MNbyya2NolVDSsXNcDohwMxln0DPK9Noz0yYAhhdae7e8LvwS1OLkfa9tWUCjMsXtMLaG8+P
3rUjV6x9zUXbpPznqvLtFzl5DXKDNHQZudBGgRoxBG1wkUXS8myiPac6cKG+5vQm5tgMOsBSh5J9
RA6XEMdry1nCDoPjJEpinwfgOcKgP0i+xD3Tu07rM1zarnsV1d0N8SDOJdnnayKT6rFRkhHi8QgF
70v+QPBJj9LkFgCkqLjtcsiiwGrrld9NelPsVLeHpISlJYX7PiM91vFf5Nq+32Yc3K8VbmgfY+91
uUAUYCka1J1NXqm5CPgR8tM9hZAUWkMZUluetcoGKqhjnDQvLHTMBBbuRLepkWiBh9DjzzFFBLPk
9okn7adg51EBF0MWLIYv7MyW+D8bNifXiiFRiiI9/ie2Wdd/up2iN6ltopIc5ZGvLFjZuInSYW4m
4lgI71LEl7+TLYl7unjqaxOQr+7GIRITOPeoJwhPbnUzJJZCeL2e1oNd+GJuAVb0onKaK1Sp0tTd
uEhemNMZMI940I9Ig04JknGNniZmaXUwyc1rHMh20bDm7jWlGVMxsRC3q599gXbE+NsalXEGPAvj
bLuGjzbiGkeWpIidNHB5xTX9GT0O6Wt14iJ4NipuTI5cJVXLcPdrwZ56D+cCKplu8+NZUDdLpKdF
rulfXtAHi+D66qGYfxugXMyvjXf14u6XsZOBaiiVkPwTEDz4gVrVTIRhfPjB9IdAO/1jTeeGt048
tO02ehURmfg6YhEW+/4qOf0lNJ57sBQd3L/pnoIEufajmv1KcqWut1cwFCfOoEr4ZYRMLBGKN24e
s7eyA74fFTZWu2HJhkpd39Oo5Gr1YcWyv0RrFSuU9mXlQUgEapd1zK+ChaBqwV2JaQVW9g7A5fV2
88qcHBEQO5+OqItqoM6nCW016U0UKbKBEalUtWLSEClaDHZhu75Ax7xpegNFClHiYE0bzDWNaNpT
cXzSKxr2vV4qGdD1/yuxha8sur3gk/XItaMmmTosKyJWKzUVtIKZkGOEQoQwUJs1iFanvc4qXYR8
8rvMCRw5gXApBEW+KNg+1FEWC6AJvV4zhZ2GXM/uUPafY32rwrraEgJ4S96iPNC3CjmW4yx8IbBS
9ktbIiGxwbqGUQ7Ri5EWaKPUp/nJBVpBv7eAjQ8EFm1xr9Slcqr+6fMyreoiXdhAxGNkgO7d/Q8V
9JLdM1hswj4tPtUvNVOR89VKQXYirMwCn/O33AJHNA1BmWmNotbPUHvig1IQj319zKmuQeJ4Rk30
vbPh/RKmTHuG9ARDEJM+lEteFW5zGRaAOHpR0CIWTSjCApGI7Tbf7rAGkVSiqSgFSlFR1vOOjsBE
tbQqbPPhbZii2bpcAFwkVBA9UG5Uek4wlyHyczDFQ5NGQt/uJN0SG9MGIgNJ3pfRx2CDqWSd3pqZ
ZIBXnugfW87/MAq0Z8Wu9NggzHXIm51vOm6H3bCz/pXRadzxiCKhx9yXJ9yTFNwp1Nakfurz9v5Z
B48hEvP1Y04tS6Dy6wLXFXfYEUXMtS30iigSmptz1YBmQoep8lSYiM+DPqpglGGdliDWOebc4AT9
x1et8iCRAUrxj81td1KDZRmfAeg7UhqMcR45buNHqL1RtdmxYvZRoaS787BRUWmnOqn5dq0D+ufa
JXmeqUQUMLETdQtwMwG+uMgJBYdsHJ3ygFYw2/iojaJlRdGgzyQLhajXmALN9WuVVgXI7x3hAnib
52XYtPO8VW/STRAsJAt+fDQYJNxNgwcezxThpwdw1Xxv1WEt05Vy6Q8ekZojpxBsJIrbKbJ7CAqb
EDG8UjNzimEgji7efNOMYTsGHtbk68yuhCrCPV4Re4nUrbNkP1oSltWQgBa109B6zzyfCsewNaa9
ohdOZqS6pSnvgcxkqxPIHDfHA+dcTvdRo+Vv2GkicVHpvZyYalA14X6nj15BEUCt3Kmq6HyHjXXd
t4JADznTW+VT4V8ucUM2H0IQmYuNe/5bT4557iAUuuurMTCl3koHENLDkSr0trQNnKXZ1INzswo5
v5hOJIHSAK5yvb4v38yanylmik7DTT7yIRsZxh94ZGR7/+DgtALo3ji00HTAJCEabbmjUsOWEZbx
keE8I0kgsYIDXr7s56IC93yxRhRWGSJtnECacIQzrfTzG4bp1gQt33WUBO7xzgU78RAGI/7hPuTX
boykyNeic6nu5wCdZn3kYBRQyyz2GeOfFzVJaYZwQ3H4H8JmpBMezeDxjjFaazUmIBr3Q2DzOi0c
TTF1PcivpzrFcEgzNHhmkSL1tucWc+DKXb+XlRnW+gM5anHOvM1j8/WHYE6h9psHh33ID7b2ewsh
uQTcKaTlnlp4w+Kk8s8lMsZw/iRzxAW+Cmu5nyl9oXi948V/H0Jy+O03eHDJVrq2oYdGayf/lNiT
E/xvMljrFuVJAu/Ut8uz/oMZLwIuCMM0CuPnwmouGpWpPs7Lm29+CGvdmB2PvBRvZGNYiNZrSJaG
ZEa88nGZSoRPHfBaBfFFLpXbksJz/Qr4DII723bzXfVv3LzNMNBspqL27QXNGP5b/ozI5PG7hbyP
cJSocg/+DAbdnJpmz/e4AF6xcUGsPS7/Dml08A7uY4Dxa6aa7vFQk+mEQjcK1V4XfqwZj+guEyhf
6bsuYajoEM6virDom9ohWhq7qJJCLUFs0p2ZPk4DQiRyLZj1wxXwS92Xd7S3qWFJV4xQ+PM3cgVU
BgDcmRPh7hKY2MKF5MPnC5/+24F0ojeR9XmoShoWpwKNi9wOBDPe4poTiA+YzZthxAxF8KxssZvC
J8Ouw/DxCl0a1ajklN5jd5hHdpvg4RwyuNsDColeFmLIHNVPMA2FUChtMIdic1NHtoqpkdPHztbn
uxlY6TCy9D919E8gAgInv3vFkXoPmAPrmRjsokR5Zw5KUcFEvyTl5Yapksx6wrB3ReXHvpJWTD+F
yCjnMwY+xEjl1LpS//wg4eY5pKGAyUc5icxQkUf2lgSRXpmge+o/jSsacHZgJZeDQsUAPGPTxfN3
mkvu1dzS/kdNBaC7b6i/tT6o6lu3LdjkHkq/mlzP9YTFrrNOBir7PS5Bsz1QKL/Md36rlUiRURWG
KTeJJXtbFP/18cdzwygksam49gIz11veDJCFOjuz92DjHKUS1LxbL4o3PsEh5H+LoYjPdsowkA03
DKBau8voWU6X6Vv5W16oUHRpWsCh7c8UaCcGLrYcg9qbJnMCf8S69jq3g3UG1nl+oo8hbPWT+I16
CrlSO7J8iUMaHEE56Tts8USbB4PCOWosjCz4NNgV2cyBn9Qgev55m7syJZxTgD5ehjFYM++n9fZw
J93DSP4P/D/zpFQwFRqTkObnGF56SwHJcacec7m1QcVMJ39gVBrv3rBz4vnnddV9Dzg4hjHs5Z5t
1YX/zQNoNAzvhuOVev1MDg6g+i357GXU58yP6uJwzd2xqisA0URdcfwIeZPTlmnngZIfrtf6o4sc
RKqtOJoGFtmkD8b/d0xidHNt88vMG8NqeRZncpzkZlZmtbMyFLHTUg82PV3vbb+58i/aqtIXb60G
YZyf4TvZjGyQUYMOzvXmq2apa6IE2x2WbVfgGlNHDktj989f8NBzO70u9rrd6yu1zxumtdClR2sK
POK9V6SY8G0e2ZHZydizWKD6Rk+MZ79njtP4pActrGb/Cw/Vheten/MD8Dzn3TQLCtP7pJwDBymN
RlGOLIsTxFHKWBKBh1gWe5WOSvrpf3qP9qTsPjq9Exajd7ZlC7K/T8yyTSuygUGIocYg3vnfU7lj
sUuF1OAJWcxuE7fKejq9hI34GCTQ0WcJpeBDs0mCEmkZCPUtR4DOzJkHccUqkhKiE8VU+FAJoiE6
EX31mKAUBG5pxi+KxoML8xxSjkzgqqchANW9SvJRl7taA+kpu7eEFTrrqBKPHXwGhRgFWjYcGru8
YK9TLtdJoW74A8bYIgIHMtMnNsuX38yY1dh/OyT5icMv/v1LpBfJc3C25x4uKz3OJUyOHFTFsGqi
cEs/6O+YGkLn6/+XoEPAks90rHxkNresuZQ5MBJ70cbepb6qo7cNvzU2rq8obyO7YrVewmojxsDw
qeYdhIQ/sc/ZUgpzn5zI7Xp+Lb2rZREzIK0wXeb9HjMbrtWiOzc6LzcZRUyupX6hbu1z/8trdK2q
hlCMM6WTqPv0f3wM6kWyN7JEuL0FRn1lR29576UC8hbdyt4prLWDOTFo9gr3a/ljMfG6Tv0DHHub
vJ2Nw2xlsYj6z6PqYq6Ji0sGnESqOUvV7ILyQ8s4tn1EGvpTYC9q5foavUJQ175vTwfBh6U4gkuq
HQHmwmCq+89/Z3nRe+i7oj9nXRyTOtaIUfINgmQVHZjim4ZJ7T5bPNv7zvzaJoXIq89HUO3KbC94
GNrWrte/3hy4Od88xfWvE9nj/4dEMeaY8BEYX5st3wqOqxmmNcnODtz1wIbwzdN49PPGMEHDrSw0
aQb86YxcS57CvAC4JLPS+lyiGtvgtW5Yq6fr9hhnD3UBr0xLtRwODN0YvF9GfO0tUCkXhmTiAYUW
tjlDBlIYyrpkAeavMhy5vj39BhGWyATQGV2TXJ+sw5hHP2NbO4pFm3mWWcyhx4gZj50eBVxjCevC
/B7Atre6deHqkG5H5ZXXewB7CiuzxNvsCMHlppU1yoJ+QjybUhuN1hxwaracTvxJZpbyO1/QSfVr
oBZUpZiPZ3ZmpQibcTx20w4aV3hZ844PqeWSQljoq3/uHUwZwuZs9ZHTln8LDbbeYCqt1/SFMC9k
V01ZwkPKse34qau/yzUNSWF+rku3dAKrPRGR/waVJCmPdI81bnIhdkH9qeDUXOwgguN8fI8OCcwc
f7ujVbCmedMPylSFdy7YLolqZ4JxZvRP1WtoYsyqd1BIVTsevySnXgQn9NGc/CAfCyF1qxxtyqNM
VXpPrsf11DbcdjLsWLrzNgxmSBYplfc1Uf4KwgPaoUQgDaZZtGw3BI74oAvrRmzab2kMcuphtmHK
L8/9X+q0yomVpOFYKb+GkiJM2rud2lJBvB2CyR8nljunwKoNQ224wj10mgKrJ6bimIUwq3LtD3ib
R4O8608QH0Bc8a4XSlO3I4aGTDniR3p0XObABCqiQYuYKdpNBs9PIBwPZq8hPhkim4Ct8TGxw4FY
cH3JbBCYd2fnkpOsg8uNLvd7wK9qMQiclvqbiTLu2GIAaceqU10lAjaTrfhtbIhh7/VGgHi3wvQO
/iYu+BmjBP8FbFVpkdyVo2j4KpfrLlAAxTf+Kcpacdo8O1EqjE2oUqwNMdnt/zbgTxWsy6a66U/U
2f+tqBp5tztndoQQAkRLq+Q1rcpp9H8X/Whzvsbw6gv8A/E6PEigbYmj7N/xONoM1RfY5p5/6hvw
zdaAmx0qImYrg/yLdOw1khADKpSisIYZukrZwZhTiustvySbotrpMI4K+2sgNyGjr28sp8ZM794n
wN3AUG2qVShw9Y87uxQTi7dZiAaS4KAyKGYyRe3R8oJYJlN9nwo4HgrIIqLO6oV+tTP2j+u0kefT
ija81XmYMNaBFa+LyVO3d3NAmUZHLfM4uonpFu1r84UPxyfwdYIC7Qn3W8133n8UBvm+jZGtUfGq
uiEfha+pZUIRRzfO0OPO2+wOVJlFae7F/IUfTHBMHw/bzxSLMv0pbYmm1lgCRXGYVyZyR5ge6Wva
naubE4l3gQl8hosOpWFXG+8GYP9uPxvbHgHcFtTggKGXRhQjw2fdViuBJn2ns656odhzt87D99Ay
Ipe7H/nALqsDAZ/w+nLJvfUOFj9eGsrxAsTCtDGiqzhAAyRTwUX4nCNYUO7E/BsRvIM0FMsBgqvd
NAfuo6Czx18aFC2EwKBEeRSFcMCCL0DKKev5a+rODVYOmVUh91S/CXQH6g+mx8KCy4pe82Kj6I+A
0UvuGFg7hZxHQzgvuoQpm4VOPL5mqAFZBD4jNvD8mEuHyJX13vcxH3P2wYcqcm6gmrxqfyR9Y1hp
s26tQOGQ/YoEp5fjTdaX7DIDGeXRhwua6C1D4XXRUOZx0MI2ElaK/SmfrpfhNjd0nryK4VFyURGp
IAYlYhpnXUnSRYexJx7fy3Q+xFwlbnRXrHvmVfF/OvFs5exVt42hoD7IO4tGBhZDUjBoss+TOEc3
Iggb28C4K52W5YhiqMLktVwC6Yare5gK6KvQNva5kup6NjXH7pZNSTss3liWIy9YUrT9TRTIDUPC
Tr5W/MSwGJPedoHLmvroSPiMs0edJYlNN077Jnswg5WpkWuN4ty/SzdgwYBWQgnLYpnk2nMLDOib
6sNrObck3AXeS9v/FoZxUEho1pOLEHI9wN87fdZB3x/7LfNjUcbp/k9gaPBbBUYBYus7aA5iUlmX
A9JeETGwuSsRiBK7r5K35CO6nC8X3NffPuxkjcB/2pMZ03EiyngdzI9ICW0JEVca88s7Py3A94jB
gLfETR1QhRHBLiiiXpwOgSfRG+pwQZuV8vKiprkKcbvXxMSG/iyk7DX+benrzbw1YZpF0D0fGIMB
hLrLd15zWGPmkTzLxYui1b2yjvC9n43VjpCHAJOQmvP05+QK78LvPTkhNSPke7tMW6hzQJO3mEvo
L5UDvAV4dlMGAFI5hHfqW+GOu8eZeJQYW/QAI93ueL90S/GZRiKoDTsRaVx8enwP+WjhZxVEYARQ
PhlX+WPFOwjdcBN5xHckK4R4DLvwrgOR3CNbmgQAoWMxJsLlqC6JXPQWl5PwHV1xMQ8UwZDGULAU
6sD84NlhEK+EdhTD8xwfBf2yBinJPu/Ql6fksrL4crv+10OMbQQPZsRQczXRhJ/P0lWRA9qxBDyi
scC38q7hidJiERSGzUUPEiSgMZEnXIBE0T5C9k1h18Obxr1tL9Bj6Fra89kX3MMpiJBoUvGjDhf2
biyOjL8A3fwR0Nr4FVPDdS3+Ql7Hu6B9MyqXh91RCp7j50gNRCdcdddlI04KHV/yaNpmDHz7vsiF
cNBoAdQztHEArBdX2x/BYsZIg2048lszwJtgty33SB+9IS0+RlRC4xtsCZwt/8l/04qojzKyYjkw
PeMyKJajzrpGw2xtXgoUGpDNg3fOIN1XAfPslcqFrDSnhpd0sBMqpbwTiYb/jVjCaWd4TZzPgiSx
Lj4c44leoA2DUD6dcIHiMGocAsfKSntKdgjC9nnjSpKZ9cCEG+bxa9ki7or+svNP8Wuhsoai1cjL
dGUgmICYpKWTWBzCfeCzrEyeuPbo+QtArUzOQyEFepkYnJUoqj6jWiZo8LNBjl+JDNyXUe7hwcH8
/00VarFOeyrsCHXQhx9qU9Hpde0zDr2uNHs5VgyfCYUgnqAg6iEKoaA36DGG2YeHIv0nOZsLCGnS
TOOgOi5IocChlBzgbyqDjDLeyf7oy/FJsrRWTDSPGg78pejAbkbzqZT5Ah8a73lNckM/+biCTeHq
roP9U/sWxeYQqAEDTYCeMdNhGL5x4jk92oJSpCOlwZp8tKGvjAL8aFd0TYrzXp79dVtoTIB1JkKh
KiJfsSzxRrCCWN9JXgRIiNHlVYX2Ri834wLGwjXFqhXr37a2bDNSKOBmeIyts3iaZCrGQRw7QoHr
zMPpnwT//9OY5yuuHj3oOe+hQQAlARxRGZ43e0MUo9cHaohe1FKKGL8cvu5K0boNoEcYqO7l6R9q
Wn+LQjvyUjg3uMTXqqkF/TIEv5lJf1o2hx09VYyPYThmiTIvgGc4zXtou/GVyaNNhoFHpShdhq+3
gTOWiL/H614PiJobe4NERe+3Hbj/+gEMxq3eHwztaJusft06vpobC7VyuUEYi6DLCvTkS2O8sdO3
ePjQeSYRiXhiwdK1LN96DdKzjbfi8MKJPUFdRTCKCxpfupMXNRHAQdq1yjlJFZCi33fgDBs4S+X8
FwfTy3Nh1Y8dzU+0Sk5asTijHKgsk6khD+C3xxWrergfhvDNpJ0Zhr4TJHA9f0IGdtisjeRqQXOC
FV2PS1vIfGDJCdlRWk1QnTrBOo7w4S49mJkNexxrVHAZK7JFov9vnih7Uz3c0oOF2zf9nVa4gRFm
TrZP6zf+GrN6I0in+q7k1OPNkbHzHvNTFK7PaCJSpMfC7HVDFa4vA1CNytPjzRklFQVmAxseB6D5
JHiaP9AuEXvBQd6pIcWPdmsvrEAgQ+pBclMStqr710dENfIpQuKnprK9d9KAk/mARSEyoYorV7zs
vSF2VIRCj127T7WtawDPnwc/D+tUF5hKiU68x3Mxs7O8bczHnfdX9lq8qTlXDhT1w2Sr/4EEHYJw
XuaQxcoxxvKQJdXjWNNVjqy3btrBtW+nu2NxpUfIEB5hYloRa9Oi/HhDxXd8J56sdMbgFaKzoX9Y
cb0T22+0368Gf9s4dmQ+S+OyoHjCLtOJXOzma3e6M0s4Lmr67l7b/gepel5CdeLMn0qxlrE5jjDx
Y8ijucf/x/PY9aJ1wVs5A3CDH893O+td0YKs2KLySqRe9ph0vNes9+v9fZFMoBJi5mwRTYO62Si3
ugxYa31WMKdcx63MLUxfYKmskhxosdtPoUmpIKgePNtSjo3JT3hz31MJ6ZW7mVqMm42HxDx40bJz
FQMJvIFqkTKQn3ZY0VY+/e6IOdHQ7a6Zbif5Q9j2jidYOrXi/W3v4ELX1XRLiaFORrO3QqozFGpM
GihN2RTo66YaYPNQ2VVP4UcRFEt/NqigsdfHyvTn37R+Wfp/Uc96kUWe/GUVSh6m/NZxcZ6h0vTI
oXfN6lbtV24XNzRGPT5YnTOGaN1jYRCr3NryZ159eh8xhc6ZiMLTtW1z16WThJUmF17HbEpVjpxY
iOgHULVRkkMlEIptREaGGEUibWl57f5et/IUezX76qEvK//JTr6vRYG/X7UdRKdPqpGe6F0/OSox
xfbcC4TP40oYtA8HLXom0IwN/9OCcC6WqDz7he2QfBL/K38BgwPQeFZPb2Otv2UKRdHq8NzlolA6
3DvcjV33jQNbC5VdRz+JvQibp9UMtMtT5Y7Pd2f71NRzT7KSEGDNmcC1Vdck/e4f5AmaYHNT9dJX
RqAGi5zF7QAlmrh9yDOlSJHI8Hu7KNz1s1qqU/jFtGSMvPuY7jkXetky++K8fJGvF5bGhqwL81K1
+Mz+ef0QRKZ7SjETYLtWLiNtCxDQUW9EkUtmFM/F5PG1GxBiYRQVV0Wq53a7nxz2bFSQDfnoa0Jy
bh6Dx34nVq/KsVqaO9D+xrFJHzH0eSK7m1nZkb8VFgDyOV0TBcusnFtxijHFi7QpBeMVWmP4KHR5
UJjt9f8Mlgzj5zmSZeRxS/t/LPLZUIh9iO5JKi52kAHs8XZVzRDeR+9ZLcrVCYF3SFyHImoNtW93
Mi541il1whSBZrsWo+knDKdrNItxu9u7n+38bOQN7yiZc8gyOQgAvr+Bca3YDMcP2lIOk9Ii/w+a
hzWh/+C/Ku3PEfu8rc/xoBa6pEi46gpEGhCvxaybO4OgDz/4du54epYQB5WDSyytp3/sN4xqueE5
Bwrixx2jeW7VO2xDmA7XOKBMxeKIT+u8r/O9L3ZBfx8uPvkZgJro1+SpR5J/UgV1XQfaXTfojIx/
un2zR6/Re9/hvzY9hvhoXJUZ8wyRu8TQ2PFcAHiN3XpgWtVpnEmfEXEtA9DA3llq69O8gEkoAT6v
KdpIkLhljDGZVQzmjYopKfpgI7aIhGewlA2Xq3YqBjn3HLKJ49gylOzfjcXMuv+vDA2YKmR4cnkH
m7BbFhdHywMUdSKYywP/87sSMpjkUKzOqm+ILkOTvLYI4KmUQl1OBxHduJvb/3LWpFCO2OPAx2Eg
clhrYrvG6vP5bub481gOExavsyuTrVPExoWrmD8VcldJIYY3p6zRizjEN8ljDdrg+psOHQ0/cejK
3owhjWr1v9jLQmwwgLPfHp5qcaBehnO7ProsUKU1L0Qq+LET4/9aimrBd8BAizutl00QJzxNO3L4
IOuHMPLm8uvOdGzcmFk1oDvgvecT8ri83oBhxfFVJGBRUPpSQHg7ECcq8JwM/kJV11oEMZh7MVhz
8Gtg62ZIOMBC0ikSA5SVARJPkUmInxxm90ri/TpUvniX+XFW9BOfTCvPZbuh7XSj4HAwtUgCBFhz
81snwoaJt43o8puDG13TK2/RG0FrrSwzye7SbJzo5p8fm2okW7EiGTktP1Vm00RcwYzXVXUq4KSp
2SYZIZRQxk84/L5s2smdTpSmRkjUT7oQnhdOd1Wb6mRZRjFAmmBgFwSWLP7d0+NzcrFai8hYuNjV
0gevFG2tEKtABer3PncG4xWxsCDoFwkp/s8zsBQ/vjaF4fd1xYe3Q6VJsJYJ2BdwTcxpkPqggw3G
BHDaeW6ZgpMS1ghCrwIp9wfIPmIovqz9hikoDAwmiu+UGo0XD9hKfil59DdY++yi+ExEUFB+GYw7
FCicvSuYzQ66TQ/LZIN8jWb/lVzO3fus41tEC4hB4KmhpD2sJydQUhli8JsJZtzdj9Fw1ROxp788
y+YPiW/QHiclk6PxFzmNqouchPHxFmRwh6t1JyqUlTzIb/4zx2pKemZSEVdaavABRufcrUHIv6n3
dRVpUc/tXnI/UYMBLO01hZ39UMDVIKxIlNBf14+yPAkJ2o4LNvWfT2Kh1qff05Np/mHZG3XYSpAf
7+6qxtHXSXaAoXQrEUGPLVBf0+QTUOtotzBmfG+FJSNz2ov8Le0esA5Xp7wbMPMYrk1OpeOwh/cF
ULA2Z/brv+uQzDr0Mj/kPQUTb9+vUuEfUb/8QFqEo5QzCRGZBjhmNMZ/71VpQ55uyafXFNPh7cNZ
2skfN1rx3rcZD7hjidEpO0c0DRBsjQtrb6b+3vGfiw9L1iJ2vqLRxLm3AJwMQl7+vPwsYSsSh7Sy
dpIZeNFQqBBb+LOBRgr5+gSFy7eKgHdNz+7W8bE6NLGZJbDop/yYy55Furi9HpIy5Lqfu8zl1NzC
Hm1SwcSVBbkFLAgyt1+UQJmKEvii50iyMkpFk9SSqlEnnzCbi6h+Et95QKFcpkY3vaIA/BS3JPGb
+o5veHHAjSkmpPV8ovdlXNeyOCyfxkPa6JzWI/rBtcGNM3KemTw7TaSSBbe5L/K1ulxXZJ8ZKEv+
pioedbg967Ewe8/4mnx41sKETnQqrbuoiiBxiiSON7aWd40wWmPK9YBJnbjcG8ryipNwYQSvZasS
JSDRzr0QnnKyiBhbMcMIancvF2AVfato272YkZmJCIIbQlPCUFmlJ0UIG+SBs2TjlITFIsyQhwND
6MQ91WY9R/kltE8YNv/lvehexo4/YyxaxOpGzsrF0ZNk10zsdt1sAjVYlJllu07aO7ivOs7O77Sz
0cZ/xH2UEWu3CE9/sl09nG8s9JptdAMnOTpaDmCAZNnpzCt/d7GQIdAt2x+BgyFNR/BeUUV67aTi
L+yT6ONWvvJ/iYFG4flBOo42Pl8XUmRkyv6i5a5lgAXdFdurqhx/6Q5LlVu0Yj1Eyej7+MV7YBY9
fNZI1vbVv/3OAG1i0BtRM9o3gVVW7jdj7qOxRju+Z6DeXkNRDPLM4r3OEhFFyWT+waPi8G9hYdvC
LllMAw4lAr+3cYNrrMJAKVKh4OaLveClEn+QHyVkIUp8QbYyOJT+YG8jwUUPnBE9z7oosQ8WveUh
p+EMMfVS6/JmYUF/Vv6AzyM27fp/ilE/ZgCV1g8UlGJ6qbDJQjl+OxBQpEj48YoCXnWN+WpDYgVS
vkLI7nh2E27gQltjluKDvVr4ohkNzVtdjAbuC99J1sJmfUjezho1NpcNW2dkTLiUfOtg9bXuCMBX
KLYXTAcJzUJRJJIfFuVfSzIhS/f8evsPtzDQjJb/q5VH3rEx27tq1hcCppEYVCe0LDe6LuFTM53/
Ykwvj9kAByNHX2bRo15AMOnKPE7lBdFGpmGGXw/6gW0GtGwMfvBKYvMGWRLzWQN9qO5q5sDSPE7U
Ena7YB138b107da3ILd/U138dECe1QZ8XWy5iSqN2HvIGZtpKkmgSLYFkT/zn18ar6GvDfRB75yl
bkw96ZaeAg9Aw6E4XMYFoHXyxbuWsmgrlO3uqlLRaI/BcRk8jWg7WyydWjjOHhl3QUBoD7FBoXVz
PuDJc/ovwe99y5soIgERn/XLS6lONT5jwU1RJuo3xEJm8hvZkOSCTyRVzMao1isAjLwAbV5NJSPy
alXaptmlc5M3Ktpxhte+Ivv+ia3WzUzg8BTjFCKobDaLJs0TyXWAGJNEDZ7ZRI3R0F6HktiJEwVw
pjIz2vN5d6++q5H3rnD9LpprkRvF3WbTzAx3JlPtbfJQUziZ07JnJY9lasl3kP21KvcJVBZWA8u6
cS9u8nfwy/s0dvf+7w7m83c7+zoIw+5B8oWAW14dbmmnoOCizXJqfFUT2/dlq0CZkBR2mRdVidP+
b6rabudoZnyg53HerbuGKwtjS1ND6jGruAFHVAYNdP9TwMwOn9dRDDN45fyARY4o9YdF5UEyRIFU
Px5EFod+DYG1zGOsWDyGNoQCZ3bdfdZlhoekWdqm0dWKOWMswLnGcvt57UiEpI+oxjKgiIJY21Gp
4Q47ifd9O0/zvGbTas7GtBr/MvAXwYf5cfzQGaqKoR1nx4WjQhXEmpl0naeX+xOd5tr+jitBkhlw
iMzSftHIIb0TEeeu9F/QxSJ1T29sajDmSbPYXqfFNVXdCvigH0pWm6kBsNk+h5hYhzDmiDLjQWbN
ZA0fLrEUlCqBYZevyAPWTctVGj9iWXNzBXcHowkYIo7S0/2glLUza3FjiH3jIyO4/MOWSUQb8o4y
26kf+vxdry3wj9BVBZT374y7T8CDZd41Jt4mBOHKo3lF1ujjhrspU9ffI9fP9NbOZurCP+jNhkoo
fABLEQdN1fhXvEPHJ5OnaQQbsV/5SmzsVhHHg6FMLwZhNPVoxyJ+2FdBW46ptYgEqQJan9yWTcZU
iqkney+6xE+mrIVCmxWk0ZWiW+POgqUKuqteEGSlkaecgkwpH9icTryuRQl2ShXjTqlPwG3HCh5S
8uUK9uSpxscnPj01KOqfOySasofF5k/ZsoOV3mWn8UpbXbuFlJ54vXEANC5dpvWqcggG7EXQ7D7R
/fdYe4+CJcuFf5x+Ei0LYxtuXSC4wpuNXht31rXuKe5I/QbMy3LR5kUZf2X8EMNgNYDUE9lp8fuD
X2Wdu0hqzhf632Z8gtYLnpNUdiR1uTzzkGRsLZXNfIolE0gj/xruZop5bj3aYcM4dyT44wBrgBoQ
W4ZG0l9ICQ6XZmAoaNyXJ+Km95vbHssaqKjD0atBEJOrIP3bzmb3UOH+h1DyMtxDzl7i6TN7PObr
d0niGtNskBXB8lMQ3CAqnd+RRNwRo5r4iiiDJgrzlliUG3LwQfgmds28iOyY+Ogt7pFk63/VzwKf
aiPAyqZPlBxyvMPLawSEJ9SyEjnyL5DgSW1cDUl0QjM1odcOOTeP1ZrKxrBI9/l3DNWKsOn1Pcd/
470praiTOu7F0C36qS+miXyxMxinZAJCT5GtN8YVwsqht+n1d0OMlJggjoaHsiVTZ323DKfaAJo5
FaGZfwOy4WlMxHyDoE92JdXTy3Ch71+NubZU5+J9YbdRLxev6eDxmwmblk9DCBkI6cRlNeHde5L1
jwKQU9C00KJO0lxZ9Vs/EgxpN4C0ylRREOTnLmb/qJ4sxN4XHEmoEhWXxjaF068qxXrPPvs1FU5V
ulIrq6oyXpZRm/pUyE0aUWWovrh4yWYUqJezpuNiqk2xdBh3KaGdSN3NiVCIgBVGl3UlL2o+Dhe/
4NzeWDu6JJbPxaDHl98TAoK+Dl2qKIR5X3KpsjHteDsCmnhHYNl8amTub6Cn5ZDju8aQpGsoFpLc
hg6Ifw+OC2FCENyNCvOPTMV1CartvKaLHFRCrwFhlBvB6beOZ8aV3SJOH3EJJhylQWkyRFaJyRnd
/D8ZMHPCKWDXqr2k77/TN+tG5Rm5wSIu/tfYCRMXaYHTNSAe9kCERYJ5vEoxdRGidxkUWYBJHp2q
v+czi7NjFkqWczkoVoSBWqQmDQDgY7lK6+DM0iZTw7x77PUXC3ySOnfOccVKxiT1+3ond1KJ7pYZ
6N/E8sYT3CzqC13c5foxyPNIJfexlt4oeUQZHo3tIoomOZMJW4mgZd7muodP1BK+WMhvvIMMqClZ
ESNC9Xib8QebL9EBcziItEmuKmDaYgoCJvFGOAXE843v9ALMZV0w3KtJCHiiwGIqmR4NiILAY2sQ
aMDGH5mKynlSg5jjv7Bl4WMwAdqIR9UIpXGwxPw9SFicMRMSa+h9MwgXwdpn3bPuwrHOdkSDGh5v
XMJMDJCHq9r7bP41gOCqIAa9SPvIV+tMqkrOnTxJz2P4YMS94Ts5MKxfABiLnEkz+iE2Xf0tuM/3
FvlFPfyfvhMqzlCVhH5BRkOUDSAxUmyUYhGDkL5OlgcwmnTNe87LSwxpAshAzVYG3mEv11IZv7U3
V030VaLi2LlAjGDrVfla+8hWBvZUo9FkfyTyjRMPfbuuT5wW0YD6/n/Jk5eczVetQ+UIchumu1+h
A/DOZz9Vs0/L7hX2ywYMpeipFxqJYkaHMROdlfu/B/tmYRCJ6KgAoLlAt77wF+4VFUCezRRagN+6
FWFr+AhJrN2JcgwZrI6UpsY1bpoV8CiIpdzmuSVDImMOO8QwMsn59FWGod7S+gJKbDHl9qcz8ztU
9OYSEq6B13WBolHDZ7V3kd8qDECwFjv4z4MU+8+r8jsok+LPgY7IT2LjyCYRCnLO4OQ/16MlVSsL
tqmPr3Fl7dStWqC7KWKDEZx6d5LknJU+tIOI0M3SWh1whpCTm3QUmLnWFQnQc9Miq86uE9uf1st+
3afZfTQBrwJ8dJkSZi6caYn2yQ+GdpF4+T2Kc7m2PNlvRDCXTtl5bPvfClfC5G7Zh83J6PDEU2hN
HZ8P7sEmCjLGkKGcEq0t89nj9ANfUprMNd+1qzOKiebHQzRCPmBL+mGMLvh7JkXGBm+l4yYQHoGF
+e04TiPzt05bIltBoKFKSbDv3clmT7EqoELib1FLNHgzlV3bTXAEXr8r2EMBsWWNrSmhvn7Xp+lN
ewRe3HIvgJbGuZhl/TOsEQFrUiJ0j8/8ESyQ73mhNyCSgrUNQTq4dQnZMvwmVig0cd6XtZpn8dMd
AV69Qb1w8qU4gPhK4iG76oSAhbcv2adcK9Kf+cTfaXhHIQ5usDVwc8NT7PLb5AP98cY8GSWy/pgO
zWGo8IHzqG6xiB1dqlkeBQ07RcF5Y5dfZtvxb59e+A2OiuesC6Aij0uNHB/WeW2/AkpYH3eUQQkg
phstjNs7x/bKBts7O1t6sauKg4bn0BtaoqKxJ8AusAMn+/j0gFu7m+chR5Ly5OL2R2Q+vlJrlXdB
2nDUN+jkUDmgD49f1z0R3N+F98KVWwkdcP+sYLmN8X8IWCjY7XAYfDKEXkjlYhnNLIRMEaFzfaRg
zsGAiTA7jSj2rrPU4UPoR0DiQsAAf1ZCEtkUVZ1FERY9h+PqxvWdw3VB8FkHOduZGYRZ4p8YzjEd
lw0GUqHNHQg5SQsD03KC5y8YmKfq/i+x0CtndzcLgMcBet9Y0yH0E5m21gqs6f2Dc3g6GzhGEoiJ
kQqg7nLHcg3EfKEEjvOPFem1kmnX8tfV1hI9Z6UH3Teu3pKphQdCgDVkkobkpy4VANebFBE1cquH
m66eroKZQlUt1nejHUSIsFLstZeHsk0wWzZJE0+u+Bm8dvKhbTYn/nuNQ+VY/T8+4EGXyiReL0tu
6s0/cMppGPwMnzzSLFSL/BzfvIujWpnJey/j0x9zI2RHRW2AbfJeGxCrkDUs9zv1NrJXhb2MBKGU
9fRGCNoZrC+bOHf47uy6Wv9sQd8B5jR0bUSsKkghnNUE7meceI5c2YqFCzo59vNXcUL4VER7bBiF
HrIQaOP7BiW7rYYIXpCsErbQY4Vp70m+K/vSnjwewTmQiexY+MLm1Q3JbP3oUX7RkIF+8VKtgJ35
jM5XNTDm/J7O+36vmGsrgEdZ4w6z79r+/flfJDeunm6UMPQVJMwEW9c+2uVwPnYbFP2u3R8wOuvH
MwjbKId2Ayob/ys+q0dtP23g5Xq6fSwA02sIkTBfFCGIz2+ovv04Eo+nU4QENpmq78SqFsTtfIOl
9qClX86XdDyefED0uM1qid4pYyrLBcqOpQJ7lnP4hOo2nw0jqyWGpFjuzZof3bR1sz03ZORjUlqs
SHq7OUtbR+8cjiGa2OrO/CxtzGH9/hHV4gjKsy7FgCLPmeyIg0u5hUBcpkjRJI6lxVIbzGdsFk72
XxYTMAp9XwToZ3oMzUL9/iQgZ8mqbVaV5PHjucvE61o7NyFPxZieVmPA4WaG1QP/DrSoQNOSCbQt
6mZlr+KOA3xLeSL+IFdFBcIFNFx4VaOw/zG1I4AfhjmsZGktlo6NZClD3N9695PYto+xzDae5fub
PqKrPS5OFrI/2dCa1AcIZJ8EaVreYhPycz98T7CcDzK4MCmIAW9qMQMhvSFK00zqD+TzIvsY5aCb
Zdn34VKel2Dj1yi9RyMVYcQWHyJ8ZQVgYA9LvpYGuprCGEmF9KjM8XyxpAKLCFXMVVxspyw1dLsT
MlUxkMP5cvoeJgOxHIOZt0wpAelltLKEhspKvC+p8cnbVn869PaeFw/A8nV8OA8VIsNcum+p/pS3
SMjGoHwO9ItcWLvghdfATfIBTpyicT5G8Qx46Np2aCxfxCHUE12ulEWo2kAw8xBE+l2EkjHxpYu+
M1V+lM/6a8MP3uv4BUiwZUD/LnPo5jZlAJEqlfPwdOmAHmwnl4ePbZAE6R0UC5SuHtJRBybMEDeg
ijDlNVkjdELxinEsBzLyY2C2lPdYbEJ9wEsksBWKBc10cSWkBCMNShO6OAaWoSyKUhw/ta9p0FJF
BzGu2Lrxlq4rnCtjWoJcmqO4mB5sXRE06wwuMHUvuxHGIu/t7gna1akjUPdRuvK/I8Ob8bf/hyAI
86CsBwZ61WDHzrFNGb90lef+P4biSrKStalc5ofLBPLQqp1SZQJoCWAa2DiCZASgAPwWKS8I/hZc
uv5tsC+fqThRARHZ+Om/QtNi0hMqSzKTpc22o+MIePS/pcP61zl8NIGLH2GOGLP8k6YXSj4xQYxw
pT7r2c416omWf1Sqb3ep5QQby5dSfgDJUqsJZDM3dYNCHFVjwJm8KBSK7hKsNmqOs3rNj79eQESF
61iTOb0RYZ3NlcfyD5uH/vevYg9FEhqnR5H7tvphzZh6cvITyqY1v7VU4aoeZvgkrFxMXVCD+T3K
btXQz89wd1y8Cs33hPGNSxif6djXz13G3vto6lppzZS+5Oaju31IolAAcR6KconnF9ilgUGiUoKH
337iyFS32d1JgK/OBf+LrsA5OPJSoCJkC8KiWSWhZPKYHJOeTHdgMweJsarqsVqvBddAheR8udLm
Htnyiw/2cEvTyKNFNGlj2hlW6/FU5syka2o7/NvJjJ1g/ZZkPdOzagRZNmLnxco/+zo8mI7CGpQr
A8g80poyX/T60FmAaEo0xEkKI1SYtWoscXFA1309EACG/DZA0anOpS1LWZJVmnLlSWVK0jqFJq9H
Cbe1At60hySFe+rdk3XXgFZxfj8vrn/gVGViF/dW1p9wxYoxuF8u0qiUF67sr0Wsxi22EflY9f4o
PTRGHtnWW4/31q012oI2+rq9Mqu3vDsBnihJ1VllIvXKGQjv0MbnDvUkCwG01lJ9X7amlrW7fze1
SwB/TZbixZfPNdAYQbly3J/WZeBFUPemeUknbRvhbJ80TWF2TXxPId8UzyEjjQGMzbprs+INu4Ar
vAFc510jOUqQvYnBCbg13N/MipUtv+s/BbTwCeIEWeawTjRR9RURaOXZt+HsKiZ+/s4YAfRoU3zz
2fd6GhO86sbi2ShxarfwVonm2QpRnSHgdGgarVhwvQlUb2Y6oyql0O3QYv/X3BVo4mW0PUgQU1ee
KYJUhwz1mSBx0ZFzvpAMztEzbm6gedH3IVPRan/v9GsCpxmNwszR+hhVSWRbTjUPFbOHJ0N+WdUs
e05wksFgzM509MTwRPoUYeyjlQqDbGKp5rT6WTSLiB9wAjFyVS8HO/JOTUfCRJcVcl/o0L8wEHcU
Z2tPs3ihi5HsbLm8zsQMVJCTkSTlVj39XHotD6qCIwqdyrKcwq8BTvBS07Ta796tBPj55by9pGvh
AWQh8jNfHIf84oKU9MlcddRIOg5I8+t+pb9NL0owG8+gkS8m6Whgm4pAZEBxI65VYUr64e+SPcgk
MNzfD/oksQl2irP2zJSpAudUpEBZHKznaWPW3pb8f1BmWwriEnIBY43Rj9pX3lZhxOWnmjsY+l43
9ETbcXseWzEw1i07gI4IN+uWTO0Y9nYNeJeWvNAqcpx5spTiaa+TYKj76KupUwpx+U0HrFjDcdFj
Qsww5lm7wT3L9vUz7JERM/fvh0utE5FhVaK/quXfggEnkHbVrVW0fIjNuGn1IKUaP9/6c9zoGC7M
893IaCo25qk4dc5Xyoth0i1o+1CbO4mQ+HdwMMj0UZxSr3y4ksnqLq2UzcMSBwmet1ZjiWSkK0AE
PZW2pCMQZu9eZI6YnnD4N6vvg6GcTWlDDVRy5y0Q6fLD91/ULDL7ZKBEvSWj6zaqR+wfruSNZr9b
LE4wvTMyxiv/fM1j4sEGKY8Wu2HvN25adgnlggiMA32G71ZlHLJdMsGLnf05a3FK0//GT8Mbr8ra
NSkwle2Rcb+5KbjmMJ5E5mKjzGzpZl9/tpVr61VZERN8XHRBJ1OmAsFUu5dm78DsYqH870F3pFxx
ZZMMFaCyxKyLixFHxRFsduuuGb66/khO6OJ7CvEdEbANrkcjoqKjC5BKeEEuhFjnrp/wQo9ncY7q
8kRs8+pXD3PkZkfDF3S153FmmeWtEuzE2JB1iB4cWJ3F0/+fs/4MP0CN4MpiDq7YCSwk+grEjtcN
7GajdAVfZglTQin0LhYRrv0/8RB7f3DMB1qF2XRq8CY1JJLcOcg2JRr2K9ErWHqoYGRtBAXhYiyS
6SYsIVFWZs6h3hMFPPr1O8pfF6CgslENfWWIlUF2uOuqJ3tJTowJmOZNoMyRupAqUReDeGnGZTEa
Vz2Ng7bIF7GRWtcVfYHZ+4wfyvlTbyML4nUkkPk2G4ohsA+kSRPOPtPU81SPi0jYAfspO2wKsiQy
WAuAfuaxDTTlEiBam7MF5zoOfZxbRGi4xINEhJpaDl/e7nILQqp0wxVdEF77G6pjpU9Zue2mMSse
6OEA4+Hd8NvGRAi7IJhQc7ybh6nlZDjd01NgWN1QIH4bDgsyFa6wGVL4RbG58cYQ7Ah+7K7+rqJY
uPy61HbkK0HNxrVVW8BGYMfUxtI0EMHaixtow+Tmg5NRYx0nBocRUeYj479zTXI1x/Yu+2QPGfPR
QBtrobMMMduEVAego+o1+WrJKFWRfsZtpdve684F81S8T3CTk6eBNt+AiFdKCYqHcxandkkPKCpE
TuXofVAvBkFFziB7ox0cGdoi1uML/VtW2LQ1wggW7iekXuY04f4gPy/YqzXUVgOTgjiuW/W3bM/I
Z6hp3sFFZi3KRyB58HoIOLFdZ96+MxkncVcoD8pzjI1GokzG/hUCHKRdNqetLNlyNjdLScstmm2n
BXf+CslVFCxzB+Aj9XnbV8sHcPlGZ8sRcTlPUiA3SorR6anfazCA6i1ZyQ61Eqh0+SFLeVLgoMkZ
eMtu0GUiOp/PgoCSfcoS4zvTBxKuWiy5LDK1N4XOc3e5byfyvdu6of3HowZ/4dhvV2/7Ce901twV
bQNz6lRGofzlNj5lfKF1RnbErz3NawYf8cWDGetCDnoZQqEWnjk7DWGyqHcEefLTgZrav7cP0o4t
vWZgb6DnPrY3b5fi2UlOW0iU0jzWqpLuQ0Gtn011QetMMUAxUIYkC7DNi9RpckhkufSV8ddlp0H/
Ssb40/c0pdlRzriCE19oxjo9vrx2gYYIKY5bnslfBnbsdlf5Hz6rS2z1GIeP1W07vHPhYk4yE5sq
ug354D4hohQiuvRBpTo05p3F8vqwP47wXcLddWellmIifs0uiH6tULz7oRkSCa1loCJQ0Z+csQe7
1lKH6b3Ts+aSXHys3hCnDiVh6tEhfFpUMxtL5bY0CLsJsYhR+e14EGiexJJEu7lTQHiVzgZxTH7K
2Fb1sCWiNtqWAlxauI5Me8IQKwRBx58XJ+ZC4JcRa1zkZAHJAQyrxZ1oF8KtQpbLMYyr/l5Osy83
/6rJzEp5q1jiJxzojVxG0PpBbot9Wjxx0/2viJeN9GFetk+3nsnLDsWOiEFfWrI/oH7YCmZyUmD4
JUFvXQl602LCiUOz0V6zpf3LCikNC/Y7RNO8FzykawARqpHbRgiF6F4zG6Zju180sMzJpbJv0cVS
/SvloHVIFajpJtNON1g7tQzfudR4O6680vpxGfN2mfbiZf/GzNYc5EGBT3EBgrT7eVg55nWfyFRz
I2MXAIpu6dURwOG2w1i6HNDChxM6aWPP5MipEF4RRL8fp5Q1XGxINL+/VBkYdQbPTpy9NVKQNjHo
L1awMKsGJ1XY+RRTKUMpB9vfP4DxwuBZuhtKvDkqlVmie0JDZ57ssoU58LBsmKEQGvbtPeLo3eKY
UwY38sgZXl5k69NxNUnwMSH+FA/Byd0DAL8BEEUeGapktQO91lrfAWxXllwEd+1p9Wm7zc11nzo5
bWwlsGOwjiO8+t1zE/EjduVovTJ8CNMGhNFzzBOG6aaNx6OU9F2PJiOkXwnuXmEiEJ5PcmI2+lfc
XYkg6cGqO9YHKP3NkbSpIGpvOYeyhbVqfOhSDKvKMfzRhJbsk0k31CpOOqbR9LO2cvnzaE4c3vsh
LTZR4FtZ6dDmzhs/ZVAvTNxW5xfwMVjLgU9jCWQbxg0Wca9L4uznuYHJRWk3Alj7xukLDcarJ0oJ
a4uBe+J+0ljwaDcSFKdnSD1r695GCn8D+VBWbD1JqduRlYEm/57+Z/I4XQs001JCU/l2NiNTkFI+
kmfRygyPcM0L5qsRMMWzTzaNg0J9peaufb31YIAG0Wz6Krcy7jpbZ0b8NiQvHrTgqt+YoOaLb1gu
tJyfUx4Ksg5wWBYaTFdNUHQGf/6qjwtDSeSNYSZYPwnkHcnmGUXJEz0LcQchOy6syWk9GZVN1MCM
Tc/mHJA/wRxWCOmL0CTZW6sTysgCBJcE3NITbwyQCBLL5VeMvqVHTMJO6PJkfImWmpzMQED8aUyD
HmfjvdJbKGDl0qDhbTzWyFmrNOCjqruptgHEhufcBzsByrXmlV2DuRKYdq+Xpi38G93CdkCsCfi1
ShYXPKQfiQkz5u3jXs9rQqdmhq/LQcxQ+CeI9bKWKTsDMtKVMq4mcsdWwJRuYVkDEETo855qF1zc
bfxX5T3cC47Qfo9GjArgME0cDb56EaIlc99IrnK0GasbAVlwQXpPX9uCDgs0a1MPfozF09o+Dsbd
JL4b/BlZlEKb0S4I5K1bRltRHsaYOPmh4cxOC1j4knEmXoJ6KYv6hulIRobvCKkk+WMODrwVrkGE
rNaxMHwW4PlyNWBJRecvU7Le+3q3L1QX/lHZlP1CqZ4qLOxEbDzBxMBa6ZgFw5iLEMDXQpuz7hTc
4os7JrdV2NiGrF1TNuBqsDkeoMHeZJFn8caiXEkrh6CSIzEEbiZ4/QL8a1pgUTJc+QipkwZRTc3x
Zykws9WYslyuRglP9nGrUvjcq8Xazp3Afr69hAcRduhN6CzGyNEz49yoyZYkzsL0++c4lPkl7BWd
OMAncgvz0AZuHlJ2xIJdcpLkuRCCrzo/cVbxD6JONqM7hSti0v2Fk3nqNAWaNrKe/Vt5ZzMvrxtC
navwEMhM441kkLu3cjdz736gm5IHpDLoHwKKtVysv/TKrhB+LlslJjIiXFqp49VLfFRQXAURXgXe
FFAUZ3IP9oxoR29uckUh11XYcPft1OBtRqjOSDIJMPNhuQknNOmEaQEfFnxe2W5KhFgNoC0CFfTz
bYz4b9ENyYFqiKiiSiTYlswCR3n+Y45umn17+NUX6wN7wEpsm8hMpHCYc4CV5SBSQueXycOSa921
h1XGbjWpZmcDMx0n8OzPhJthvkciDE7umWI0MJOl+S7hS7fbzAuVIawvfHpG2mG+br7RGciwxkPj
u+6EA3ZkZYhj+IwPYAVDMJZpJMmsUz/2KbFzgGjxMRhCC7jdTmeqVogUX4sEUFly1mDSuNm14wKr
/X0erSyod3mPVyaP9UuZC6pRL8Lkob4IfOnDKGGPLEsC26iNfzmi/i3h5+v4Dw8suJF0xIzIu7XY
iSX9+nF9TEiyf21XD0MMdcU/lgW9UOsIwd0vmOIdhxiFZz+1bmV8pYCZTZ/mAePhoKxjjiVA8I+0
4Xy+ub84WDe18bny1etaksJnBmrcFvw5jDvsomSwk0co++jvS7oOt3MWzlXaB7UTEowPMCohczbo
NIu2NeraMjIixNYQxQG8AphpW/k76jxye8On+WwDFGFPBql4/N5sI2OZN0wsPc3EUTQrow0l9IY0
ZhwqC+uOYmsd+UCOeWUeJ0DKuB/M1ntyJcMXoOtH3ykp3K6UHpnTIuKAioF/UQTyn49ECFmKdJU5
Lq/uSLs7qSxDAKuJyl7aEIIIC5O2Qc6kywv0W4bJQPtWE99D/98f9Vi0OQ5SQBa4pW5p07IAHNmf
3tKvinsLwYJmLpXKhs1aUo2agOUg9y0Sq45K6VitLVfa4zy5Ii27DlaY172sI88yPYlW0QaaJ+8S
W0b/IBxRwFMQsLoGzurcHR2sDNT1YQp8E+MabQKt5bpoI7yueG0vhZcn9jOfjs8OkdRKm4twRHqA
3NvYDWU4EkQJmT7OrUZD5y84/Oun6+9e5Q9gV+AIoLokDSJxFL3lPfEBb4Kd6ugsD2X1Pgu7dBXT
tim3iaSMl4Q9iUzoccjxMypIRJ62f9H0PsAJbMS/w1qa/CXQwddUxWNdw2IieEhL4xTgdSDJAMAi
63bPTtMV2P7NchEh3wzFanazKy/Pf0Ecia39kpGy4CjeZr8Y1+knSPcvW6Xpmq3dWpymnvAC1Tj7
K1NGLHXcfNwabP5SbDSnm58kaqRPRytXFV73YtgpWSbMaCjA4SdQ0k8R+Ja8oM0E5QyBHvDuWaR4
LzrJbnu1R8JYlUxz6SG4g0vt6rt3V2xGivmU7EPMESzxmkJe/NNyWKAukutT5nS+tsUOJMw2GuEO
OxfDXRIgh33uv4Q3b5QvughaoY19I80Ftt6wyiVWi1pjH1kSbzDVElbWiNn/8LfAq7lEOm0V16uk
Y95WujW2pv7ibu8/2JsLMrbIXV7ZMSQCpv2EKTQnuCWZdv1LTMTFXOo/1K1v1NG5zqbJlz6VIe6B
Bcz208BcRBOA5f703DbhSGhyh+htl7vVa9HZvbfcTJZlojfSovCPNyRGRT6HKngXNnpVLssHsrxm
6dkf7EVVnBn1vI7JnW3iUZgKQXJkPfe7gjEEFlfeqPjldtBgtl08qU/2atSkV39OpnAYZkXj2Klt
CeYAv7Jf70PinxHw3twTDHz28xmZ8N3RwJ6KXsPlSnJWdi1cTKW+VWK0+bCG8Y4cDNZ86JDccRG/
zibwAeZJbSJO8y5IHOrihcl1df3WTx2LD2brcPuT+Iha+FltTIR3K94fLBjc2PfpHtsGhnBy2P0r
6+k8KhfeKBL7pOx7E8mAeRikAhAuGiRdf94H8bZaXL9aCx2YpqUmHXTiCzul3tViXem+14lKBaDJ
K5aFTHC1EmHvqliPYpR9OJOLtNo/YT0UrwycHXwnIrhhalS/QYdT96zfLpsOM1IhKv2Z2VYIKIy4
Sjhxjk+VBDy1pqzM8qBz6Hp9VDK++4mIxbswnc+n9ZViXHrwLI5rg1YHzvIMJE5O7duoVGNHx8Zc
uKMMfNwqLsnCtyWG+Btx+OtQwTxnG2LpoU2jvYnFmdedVIr4jU666DxnyFyreDz1IbgpVD2F5E4R
TykvVj+jr980DiQArGjplhTtYSNtjl76QtLd1RKnjtdxFFYQZpXZRl1oUaFJObYBYBMwizs3QBJy
l9Miwx0jMa0LCPhkkKmVCsJRDBQX4InC4zEaqJEhrXZgokLPVk8YAV2Nz45xxlv2AopCrE/FlkK6
hYNgKdlkNIxTrsyRzUi5Vzvy7tSsr3wJpsI7vUmplRy2KNg7kYkXo23DpHMozVkdHx/o4wcp7Ke0
Ji559H9KQpLlksqEhDaljltbk+aB5YMGVfpXxEanE2wrrIBjwf3NXHl79CxJKmaWzzBZsMZT6wcG
4CoAV0ScQke21zYP4B/NWSgTg9cxHm/2A0jRfbscJazAobTxKjwE9ehGr49jCBohYLCz60znrVsq
72iFLsqXatTyvh2ei4hMBY9lv/2v1hdUXi8a5IQzapoP2DHzdpJQL/Ls9RgBNmNBD4J7KzaU4jsj
W+E7ZDX3yXY3swEL+Lk6ODa4+hGgqDRxhNoLmT3y2tKjPuNUosNWpHBKq4D8li9uP3+PoX9c+fFp
we/nOLIhaFDBwt5WCZrWp+UB4/eOzKFiGtm0m9a/31hazQ6/ZgQmfd15dD/PLCehpCt00JRvG8Ko
HLyI6bIkcS2d0kkNxyBGr4UTxhJT8V6WIP5aQS99PzUPy8whui6M794EDEQyiKwevo3kFGhQnqLk
TOuemLOc1wamMjCuO4ePHjiPFyxeYeCQ4lhfNiG6y+d281Enbk8st5vccjYNJdXFRlC2WTn59DUU
Zw55zARK7MFW2ijh/NBIdwAReEX/Dc+3+8ibvHnfzcoEntl0XBGpxmZmQn1l7p3UYnyMtboVy/s7
mTh+EYjdiWj9amRYdExfLdnZCb6HesOPHzHaRk80RoxqRcFU4GMN5oEA5oUWn0lKnU8IO58eGlWl
flI/souFAMmHHBVI0w5Tvd4sCQmgry9sNRgfyXOCzeIINsEa3OKVBBPll62jwZ89cSU/HmME6N/E
saKpwhjOYciH84qpP0mHQTgMJVIrNFkI8vngfAMKRKR3Itgb484EYqxikcIcCNOeqvc6f1dGqv0l
ZCOsfH0QAVGA3C0OJNrTmaoWvjJ94yZBUVzO3arsH/oDx5bKJdUYUjzxcwBvUT5nax4xH+/u+wBj
HmyqL1dlyxT+MbvhDEcmn5lSUqWguAYfFghJYFRurqTH0G69XN4ukfz/oZ73BrKVfccbrDktJNVC
PKRORGsnzNueaHsJt8P+XRp3DxmYEzTSHe6OKz6v0DbnfOWPqp/widkgVRGjBT6PdsXXxDqMtg+n
J6YFot843krTmrQqNzUh6fe0nzRSnbLEzDZOnyhugpui+6bwGSf0zMlQwrafbuYt9JK2R7zRaRrp
8jEyQKCoZehrM0Nx5nGtZrtNV6NVgz4mqntDcdR/JUxHlCn2d4PdHmUBm8KLPp3wnZsJVJalDB2A
Wfl+w3SqSa2zHBiO1WkDNtbCx+AbHW6a93MEZq7Nr28zWdmULP+F7kaMTqnCrsOQ32vil8n8M/Bn
J904wkpE5dm0UzB04d6lLw6BqBgUjHezkMCiY3x7F7DqpsZM0fpdZ6Q3KVJXTYJiPR01Y7qr6MPn
Br7nKQ7yFCodW+t3vv3ry+HjJD2icor4pg2JIeVOkmF/M2XwY8xAkN2ahGKmIQnGzvBbhhuWt+9H
trw8e6ltjMB9evP1At4vQmFFJ686T78zc02x2Ud1Qf3U4NPfkOQC0fV8HzwEk2hE0/5D2CeVfwZ3
bt/qrO+MYbuamDpRbAOBHrJEM8KGd2qC1tapL0P/mqdp92U3vCRgacn4P1llAwn3YIHrOUv5QzT2
1tmt2VsIcjaSqSxGX0SO/GFenrxItQNq9gojklmRzOuUoD16ZD1Se5GFLSvRoWcoap/jOMDcoLD7
fmqPPV+Y5iHD56KNreZCYbDHcoD4d5CFwApXlFgcyDfAdhmIT5pPCT3mEBVQwtfKgu1dkKzZmwua
sbFvyYhFJimd/tDiBthhc+oE2KmoTvt0YTxoQm8D4P0bzRXCJ9lVrM+4doJxBhw62A9qqBJ1axEe
YX/SINJqaEp0m1F9HDi2Uuat1BxsNkxLiiDgktw+xRxJKwmw3WWSM8vlgT8HoDoh3PJCvOehA/xU
Zvm3w81T93ejTR859g2OYh7lWojYh2daQgSPGJcHxuSJ+6IE2jEzb/hLtRaJJJP6wKVn9SAyc1YR
7+StpH72fiP5kCwq2mJ4R7UFayHzsr3G1H7U/dBeOeDo3DHZvccHhKlLkhJp2fYJI/dHAajnRYYC
nTbIMKN5rdwXvMM06d56O9IR1D1ASHK37fw5v5IUXGbSUkojr2gjeQPLQ9CWVx+cbr9VzpIBl7NO
8DU8dLnyfU/7medFf0xPGLFMeMNkHspHKrQmomg4xlZVqOAortnO71rQLdTbqOUJjIvxxKqRfl6O
W2LOJIhCSEC3r6NTHc0osBtetOOA1iDfDmagBNakPOGLeFjSij2HTCRtz8QgFYLkbwNop/O3s29S
E6NAVCiEMpbETIW00Wy+pGw+R+jYFWoWU45xWy306F+lkKM9zDQzTveSh42l36/lm4nHIZBLuTDJ
4z1kpOgIgpsaE5WKdYhHWL9mZxOwVRMWza+PLJbOSDGncSgJ35uplFVs2H/z4Oydu38Ep2W7j7eG
u7NJDVNh0MP1GDm0E6qZlNuUZ15vWhTqtO09Du/8jwxQWhpofz9rTHSXcbSaLwqq82tAQpU1a94t
snhsICSvlUN8eFrP7KBv1Qch2UaHgZpOo47yNFYCmmMgvg27eGBW2nFYHpFOvKUuZ0rE5DZBt8tl
+w1HNin8yrX928KOrpaAQbZk19BS9v1LpCPrlwWgCZ/tSDPO64+MFNBeYaAsJop6LZJ+0bU636ob
4eFPPgvF4XZnRUtvOeZmuJxfy/BY6E0ffm3KB77Bpyd5qEZwDFDUiFHMSs+UVlV+ga7kLDxOsT1E
Jhmug5JJrdPgXlpa1r4RYxO+QbFwIULOKQigkMjdRJ+bxwiteXQ7B/z32GiB/HGeDBcFD6ziGYHU
wKRjodQKKhuey5T13F0LHcs3FIl4s4pToJZ1sLAixYwPbrCP8odvAr5oMKBFl4raHVzWUuH6/9Lm
AMXaQWiJrwHdPv3SZsGNBOCeMOgrcDEItwgzL7tyRrX9vpG3DXY6I5jk2Fk9MLIgQycuzVJE+Sy9
3EKj0Fnu6kWGRZBEHLOPoxgHzNXvH79mwifVgwhQjGzcLb9P2BhIR5d2I8L6m8rNwory4lanwRgH
j2HSN4U0vXV2hMh+XjzzcECrwp4abkm0oBYSWM6yn0EEBZpEyDL+Itio2cO6TAWfunmF/9z172Rc
r5g64MszYV+YuDcU2BWd4Zk7frEUHu4QlT9iMyPwb1aYhKtbQNY5mlOfVwV1rP0xMFMS2gjjK7JO
cNzaUbh7RUO1Ge43S3dtGRz7iT4P9i2tFFEzvA0QyQiq0NIsskPziR1s2ML8UBj1jPBOhxAKeOrG
E/GuXXbuL1PvXjdPJKUNUulfg/YNyzdmDchAix8t9UFxz2ZK7+gcNve8YJllc6PBEM9B0pkzQ9ZX
PneeZwJT4yGjRE34xro8rBrSrK2GrFaGkxXocNrfE0txO/rS43RTOPiBMSdqQ147qSNgHSyCeRDp
oyNIubtVHikpIJ4eXt1EJCo0lk99tASKUcFSeWC92apfGEutMvQpcRwZMqd+l1AtotNtpZQSIPlB
jcXzBtd5R8hgc2HLyRKF/M1CznFLASKFlHRalwfuiMdFCb0F/0BZwuaTe9cMJadU0AHLm9DW9k1Y
r/Q3dvZZxQJH6cHGH22L2drtEJkaL1k0sZMuUMt1EgnpTjAbqXslUatjgPqXIjRD31FLGl+7vzbA
ZZdpa+RMVOtVnkgrSbJ19F4OlO7wS+6rGxYsi/L2BBexOwwv2TMZ/kome0uX62YU9m+3vDuW6gjq
ooMGv1jWMvks9MVcSpdzjp3ibs2YjsfwvX76fFFPcvBQQ5WyrArV98o2XA3+MT9HBOb8eQ2m46fe
Js2ZP0XimNnaCWaa5habRzNz2XRjqcp4ta5LksRFgO3oOPsUrTHH2Mi9yn6waVs5Bg7cF4CxxhGD
JTM06hohSHWrL7QfKcHhzn6VaEqGXarziwk20sreQpHshUhh10U+/Pwpy5jwzRYNBQbwqCutG5IO
ldqW3He3jzgrmYGE+IX8z3sWQ3vtXM9izDZl2QA/RXYtN3DCaRSP9cFCW/lHHnVt5JcGC039tE7x
KUNPwg1xWvObDTN5XMUZwkzDwsK22X0mlsUkW9pme2Q76k+UH1HW/Yk06bwKiCdEesyLlOj7ekE6
/3bzjE4lF1lIVQk87Ilp32Tt4fRJbul++3mADSjh4exdv2F0stqyEpQe9NCB+aQbZaRRlMga37K0
z+LtSeGaXYNTQ2xTzfXeA6GrkgnkBpfCoFVdPGkZlALmdOA5qSJGBPvWiFQk1bruuUV25GGSgtbW
TZnck5roSDd8KsGn3XTyCTSCh0JGp+FYOv6bCpFV6Q8mFBQ84nPcGiKSovy29FDq9h1fpz52wI6O
6rHgHdOJcqXamVhclnzznDL9Y90GWBOmJj4Se6+bWQtCuzWoSADgO6fURIym5GkDD30d0FpiSnP+
S5iROzwVVbyiSQv2hUPXn+n2vN9q/BrxDb6FpPqEAC7DXVnyryUcvV3fRXfDR/YMpxjQf0eJbYxb
1bITkmpzLSUQ+Yqz3nLZgQCUFSgkC726U++GqXRgCc2dJ36T4lXB1iSfNRTFBoARnvgt15i+4RvX
sf3pB5ksXsbT7vSFvHS47xoPHnJp1QkCpOVKI/xgqN4nC7lhiV9KGpfj1xla/iZIvanhDg7uQzSe
B7hw07bRJh58Nm8+Hb8pgTOxw+9VBZJcmQs+PtrHPJpi73Kw2mmSyTG2FdEKw3OGGg44m0+KgxNl
bgJY3PKcuscmND8A8M1BYLCbTC5Qz1es3g36to8PUzujb1FkFv7FSwzmlrWfsuLb2NpOQNZmLO2q
xBZUuq+4VEXZbBPzhnXAj5l9ycNttBU9UImEw0P4r6OCNgK/7NgaYMP2hT/Oo6y3rz1oZhyQBj8l
Sa1ljw9GEYXl1l/JMwa0bLJHQSnglDjHN2Bo1FfKTpeL6tQD+aiai9xhkaSm/rtCF8x7+7gdzw2D
lB13mfUPzHIB8j5CLiN5LpkCiA7cTkeRwbHx75V6v7rffy/iz3IYGJW/hUJ4zjd1CI3WdI2ht2um
m+Uk49DaPo/wTmyxcXG6iBYrUBsst5FXSFe4xXukpc8sCPci86uSYf5d/9YooVrVxam9EnZtwIgm
EKQKS6TtUSkjoVjgfDAPU/gXT2m4Mii3GofTgC3faQNfyi1kEsGHlCWeYRwi+mm8OTWhdHIMfVS5
m159sU4rzy72PWW0lxTNrDZH4KzViONliOApj3ve6uCSYVTTBhJlFrUtKUVwc5Kq5S66Cv2J+/Gc
O8QVBB7V37vMcyImEOMpL5b3VAX9k8cFy6IZfkoGRAVkpZ2tqG5JO/D2F+9gUeMACNZRoa3Zr6SE
IGqrBzfhOaw1LDrPyeRI6Jk6DaopfSjdkLfMiP4fHDzZEvHHZ0B5Sadk6r/nFK4z5N7sMZ9fJFrR
DA9+XUIKwZLa8od8NoIYhLdKNvrhaAsDjDVN/TOATqcz7ZkJtlb6Ta5IuePkNeCGG7qZK5tlfOto
h4dRAZ3g4zRMtY86K+BGCaDPoRBCrFwOiwp8hO0zuLAAlajoM/wqAoRix3QdbGHpnWMp5OCbEq1/
atjCXdPcJn+iwmI1dRqBKWhwtodklmx03FdIX9xvd0l+36ZD3+tA4tsXN5QzWIVaUGCHt+je+DFo
nMOVHwpiITNPFWaQU+XsZkGd5ZD4GN39U13Z/M0k7YHZjCH1oOjkOaPe59U4feCRqQcFAhhLMVof
+5JMOx/wziQeMJiu961+MKgK2ZifOMRylDPDEAy93oEBj5K8EhI6BhqU/zwisZAgmdZl0fW3xUAX
5igJY+DGDumtU+0KTs8QXdl+Kexxx73/x5Sv79ZtGSmfh3K3yurE4N+1o3Ep4co5XDQsyy4n4Cwe
p4dh9iRwsdpItK93kwcB9SVwZ1f5WyV6IMhDi/WsGR1xRMvHueaOpGnZ36NQbLF4cfBjbxjZEDOS
Zml6lk/5VSH+nazFWkrzLBpNbuA8wd5d6uIj7F34uVfnJGMQOhfVAa6TCXiVfR7jvUSTx4v1F9zY
NJJi2RFDXMfXrpw5/SBLaqXYysccBGao9oW5y6qYLnFR79SmlqObZkFyGeIhGdR5vbmr9lj0rGuS
fLe8yioPy4anu1e7oWJ0WX9S+9SjafSCsLNvmFaStcFyUnNyEp+CEzDtfbOiqbab6GblOUdxTLGp
humSBISQiJ2mLgiife+TSVQfIOLilgbbXmmSGQfGArj5QusmDr8+B1HpgWCXzzpJXts1Xoc7komo
7DBzz6e6EN0l+g/XyBV/BWKkToRolF2IKD9Mhkdk2ZluvCYJZfR1R3JBcgZ09RM6VB778Yey7Kmd
2KFw9C7pNVCV3vJIOqogC4NWrrdl+gzA7Oi7o7VtrQ4k7+n68VIAU51NaiSTpdCMcPNsvqhsjbXD
/RXStt2rs1OTg+xEthOiH0GkTmZep+FkjTXyS/A16Eodnb40+gZq/wJStgbv9kmWDmeLJXJxF78G
10DbqxySRr/ht+Rdct8RlfGm/WDCs5KpbbGkcWHiyS/8SUtiLWbu3i7cPUxIfW6RWnTLufj48U06
ITIlNugcFaVvMz0V2cQPXjKzbR1yeRIFowPVtH7XzpJpciKQsS7Faer/Yd1iemWtEu6TouMP13f+
/7yiIrU0NV2cGT7ydlerdknaj2ezXvhJd9e6iDOpoQmOeE6u3F2vmGMtrzHys65+IoPfgwY0q1/m
nuwvpTyTAB9c2MxhfnBa8sH5ViC/KBgD2AHtvjeNyf8VUCSJ5eVO/89FBszhaj4HeRfCSLRW6pWU
sP0+vF8PJynA+WfukvC4GiZazyKW5x3ydrwAKynNoE3WQS+yrcvcCp4Cs4xBXvGIO5iHNJvo/fVM
MM4JkskkBERdP5uitGzTCl5hxFhJZjZ9fEBzycqSJzx1O5RJSOk0lTln7SrK1GRZInrhArm5/LBM
Yl5i5PPKVMlrQNqHu5nvRsJo+dGqO0XVVwu1wxyy26rVfg4JR6NaAxMd7GBKSF5a8DAavqvEQDnB
4UDY/uk5rBPEWDVccCggl7g8rxP70ug+ZlkZpdMdsC6wUDzQqkOtdgT/XQMUy2ZrEAirhQ6lKh4U
zej2vD7axroxTPA1+9k/bYhD+sBiP/oenuBR+7QXz9+SshEGrmLB0nw5HDZ4YPFX4F6U4K3IPglZ
K7tZ20uGhuyX+VvFvOwQZ2R2dFf8ynDfEQZdPhXsL7WAvWwrapx4XthkMZln8ojD+tYgkan/JEY8
c7Nd4sHFydN+2OzVNENQ3/FjUiBcfb7FgDNwWbgNLHhL8doAbBT7xnkD6zpsTw9Qqsai/jjt2thk
+meOrkCSvZvKpGVi9mNY8C7pW8YdFezEcDuKBulhK/7i4dqL7+SZN+QVfti+sdDODa2v95t5zYii
FR9C6/pXxu3vExCtqUCs/vXLaFF0zz68rKrLcMKgVRJUrsdbJBliAEgRrkCCR3HQm++drFSD5/Nv
OekyWIE1S49iMcj2AvavskGZKR7lviFKt/1F/1XZkc/rmRn+KWsAv+5tngwIGdSPavaxWQpQ5Vas
0MqKdJHJ7aWSatyNsfuGmw3q1qsqqLS9kVr0HqArqAbd9RMdnpnnvGKNWLaM3RSQeO6B5GH/o2nv
GoAPUCJTqa0ulGnazqqPCgQZMPRBe68SUpAf1I9GHmLU6gri4k/9IeoWc7t5/eNHa0Q7knSAMrYO
Qr6nR+Qn9dXPQDkxHQIr4otXq2fvz5oG+cu0ZiEhF8AhVycKOUrSJZMPl8/hRRT4CzuGxes8Wgl5
QA2bWTC2ihi8ULjT0BSb/qNnslXt4g0EautWIAL2Cq+nkUheXSHlccx7aLSelK02ejI141dJzahp
1spLc36NvXIw+bcFn+xAE0N5iE/hCWBXbq/3oSz3W3VrKFJDaptWDpQnams/Z8GcHwXhG5v6X8ld
0maXKoqzKzB9x6i+BqtTNAZAVC7TOUhCL7r6oBaQ0HcuOkxKyq1fKn8vU2POBjZKxgPXB8iX2N9A
VLrZWAEDGEwE8z3NifyBIVqVNp8Alh6svjzqAj5pYqieuYiMk8P7m7+YSDD+uNmyEIfEGUoVzNLL
2+kcz0Wca6sSEAGSXvO9P4Nfn9aHGxFkjD9yZBcnstrl6fy9IFZUY+K6ecU9yBKFA2Iov33lT5ld
sDYyQdUbmiffkIKdJK6SjFcSPHVtELSw+5OWb4OYoTCPDwd75mzW/k6v8tR62A5eHuD7vVqwTndC
UpH6oMLDxGEx36pW04spCwHMjVS3QVY/Xv830H5A1pABtwKEC2/w8uRZ+duIav0r3GnYJlg4vf51
tK7CR12vLJjHTbI6xSDZX4lzZ7jQ3xiwPdkfvVlpMmpm1pp7s9AisGBOMka1TfkcMklZmRbwYh+T
77DdUhpj3m1LifgbsGYD3yzgtCysGX6kdInEBqnlSsrgWkLffN3fq2K3QyGv9OevtHvMgke2EP8e
LgC2oDT2uzT8/HGAzmkdoXVMvH2tRzHGNeFes2aMVBNIZY0QNZD+k0ZzYaBPyeyWFQ4lo1vcL9+U
qfOGwMd/QsCzg71ncBmzDkK3JSM3xKHSTBO3nsiQNCYEpZMS0Olqi54sYloUM8nOj2WnPazlca/0
0iVQZDuY38hAOgBIinV9h7jub3E3sXwNALiB1wUzs+CBuwpwgL0YxI7iQAv75NJOaKOn1/NjAQFH
ndT5brsg3TfZGG8zXQM9eBxBEQnefG5hYe17LdwgyZxsvB5ZL57bER2Esy5Mptf65IR8dt+xWERH
UCkhHq1EMJwBAnfsSggTjZS5pcsKzd12+D8h2m28BldUghN1kGnM4mpTSRtebv68wnQkFYYLkmLg
C04oaBz3Ur6rvFs58m9kfQx2/sm3rTMAYZiUaIeTt4WAiGETRzGApaX0lz/k/6BMifDohHGEIwRL
cMDmbUjHU+JrHpZVwIKKNouVKZwgyvh/dD4NZ7igZiGFw2AdUOeRHsW3gStIvYeIDUfnxC3TpUsZ
mkx/uoA6/kVXyg9KJebhaqumIfyBM+nGpgRn0v9QH5WVLULC5vtddC2JYUIRhUinGNA+Ep2SI1n3
uMYZGxudKUT/AusJLqTtSP9kUrn7EXGmIkdunr04m572AVPJ24fosFhQikCkQr5r3Ko+OxiJ+szy
khrXc35FTcm3VS+lLb+JDg4NY93kAFJTd+KjT5tOU+xH6qCfGjsKmCozA3qjsSdCWu6/AoiFK1bA
NOan2TCv3elJ2YqZYOBFIvLQK/R7/OVN7qhnSxsn2AV36+L7Yzg0ufDUDbpiGZz4qxVP5QfCPYjc
SGefNpAMODZvi9YZEqk0xbmrZpox9njBFIdENWhwA0+KdxC9xahoM5DVFhgarVldlL3f3BWwChv7
p4lH6GIhbNLKrM2iaGHDPhzZNI82a8EtCT5sQsEXf0MCOezuLXUtd+4hnz1opU0ONgJHXX7tq2nC
pm04UYZYhZnLFBax+MVWlZ1cmDbZqHn+dnnAfKZo/k4fT1M+j/5sWTionqXDL1LuZzGj0oxTKf0t
t60nCnerYpgUblpnutBafOqA7kA9aLGThDxNIMFQZMGCcQWZ/F0bDrBD6pfAXwsrsEtnyJaB/H+C
91E/MRBfmkzTkDQ5e+A0RSz25nPKID42T8+KKJlb10SJIOTEg/s4Q13gjQyQF/lt/oYJU1PL/bAh
DYjSBAgzi50rv8fzNyqMBcDy7S+GPGreiSTkxzCzHqKjUok/rvjzoXr8E8UWVXIZYYuf5JUteEPe
4Dp/X7g7kI1BgKcsHrFwFX3CXjpez7OQv1LNU9Kwb34/E2s72URGL61uXEOoZNuYU3K8GADm59fC
svJAVQ58pRb9ZGQwVTKKF4npzFxj4lnC+ulH1+1ACe6k8x81uYBliZpnds2gh16tKVOfbU/QpMXe
lpmqi8i3u/r7dTwr/cxoah2TNA3WWcrkfxE2JXzHzZxHHm6yUWV9MrT1MDg7/+heAjqpuEM5XrjX
j2q5zS8QcxWCNabWeopcEzmVZFScw86gSv94S4awFPWNKAXGMoyu7VGs++WyCPQtGVsJaAGLweBe
u9bY4tammTjH7KbgeDnUgUCkMas9nwUyJj5pd5K4zsj8zcIAKP2BqwGS9bqeisUWx5ZxkCwkLBPI
h1EWNnwE7mHR4mHcw+WA4DwW3C2iooUBE8KhricdHo4SG4wcnaBS8WiT+S0tAevsORcb5rXdUznL
SF0edrZixirCEQwfN4uzaFmLm+2y6FIa+ioDuBLnPOSdEFPbSPHEVIn2i+6lO4l6LneYH0uxAsHX
SP1oFrI2tT2HexzfYJNf21x6Sn2EKHqxOGGV6ZjMYZL3MQdFFOzK54j/hF2q5pn8ZSo9r/sFlGM0
yQnGVvyrjm+Pzb1OfbjrdCxzqPceAwdvZ+o0ff9LOHmHKdp+n9LSmMjiR04PqqY/hFNo7VQ9pDC3
ihxGpXPR+yiUZ8TYCzmhk6xZQAAjLEMdC3A8jwUQnybcJCGQzWC6OwX8tBdNzLCIPTX1lYAwwbhF
FpHkujVa0ifYbSF9dZUsTNp13bM4z3xTBitLNX3jAeLBfWPr3oVrgG/C0xzjoBMvC6HZLpg2Lt+0
zuVBg5WxRmzMy5agfmLYAByqahaTh5+GFaxzFaD/CpKWN+nakQ339k7VQAJ3dbD3a+bu64py02wo
+QqBQ1371GRHNAqr5R0bOIA3EtT28/BErkpCDi2jWnJo+K0tlCnKm8eMnapYZ65vjMoFm+Znul+X
eyIEyH/XbkhUUdtwP7vjx6rRL5sk4PtPC4dHkc338j4f8xyE7vqQ0rgooYdIc7ohqtpdsaIkpBaY
giGm3PxEbv4C2NOeHhCIVr1PvvHmBGHuEq4cI0sXVjRagDuZ+f/pNzfeIgj5cVBn9wxL5KxlY4Wd
J9Txc5uwO1d8SsDdPmiB1hD43zw87sFT8tMUCvtwtVXJJ8q7vYOcLYhKPpNG0zKPOfc9C9ZdADAb
89IoayVasGp/VMfgwZl/HoZ1PZJEy2Gun4tdeZJbVBksYrc65m9Zw720tRVzBPO8ON8yH52kk6sd
wivBli0YBspWb5u8g0f4Ygl/2I1ct3rrpHSl1RQaMe0wAErOOkygryH+nsxPpoZlF+Vy6SXPKH9h
ECZHuBQaUIvNIY3knqSlTV63K5pSxOXbm7tOevXCC08Hp+XVLTqUwpq8OxF7cSy3wQsZz5ppFZoP
xRZ0jVOD90gKbS2n3hd+rfgIXM7fKJh3zeey8eFxRzcnDL9Kr1M//kWNHyf3FGIBovSrjtYRdD3k
Y5CPrFLC2ySsv6XCuE5+aoxgvPYBNFeCMG7bOK+Efgyaq8uLZd7/Ogp/LfSk+6Q9cPTomUYTl2HA
cxxBr7xXyQdXUNHkkmgESNUvTzIvVMs+3oNJzbdwzfzFmgAaMPAA6m4NqKBbpIj6dxv9oLt0g1pk
vCU4yEJDfLNBZTAVjM4IgkS/LpE4p3Pz0qvq9pb8aZl5KXl07GWzGyEGacih+vDCvJAJNMAY1HKM
Xq037/RmvLv+bB1eZvcphjSd3cZ6ro5+ddW0yvgeQSzx8B95vJ354tUuhp1dT1b6L0vqJD4iSfhP
BwLOE50+0D0cGSZ/3/563ixIKb3TcafBPjQukQ/dLlNgt1yy/VC6wKfgpvMqdUmMez/Ao30SdyGZ
shROS6u1U/ZwLqnRyQeUvkCZQn40mSmYyQFlbYLWs6jPIaQ9Hr4i7wTU2RLMq+XDDshKu3MIhwpu
IOF51VnOP2ezbbLWeC1NXY1jVBqDbOg20A+G22g4zzz3AKONWKfeUcFEouJjMJcVJ3Kb4LhA6Tzi
6cc+QJ202lA4oAuicnTQkLS62uurL3zHsDcC/8iQ01yk7VEOZpBLrL89MQPJFw7WsSgXNm8TEA/G
4whX/GFahOzj0BmP/6PygpKDqigPJhUl6Yw6ev1KOa3ThVJzFadGfUh/iJbx3XCiYaF/dbOlfD/B
06FU0GhR0nwlMywCVyJkqSf80Vkqv0OhMooFViXBueBF1bQXjVR1D200Qs00hH2iepmJlBjqaK3q
qbYGmth/0lBjTG6+MyWRfw66EyuuYd2rh7ISsZsQh3TXocoHIGTTvAIYUn67pi/OqNEktf6OzcNf
Y4arXaF/sXIfiibqnbr0DtR6isjvGzHW3mhzLfsTZCWDydE3xNd1kjliOVDPWj5fegYgy4wrfLaz
+JDHrR8Cdr5lE2Kdx1yE1ApuaohYuHjXsl9TB9rcCOWMTSngZrjkLCLuzTBnU5U2Axh4yWhhLayz
puitxvXcY1BozzNdH36uqbwxrZ5ziOLEnjO3uiMWui5LgVF8fvvNiURZrtHl2siV/JhC8nRYDDhW
oxi58d/hlc+InC+6KoLYz+Yw5vvGsse4deh9G1AigwWO0sHZg+DlNN8gP2gnmWo5sBHiFKxZrSjd
NZjpO3pyHaQpDpbNEiXJSznRPd+NV/VPs64yluAi1w4qhtWZTSaADHVseeyLYf+/iuJglY0k6ShY
40xPL6zjMHbsNE5SHXauBmMtv/6psSN99o6VDpfnlJKpRTQC6QnqiIAmeAaRaS1ZgcHVQ1+27G9C
1IpC0p+mcluT/8HdXq5ga8U2cNXjjylzn5Mk8GjWy7evCroCI2Ch/CLjsmWsfUDilTchWdHZ+udi
kzyA5iNIoFamPf3TenU6aXRxRAu1rpul0FVJwJRCKSofVd22/pU3fq94Cv4fg1BwEaGiyv737aww
srSaPwgwqglgR4OhNDcZQJocfc1uJEyHAKnFbIp9QGMJnxn7yaNqYURXtjv03AIDHlR+ABoQ/Jwi
F+L4TUP1SwO7QnYmIjbZfMuCJxikOmwefk5QScPio8cQsaD3WtIr4p4IqCo9imZZ/YLQWE6g/RpF
hpWI6VPXZzEFC344Cd8SJnPJrWlaCqgF9Hrxlx/3iqjk32bVIa0+oH3yS2vThFve95FwS1AHssQ6
rwtm1jJNMRTRVsWTNPasKwv7SrJPJ2SErWS458jYRiPBnpxUfwhwMpoxCRO39+XKhYP4fr2Qh2Sv
R2t34seO1nDduXjeW46gFkHM77uHQx55ffdIFpIjZPbYVZB//hjJnjl06+9U3egY4GrqBfdrQaH1
/Hevf5yiI7zhA1eTIBWXy0q5tunXccHaKlTvDxhCWtL5NMGH+l1nMA8AK4vfzOt0+05ANASSJMdW
/8jZAvI0D3XjZG6niCaOoLOwu24CgBEUSk2FQejcTQ1wiXjVTEZim6SsApuvFcuZtslBHcd6R7hi
dzZJZ8Eh9oXVmA2ui3+IhTuDGcD/B5wyIivPMTcm4AZUIPM8nUutnNnery4ko+NrVyRUAjXPtYUe
zTE7SGJZv46D4kni7u7t/sC3RVo+pnDNpYozu4X0ISnAsAAicRGorM91rhZtYKvky3IO8sOJ254P
RAQ7tGODxYgT11/m3t6M1YtRbrnmZfUZNsAs7RV096jx
`protect end_protected
